`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
FqauidulSSdno6Qx2+wZ+9Q01Gx52At6fmyo7SM0PROVmOgw2xtejjRUvvm0XAHR
UGxRAzca3LSJpL0PDrim1mxBgxC2bmhRfjtJ8+0WtT0dhJvUYTONzMkIabpaxaVc
pa1nfRbW7R0FHg+/rqsOesKNEZnsSgE7Pk1X3fH9+MGyR8vymszyftmsQmA7a0yF
QzYKtm7ou5jym8HiMvKYRKllJu40otj3/6othmgDoCbiKkBQyZ+hVHK43DVzoeM4
CCE92eZOvND4RLctlP1q66IUxBGfF94Q7hB5GArnBxrmK5esGWsrOWClU+lybrUh
U70wapybajo66Je/I4nN9Vuoo6gtNuroc8Lb4HZeOdImHG+OJP1Mw8HJquoDXo3p
cNrI58WNN2l4TWwzIDu612cGpIG+GuFmp3/BpVzaZbV2A244hJtRR9xSeY7PGvu2
pB0RzUVn4PNPKaTQr12U2CoALlodQDk2AjOBtJKdniivEB3ihIXNSrIiNWJ4cqOv
/xF7efZ6DOz3sbTU8ZPhj4OaHxFKLlP1LmkOZUDNdPY8c7X/T6isuIuH6zmbQNEm
GPHrphRmIhgXzlDcNsKwNMaevV1lplDvWb9dCQj4HkS2XffO2Y2DdW/dGeEj6sEH
K7RzBfzhh9+RQ4d+IPDshUSdVQ5YsVvNluMnQrNMpmoEy7acgfbZhz2vCptx9uPN
/ohIZDtVlIZl4MqkwxZHz7vivOe/jCsoloF0B3cb1Glt1Pa0zWLHdYiqsLnAL9zC
eZKsW4O5qs/L1RFyHhzqPZmNhAqx3O0gBuIAt/edon2suKG99JkmYjuuMHjwBXnS
No/DNaXhAhMOR6dJQGl8dkYtjg7+pN5AWm+plMfc/2+T3TCuWwfGdw4N1AuUJUdk
SqnxtJKC5rviBHWayu3adi+p5BnMsTO1wPfqGgJ4X6DW7OYB3Kk4ENQpnCl5Z+yu
oUKotmX8lNFDY/VMYgXPfGevFbFXybpG+ozOMu3RAff/p7a/s3LrF+5Df9Qcn+TV
eLa6eE8oEgvl2fKxX2fYzKPc9MoMq7e03VKbiEI+RzR1dj4GqQeDwGZb7qzf3VTI
nS11IAVRvavLMHacK29VAqgbM8DDEwK55PNmmDYHCo/qQR35Lh8aoI16asl104CE
OuZ4v6Ff90VUl8zSbE6DJue/gTs38Q14KiCWMvrF8QKHPZf8PE24XV1mMDcF2wes
/Y2jDIzBQWXYxyeYeIwgFWa7JEAYQCZohu3LoBMXbBhFJkfnrC78BB50edU4GjAG
cyo9k4zl+FpGO0cvCLS+Kq4e4/KWM3h0EJDVT1+PObTENTqDmmFIVz0c3YL1pxOQ
edqi9avkRC2o4VzReCdxoKitTSJwVX9A9nJKco863NvF2mUa2CqD4BRHvCzBfF8d
GJoELo5RugxkszAsPD7M3L1qFyum82qnNsnQUrLpzN86eTvXUR9Ti8/U7FZDLsSj
4WDhoG16GqStqfUuvoxyp9dVpHo6TcMRM0nduRn1+XyPNUpPgN8Dx8L3OUUWP7a0
JzvloyG57a1ekABQ+8QCiRlshxtIRRtiQu8EGqiezBgMpVu18KLHYzTTCxXd3hdK
82/UzA7ewPZJ4BzACBKcMPLznb5tl5yMkc6LoVrWS/z1pjqALnpfLaxe+Swllp6E
9nPapF+n76kqDWSmcIK3McfCGctWgIT2a17DajiPRPGwr1JZSshjQozpt23Jac15
/wNhsqAXq0EDO0kf2HHRtzXPzGiNBXsmzKrFKQysA/YGofQl+Qk86FvZTMRDRwyx
fX1c8Giq5gVLzD3qrcNJ7eoe8v8K4dlKuAfOt8F1MFqIwG4XAjNlVW7GfpOWZk+Q
OkYCZ/WT6nSYORAZVccAXFkUSj21EAyhpFqnyIKplonUU8YtyZDnPl92TXWoOqg7
2nbeFydoxhSwdqv7M38TisBe6RMmpE7XRxvz6BV1fAwX+GjtbtiBA335dukIDWAH
uqRFzrNcbVLM/+x5WllHRKMCPPVdpVbWoKON24ioGPure7muDCI/w22A3UVypuFs
m933xXNIs3m9t46xqzeJEgQT6zjeugip5rraE93TxHJZ2vllYLbdIw9QMXiRxh09
FEharRugwK/M5N1dDnCI0HNb435WJcgEpRNj5U2hZtw=
`protect END_PROTECTED
