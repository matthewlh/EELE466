`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Hj7KKEgRL1Rd1LUNMdA5hl4Bhb4BogkBjkmh4UPjZcp/0hznVCEHyxGkdNoU8PZS
qxieyfH7dBkYOm1KMl7v0UHwxuq6l4sFtslImnU6mBYztSaEShacAEHjNHcAxppi
GpewAGLe3uKi5hNvlVHTPwup7YjU00IEJrk7KIKku9NhIDKmSDEt5YUKU5Cu+JJf
QhBpkTjCrqTgBe+INHQxW8vI7LAXvd9Va8FfBqGo3+dyVhkhqoji8jFMUVfvLqdS
7JtFV5vqBLEYz6M4czy86VleRzbLfTrRak/tbd11pjX8e2LrVLDPjgu9H6safbpL
13Na3aXS5AwqSTHwnK8gowJXykJyqoHTLVeWB4YcRuMpR0e3F++fRl1eb+xDGfMn
`protect END_PROTECTED
