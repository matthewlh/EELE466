`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Aeli0cU/SQKhewCUVzVSdwVITiTjeQHBfg8HhOpuAEyY1Z61EuhkHfaZLS723M/J
BOeeqN5THaK0uJ78+ZfuWh8P6wK/g9/QkLASEKQlTpb8IxFAPd/VFA62KTyJ8SC1
XYxT/h2ISgSVCJl9nr/tziny7RmlpZ8OG6YmEKeO0xQhpQPUT6BGSNd4pJIMe6EM
4qkwdYPsuOMGwxuVw3B3L3sCe+oQWaqfZpzOPsdgiaZMg1qtsPbO1byTMDmHMp91
QjAgzHBIlUloAh4FFA3ezEQfMb2PYYlDSkVprg2TPf0/nFS4hwQQHF60KzR70sf9
axD8nbeWtV3labn/dN3nJFzUMQgiUtpx27eFgudgAHRq9pcMz6hTQdFHXybYz2zs
mm41tgprn+5UrfRe4CLrJUNNMlxyHyvaau2ph2lyaYygGOQdfoK7gkGxN6hMNXk8
+OGpXf4b3hSqgAa6LxkwbvmGQo8a1+H5x66r2CrK3RG4GhAXKMgLv8ssIkqc0ixT
8J5yxNzSUjxBxYqn5z6KbJQQ6MoXnniE/vTIRuF/VNyGTlVv9itzuAzM6Mz6N16d
96JAHqd1g/632pt5bRxbdsENgnJjDH7SA5Te3uloExvVzSUCD8yVU0dYSw0lykZw
oPMo8xXwgZZzom5hR6I4WdPhpxaChNMtUG3VLPAGOh8TFKcrgoalmkbx/MP+vVmd
B50pvd1xZUeLgJxPlEsLFaccqMaJ/GsU207w3TcvN49+nSps1ZwtJoBE/wm15hO1
G6Hh7+gtxt+Mw4nPwKll31dyf9C/+4RLLx0YhIzkN4apx8rkZCAr2pSaQEPm71bV
OKnGAybjUtFv24HkQ2awl+grkIIr5OWOYf9Ok4Z9QxJVOI+aE9RhYdTmUYR0kpxg
KO99uTsfuTQkBAJ9YPqu8d5iGQkGXvwRW5I25iS+M/lWoyKvqp7FWLNj8n4Il7zc
AVtEeU2oVEiXmAik2pMtaS7zS1y64EKzzVvcFSIR/pUbQW4svJsA1GxhBkwLcHbZ
Wj2LB8LCHP4LiPT/GG26ICa3RH2JN4WT5fWdOE4KgVpW3Sbds8JK6LzobDX0kHnT
jPKFFYPsN3EYZFRYGQvu56u7zg3T4y9qAVzlRQTFHEdJzF7eNXa6LlgwgXVU0/uV
WfrQpzIVCvuqHBu4h3Vs/0kNXfEZOyEF2EDuI1wHQRkS98TxzZa4eXaiORpoWA/J
msLlaFoALGd4r3TqW4gmABTtCUREAoOE/OY5h/xmheFARAq8lzCeJCguCJFTehGP
rAoK72MsNSyV96XaPuXjp8bk+Wns92u6hL38QiPfQ8rncRnm+4NpkahFIv9gJITb
w/iRNOGUU/c4SNqOzlzyOUzijr4KG47psDQKAcJoaJDknYCZu3pinU0R+q/kTevz
y4V9IUoDha1kaUSloENiFIGetsiyZNd9WPWuclqWwbFf04FSy3DmmdTDgUUVgtSL
ROui331rjZi8OcqQ/UUr0FoNqoqNPWCPyv6w8gdEaUEXaYQryjRQ//mzpi/eUQmp
H4nSD5TmQT6DujGBfZGF0sggc2MnqqzEGIDjuvMfyuntQsc6hZSKouZ6RqI31tDt
ne9doU7a1Q4WxunQ5Q+iYfC/WNGPydtker1oK2N9vnRqlR5x3/cCVvF6fP0KkKa/
gde8AqpeU7fyOvgF5jlJoSjYBVSRB6UpuNYhsQpPH2c8XMWGh2ThrGRmfumE8qjr
zjfKUXjILW/oDPxXRfS7T6DjsY3b5wntUunSIQJe/NAbbY95y30FR9Pjq46MQ6kg
TT8xREASObdxk+EYz3e7DgIiGHQEN1Kr+6qyGHfZJ71nFNDSvuobW1uK79c4VNCU
B1cQEbJynr8Jld+/GbCdKs/qSHDLG+xgLZQvh8FWi30k77zFoJchlO4mICggAucv
QHKc8U52M+/xxsqm5TpBVU6dJLr6BovuIwA6iAkGF+Qt9FQmlxZJmuPJegUIR9hl
xfZA/QiX0wT1nemgB1DG5xNnFV0XNQ0yXXXvcZ9IQyIAyWDVIfM3YvojCGtrTU0x
XM2TQJObJK/3PCiGxMiUWmO315WHSpSCgf5HTOfwVRjk0prkC6wUpi1wZQlYMQ60
hNeKHEi/rDbh54fdSJTOdz0Dpg5MMlXthMW4w6L7KXPzkeuUb8tHO9lCk3Sc+J+7
UFNHt7Y7PJhEQ97hXq18Nvuq6EORYG+lZciX4uyHbrFAMEOtWBVfOnX4yTvoNjxA
eOidJ32P1hYeyXRHtC5ABZxqzktj0FEKnsO5zRBQ/2XwH/9nXZXNJPEkE2OF2BET
V2n+S+QItAOVfgO6YZcvcoSL1+ADyLmOZlJk872pea5oKCZgWd6r621ysCNDD6Iv
/GHF7f0OKJGAw2Ov9cQop9IYHZyMV0Z/ZaAsI7oPnrlOKnvyq6SWp5tcuomBJnOH
WZmkRk8PcmCj6PtzToiItS180HP2ObffNUtpP9sJsyRhHUJxgjYlDe9V0ZOGGBK0
MSx+URT3vUvL6kBbYkTZqjVKFibnb72oFV9RvGMHd0O0R1uMKpaoo8H0C63atdEO
qSxHnZkoccZwZRHXb9Ia4uWSUfdDJYwhOYmElq065MM+VQNZbeImsUG9xSySR1PW
FhQePJe67qKdjGCvu0M3ZNbzk6z0gUHgJl4tQaNKCVQDzW6Qo435o/rUcTkwx5Nk
dPCWd30lh4yVU0H+lfnefsr+P/tmtoavBfEf9IgAUQGND/Fy4huIVBYW7RaHcJzn
rkIZrBtSOWQ0jEQ9Nax6r4Mm3YW6rRpy5UdoBkSDNUbiTl5rLAwTz+yhkD8E/IqE
a0SAwK0RxoMNtXgPLgm/xHF2aB+vbx846ZZcyjaEBkgwb4vDte5Yf12FeWhBC4c8
h01wh+aSkFPBqUZKIE6AOHvjAyLthuhK9DcOAvR1ehpcBmsjzGTIQf7jVuUE1URI
V7YTOW4RmcvHRSQpS1R72Q+v/7L+yD/K/NYomViugxtrcOj5/wpKOv8LBII0Hy86
nMS+b1SJ9WNeEHQK3tmT1CFhu9fztAn/bHfsy7eG+nB2qbMArmSOsoe0G8lB6O03
G9a38zNOm0ufJJNuxhwgxv3WEq00edegaWF24Lnmaj12YO/KKpQN+FlqzmVX3VqS
cb6DdpoJc6iC4Ar9fJ/WubW6UJVW5Bqq7Cp/5GCNQrOGtolT9vb8CecndyVgcyPZ
tFDrU0Z6bVcPXDe96oiMS6hsmp+OMSNSCh52n0E5Kh6vWyuX89l0bMviGwgqj1Lc
Ybl9LFjCT98yHDPy/nG7kM4FWAIUWBg4RPWwToGCy16knw2T++CNiqrUHozELDlr
+sz/HEiKIslpdi8QusJtRW8ZFsXMIQRuius4aBEJ9RoY/zEWx+6GaxD9UdieGVrR
OLR/suN18Ba64MPb1YghKGkmiKWw2eqQWcv/NhNDcUAblBfmaRLQwO84Cs35Yvuo
xQi57jeirooct3SFqmTL+XekBE078yXWjD9Kuz57h7bbr/RMFdOC/f9OzMuKqY0U
3158uzi8kXqNluYCE/D4HSHOjQjsmi6XvFrgPu9x3him4tOXLoNHZhNavLfDLAxe
FBYopcjN7SqHDCZKKbkDVOZBLhOeY+2XYoqrGtObhNQl5s6TSvYhLJF3k/C20VlR
qShVN31aBPDewYBwXL0CnPOc6yN9cXfIxgl/UNhN6OSTfCiQuKh5FUxkSNysZLJl
bS30UcGVwoBAG0YKKS9tPw3WELJswaW0ktnlONn3ESJMPjwEBaPf/ELegPA9upXv
PelR0yZXje4Yxn9flNZYCEjBZZ8vvWkPLBOkEFUnlIdqGoI3+Ll1/ZUi4WmDyEnt
g/Ilc43aJIGpLLkAg7C0cQ6qYUQE4oAWHWkfVsK2nf8h7MFwkebP0piJ+ifDKV8L
HupzozU/3BNLjvh0teuDs85WD1fwHdUihYbnXXPm1Bp50vy+gyYKw5ycUngm0NLe
VKYukfFaOi9wVAfr4mSWFKoaTEOONk3ndecrrnjSBQwkJ6L/rfj0tnqqYvi18oNC
2MTkv45cWENbbA9oP/xGwyLMHRz2rJMrTbCu9oBzP7WHg0YHIMg1JnoipFSKk6eu
fFl2jRWH4KoMV5cLLbQ/bmKKcTkv2lGIvVf46OhxwQfQRhP8ZaZt21rFY92FDO1L
A3Sd/Jq8ors7Cdt3ImuIuOxgti7c1yPKJA11mfy6QrPtsXSfYo+YIyI2MqF1mAVV
slRN22AbayUUb1asUscp4Qpz5uhfbhzxCZRHVHVFjZBeMB2VMCY2wglJXhseeFmX
uAiyF+r0AT+8WGzbYb2pAEauOwNE7jPbln1/rFT6WEg/dcwKOeIoKvYnTJxgTjtw
lysbvyDBRL7r3nr7bz8I1XLD9lTS+PSFiRTs+GG0fJvGlCg5rKgrJLA8Utyih/kC
ykXv7XvxCcBTM7DXn4tNzZ6MzRISIjtKdh7MQNYpuH1yVw0gNw5fgrgIhesuVzZE
zniRMmIImaMWeiICFE2nQbEAnYuA1lH4uX5n+6B+mw3umWryyGCYYR2YBJdYN/M1
VYLzt/8xZDAqu45OEAcHvpf//KmA9nPkFz9nu91y0cgkAprNgc6e9rNFCQSOa4s6
jTh71QnFASCmpVkVQp+Ia43UHCg2lPtUdwgeFlt8T7kpEWH+V+z2B662+cyOGNZQ
vLPlp+yOVn5/Q2xHog37YcCAB0ShWAO7/zITXBt2TPvH87m3RZKgGMyqGhnD54XS
YCOJIBw1YsmOIrD9b+fEtxj42QCyFFEJF87bWE6zK6mlU5fyP5nPIJzdjoy1EvBV
a4rFDK1oX0x4CBM+UFJcqSZGOdmMLoEeTQbAgz7FtewJjL+ChytLznuwyaYFuuEQ
1eSujCJs33n2/Tz2RuOqYsmEZ5Cr7F9AUhq8/uC+HRYucYfpriValJIK64AjIFxn
nEt3xtsXEsHb8BQpTCd3pRFeXkeStCW7uvIQJeWfq5DQ1/W0FuUI+FQommT5oU1i
MhZK1DPXhTyyiuxbijaOXlDqLwS+PtXGOoObq/PVRw3vuOvJWLJgKZ+zGtBSaNRJ
Rhdb+dlQLIcvJeR2+Yia+Js9d3xjszsdNa+44uy9bWhTROoo7Ixc4q3pnndgkY2I
nwNF2MtBvYawE69O3fEdQ4/45fkJu2ajs9siIYocCdxqquTK5rSbtpbBw68JNPPU
C4e1dwyS50KkIK/grArxQF9zIkTcMQZJQioZCdi8OuSvSSgWSdpqLMGv2FtsCwfD
U0nMQxt5qh6KTPCp5Au2fiUiOhApA2mS3BEuOeXa88cD5AoSPDU21fT3hLqfQ2A3
uP6Z8iSTL/dZlnYH/91e/o8D6r+VnidVXnlj8Qwg57tbIHJ0SUPAj7ga68Dkk27d
puJIgiXfreuMdCu8eBttMO4ZG4AqwGAcwlq5x5FyBAst25bVx0nD5gffnPd2N40H
/w9i9NthIsvSeNL80Wl0+5lW0fMuYtobLo7//XjLEjsKT8tU/b01A1+QcIGb0ZMB
hsRh2S1BaXts63v7iefwV5U+kJPIenDoIzIttjq3ZurnD7Y1rdSdpCHwVuWye20+
4MZ5GClDWj7sC2xN8xvkUsriiX1+w27TN3v1rUF1a1zWWhHBgFjtS1Bgpa6yaWdn
7rQeV0nTKsLohcshtlAQzjzdHrgwVlz/OmhggXrh9iz9WI0LKk7XQZXtHDrFQ3bA
1D3LL5pVISVLKWLsIPMYfmzAA2DrkJ7AjE0jh55oPazF0hebwXhCNnPMgo0sLE6A
SJgqwxCWSUmtEvoh2bWIUs1AO4iCsBTSXlNQJjQPLJetGW+1TI1ukMLNbjswYgy0
XciK8BPe4qJd53759Aob1NxbRWel/ikV2RV+O627fz6L4fWKhf6y48K6HGFcXPEy
7EXRbFg5gs/uTCf5fwO0AuvN6rtRrQ1CgUo7QflB67LtcStj0J2D29VZDlcD5SK9
oYMH5VKUI/xTJPMAFCUzsO37wHBhltunboAfjGwgupC1yCIeU22tQhQhwby5hsHg
qRgKWGzEAGLeE/tNYjQbMMa1rEUTyTNygiwqF1YkXVWWYjE+HaQWshIToOvBTbkT
WH0Fc4q7WYdP2GitRaGBjsWvxh4wnoCGKVPmx78vccStk2hFlUYFgueBEK2Vlz8X
glL7jpYks58yBUDrAZsEK1oLG4C9TrGfnXnVChp6UoCsymTpNxhpMpGNuzPjtLz7
Gg6Kexc2Ngi10QKS80XYuTSHSqrtlaxdPEA+te44SKluFKxpYBC04nK1v6PfFxWn
QNt1Mjwe8Yw8cQun0YMLmn/mvThSzGMt0ryDk2YW3da9AjhNpGE7F+r2nVj/YGc4
GpUmtdJBxV1PtdiaTqMZswgIO8QlaLS2Ygd/fFHsfFIiPPF0UuHwfgGNWTiWdo8o
6BUnKkOO/GkLkjPK2lf0bv9D6G5CWhxKchZ0uhZPCNS15cfqb5TiAYvBu4hjU9xI
t5N5EAI+l/ASSzQcqEyuXKyRfahFGRVsIEnDnFEEGKYmkl8NMTRaB5E7zsG9pX+/
H3Zmssnwkftco1sXvRxxgGdmgYLMJvQPAxqsttW/cb2VVJ0h3w42t7pYEcqrjhtp
iwbpZRW1BhQ1YbENvcDiIa0QrgeeAV7Qmgo34SqzQ+HWVMOEvUPYV1vGG2Le4AVu
QrwfR4pyV14TsF+CPoZb+tcpC0tuRyAO3IYJYgCqiYqfh6rvj/bm8vRKRXKS0TlH
1dEC+DRjZszEbYI6toKb87eekiMjASQuY0iwq/I1zhYFu8Nk+VB0QCX6gEwQ0vuK
Bi6BykkagdrnAvCWSPJNj48sODOSJSN2T5no9oU6PWJ37Ccl8fpwe6THcmWw/frx
RP9J2hAHXK2/1cRiS13GhxM2z06qxYRjO/wTI21dK21t7itx/Nzptabl3HU4GJa4
2nqIITXIHzPc3/PMKoYSASbsJpA7vwsvj5oHfuOdbaPZQMc5L/WhdPbjvJPEm9Ie
vVKUOOOjjScvVE2DiJn404VX1GZqkrxMnb2wkwsHpd1zjBwkD6ejeck/YetI4khm
Kpq2XOv5R5MKk5yrzoO6Gwb76L93tPjcK067P0Hq2KExjNTK8IvM+0j8W/aWH7Xh
1xXdfkjvOnrfq4yzJ7FYWYVJM+FsopVeAiYOBvOGQMf8YcgX5h8S7FGkOHWVTK49
QQmYSNFi8aytNg/SsIPtTqaPiuavl+vKpLQ4r5cWEVSPZ6/w+5QRr5xcahfy65Jp
8qV0gteHGgCLuEpLoaQQGjRy4izJqmCOUK3xoJ77WEJQFkQc967nnG10WFfcgNKg
P/Rihp5NUD4QZ+YyyosRzZNUk6ltWFbug+Kev4WphiCkgS3bObSTssmoD7Pt2fts
fivZkBCbhGyznPFpfpVRHsI+wwAMV0WX+3IXpjkVULtJOktFHjtdRXZSkvBTpGMp
P9WgCHGTiAt14jmoJ/6wtxzercSHk2PLYdGd5WgnMBMV5tkBqK03tKRcU0a59JsL
tsIr71sCiQHCGGsDnpjwdsWKJxKuP4MlnfUSBoxra3stZ+zHxUMU3Wl7MjgOX2Qy
ijZAw59uRSxwtNuf4fm04B6DhvI/1PNil0grmLOsqqFu4WrTvsVGTrnlZ4TH8Nr8
0OWm6N+MmMrmpI7VJMXSRCB4i9jXTMnU+Gm+ye1SkLzpNCmLPIj00xbCavW5/qvG
a/OtmGg7trVf5+PZP5qVd+zH2NxFGSLixPlVPR2FNZMbVnQSiwJyTgkQtt+2OAij
eJXuEoPRaeyU4Pm1WhuFWi5Z9mMW5fQwynYfzkTZeh7suE4KU84tED4Ft4lcKwHt
rslASYGlg59uXDIdswUmydCbCbnmLF1WlOp+X3KQDEoJP3D+IYko/+qZAqADKWhG
JP7sb8af0KvkAlZnXCplpEvY774024cTiWrtaU95yiWAjsXZ7QVhBXKPsQulbrPq
rFsZ/YzcAxNTv5Vy0j2YAcvM0AcyFKvVGOGvuQN78wqzcdpY1trYfvAWIv+3O/nL
vghrSS8eeezB2KRZGwv9dAW4pxnFRtiO+ae0BylXF51WaL6WryVZ/XWbd+nluCH0
WXbPOI1hI6+qpANbro8WwE21G4aACinaUTopbpIXT5chtPv3pxayA4x/eutiXW7/
gfmWOE5zZA7TYyqYGr3CqxVPE4RbcDGQEyV4WtZ8exEMSoFdknpxMIpA5vu7fwoj
sjTmBDuEUBhVdn2SiJhgLRo1b8PRSwUT7/e1pUE22VWD+IlPwnfmp0bNRUJmTmdx
wJIRbvBRDPQoxEWvi6hcjQ8M6B54X0Gbbs8ro55Gr1FZatPKa+yxWy13I44+S4kL
p7tLRopJ02anRhjOvHddJ0BuKy9w9wqFInxfXthL6rkLyG456JGUqnM3mwUvsIMN
D2v8dMcEtRRYb82DgRtdUJYS6bqiM5Jn/o76udbYSdQq6HrfxmdnGvCKVWrmlXqF
w42nqU92foSQUJA9KvvRjqcl0elxK3dWoc9ivWP8xyR8UCP1Io1xhQWgLFcFm+q1
yoUqUZ6Ty21p4IsM2hLTIN5Nd8u8NsgOQFQ84GzWl/kay3lnj8OMmBqdrhHrOjua
u2TQ0hcNXNiwDrdYVPsTLptxBuka618dkTYPf8ZBOuP8DUv619hIiKoP7AF+Lyv9
RcmGM2mlgHJq+hnGx0DdrROvJnpXq7nrP/dBre4iEAYCM/Qw7iXns/6BZRgyyyzQ
LqNfyYjd141C5L2eTcIYF+jpvyEMG2tO7wAWiDqTwMkiJ+w0FElebBdWwBFuff6C
sa8ZG2Gu8q2U96j+bngSfC5n7bo/CASfoAa+UZWoPceG/iTPHOx3DOJo/AgoiETt
jvVzVYk2oBb4yjjupQiXbB6geeVrhNQqkFfPY+Zgo+132BRbBP7Kl3ZyuWKMpc0T
mCOmH26bGkQuhg2IyQJZPQaW1aWFuLook8XDkEMRsa301UeYrT6c5FXiFX0CO1Sm
HBgHbKiSwvlwIE7hIpTg5A61exhwQDezRGADafFWToxL6pm+9RyD11pvm3L5iZfW
YqK3eQXsVmjTsihrjpHhGUHU8J9VD0V22XYe+FvwjqLJBHv+6dEsZv9C/kx2Gki6
0sCePOtcZR8Nu0KYqd61IGH+Hk58fS+xOhnrzgyoOOpjO+Slv0rS4JUO0taCspOZ
DisYoO3z60uKz4PD57Q7oOGmlgRrDTglNRIcGDR3zNQI77lVzva5XDVKrp4TqHXd
OIEVhOVLqe0Gkz/F0a7ExUXOJGTuiO+5VRXJlCFxXCC0M+MJ3DkkFh9L5ruuXQWp
VqTEpmGgtpZzHzQpllRssi9oGhKqN+18cfC93iOziDfyYXcPqQn53rj9QLkePP//
YGMymK2g5uQzr9nnZ+K2EGPKjXi+3LKJEERHhFweL4TcBjKWt8mk7boMuknIlocr
hnRiimHDHs9jYXJhb2rVVHKH7oBX8fb0fXXlfEeX1tnYlTU9l2G7R4KSMU0vQ2I4
BUpNv9IoDdesdH2OQBvX6jJPGzCaN0fCuuFEquTTDqocuJtYwUcfm5fQz7wlvpS3
rZYrT0LwPJgS1POESe3BqB4GdgGT6VNzH60HYLueh20rpq/GmvVpj2Uq//MY58U8
cJmS/c7jYPH/AvDzKCp45dgboUy2X6kZlW8tjZU0HsA9NJQ1yuQEVCEHdVRw7iWA
vAx25vxIpmaWLSeFcEMnznXOjEkykdMRHCtOspXoNebtLpzvGWaxLnCJza6zZ0Kx
r4GMvOmT5uzCyCYtwBKGfusmjjutM12fLhuZsOn6X5fpaSu2SBQytdFl9rHZnFXB
SGrC+Zj7k19Zhy7iI4jp1WhJgYXcBTzWefChi03VLrh4Q0hy10NKk4b6PB9yV8C6
bqm/65k6M6TRSeY/cqOGuegEIMjnIvNlLlhUahQNBhfNDtKGJaDM9RDTX+fV3WBx
/RwBR8A4RQ0QMipNtlC/LkqVhVjhKh6+K2lc9WvkIkaWQ3niuu+av6PqTcuy0G/A
6Cgb7SKUtI3vHc865dSo6aYRw64lxDOpgXwTmyA/qVBe/3ueK2VEbJo3CNKqaclb
ucxwleBWsUGykHU7HvCxd+lJv3pN1aOVso7o7OOdpObr/VvIBFUHGZih2zCXDIjB
nElc/SgtrEBTBAcsMhLZ+g0DEqek7w1KXxRS+naM39d+Mx5+0jlFHPAxFKRos90q
HpKEuH6cUg8LHr+kOGXnifRmSHv6mUXs0aawA/RmemdcTvdymSuWyQWCltiH/yVg
vtC0frTzUb8xmvHhBSdCYh+iM3od6aYflMjp4wBm6uMxXKHR+SDOwONsr52VhBFx
pne7WGVtcZhZDU/9fpJu2rt4C+YqumoWVuGcaJDiT9t9/eibxiQfrPjxGCMg2Ihk
3DPx2pG3eCdBz4mVf5t9gtq6+1tIbXrDtP3MIeUs+nwWB8Xuamjs3hc2dkqiTtwo
6j1ErcTVql1UkzfbLiehwpK60+Te2YmwKvoDLcTIfeJE8SqbEYFiJ7ByNgVSBjYr
kb0KB9O2RgEFquaOqy667eUL3Zf7WAHxMv3UuC+qVFaOM8u7sRjdxZqlvgKKv3Mf
nuOGCi6M0+QyYRlHbF0jTyShh4+vjH2bDEa796+jOPi9gmWZ5NI2ws9gJBQozE8t
WAeUOi4we3bNQsSqDbTjWyM1yyJMhbJfQxHGcAJeSPs+vKaF8tesxGqFPvN9Oocn
1/VNH8Munt6a0K4K3yQVJaoVvS3Bdm5XgKY8qc2Sv1kZqelqDHafb9qUmR1Xup13
EZMW54Hnn7QjOJG/88jU/kdhGP6dDCeM4/zgRRzAAvjazyeQZ9ykJjComJrKpVqI
QK+d35oWR+6C5QSVjxRVlhjE6bjF/9oO/GfP2Sg/Llq9t+7KqEuH8zwL2XKu6nrc
MjB9A63YWFaqqpbOdcW9jmmQ2rxJe9Z+KKXVVClJfQdp94cDjCB51wY46jNYAvcM
Dalus/V+D7PTQHf349Gi63vDV2tzjq0qKZJ6z0g2jcA7Ot2XJ2HbVyRVZEtWy+u6
XE70aCJbqPKSuqh+2MJAk0NQijgHjqpbDhGWi1SSoNFPtBuc9HnsREnJhfIFMbbI
pwR6XsNqkHn9aIKioyDFKH5pE0gfm/4uDWP6m6xJDIBvvDat8QFzpw5CaWvDdlwI
+GN2F7ydRnzsMKn5yBuWP4fy4zJaJkcR7g4UJdb6sOZPY8MSE3B0QtHyUacJ4Pl5
jry51XyAHbg3Q61or/UhZXnCoY0kT48k8SYlcywpXtZEJYXDN95qf8WWrQcLuF0u
UZ+ii7L/DHk3++M8d2k5lSWoIlfa/dcMOyo2xIkloJj3REwwh7TrurOmEBhLMcy6
02WE1yzys05of+rigwNzZ1WjSWybeoJ7C2bpXobS5BQqcQUj3CymxUyxxl03Fuw9
ZA7gDsHAmX4+678OB21/d+yyYtgboJCp1uXci2ZEyrqSfk3G8US4xuOuUzQyVxsq
7QnVSNUunYTGJTpaG2dwG51ylZRAMwbeDsg32mZDk/h0ZI5j5jU199p72+D/EPZP
h6WQaLeNFJTOhXQze/QSNFlDJaGKsYfx9YdGVFHurkkDkXRO7Q1SSwB1iOHqDrKG
TrBUhqpM6USwYzInsOFW9ffSgyr7xGtpLrMz/uJ/81otixC9dmAqayzX8aRIovbS
k4tnTYJigNE4eWS2f4IRA+FzfwiSxkpJDvUQEV1MOuVrp9AWWEBrKNui2faXSBRv
ngUDxdbVP7ZlSWBeTm7I93IjGKDdimaI3Wztv8YZIlqperpk/JbSsTDbaEUjEVgm
OX4fNfdmp5EYORZ4v79Otc0fMQG9yuy10tuWPfxPnSW8eLS5JrMmlp348Lnkr5eR
5G6jGPpU6FhjTlPI2SbhH/JLItHIxYqhiMkRmCJiv7HSZj5lz1ZCFRQLmbJhegtE
TxhGxpuZY3rgSNo/YNgCvxpxoCZq//BAdV8j1NKTt21iGrmPa4ti7yo8gTzEsSUU
snpSpHHRZZd3yQ+n8o6roMYY9friIoQzF838LKjfQuGEQ3Yd4C3+psa9vmzwOzTa
9rxpeW0BEP5f0RfuFa0EnApbqZRTmpfyNygr8D+aeApFDrS/KOTRl6hWbc2bVQw5
KHWU0ui27K9dWq2WsmLVV6SQRgfT5LfbBEIN7nztUFYh/mvG3HPReE2Rsnkhe38W
tFFgi0pWzCCQipL9Rk9Zu3CCSv6mxIle2pf+cTP37cI+m2LA40bCcnW4synhAHuZ
YvxbWHC338NUvPGUk4iXW85+Z/niSVL1tho1UYWGO11ZfXFWDU7C2O8J0kZJXnBl
yCIjXjiwyFkVp/svYC3ZGAc1zXUnYG0HvSgdWPeYnIY5QqShAlsRpU2DLlG6jx8J
11gY47SI5QyJrT9mmUGpRhvaKTjcy5hrSUFGn/8bvSO6IJGf8W7dd2guVpr3Ja5G
zfk5YuZKKEOeemMRIGboYdZLB9TYOYwGsbKJDVvkQCvToW2YRFcSFw9siCEIKx+O
jUbis6qhtBvYvPC5sqS/NGRS78vpYEsd1rSCb+Kc6fr7eYet/txgy7NlSRzWpMyo
3TuAQ7UikalX2V+Bhtqm1plfPODhOWmFahj9t75kXg0voEb8BUtUzOerCpqxlCA7
Vv0KVz/FND3g9l3RBI1pJnEM0pPg+t8EAvWFDz/OHqE3pEua1TuEdjoFD9AxLlt1
l7UyGbkebkFEXWS25NoYXUT1Yyoj1bjeqSxqSV+LEgn/MH34vO8P/0ZuxLWGMlqC
12BYKioLKfo0KWCq9yl9tjgLGPTKM8wRPnicLXpPIqzMbB+uWlbkZLqg5mK42Sl+
11dfBHkMoXwYrXcYeFSueSXHnuAGiNuANul1kao2V2RGoFRdueZD57eh2I+zQFdE
ucoFaNDsTX0YHfOy29+UPNlBdldeJj9SVn4MFDp2weND1J+eJhvvjSoLZlNEevXe
gV9VO5WXjJvDnhmZR1jTPq/CFhEPrCpLCs07NvQeL+xUG1TY8gCHDxsvlsBnNNI9
HH1xiVgeMWzhTtGlau+LoY+DN+ggmPVMHoibrd0UIWF07Wc3CJmCTt9FkMhNW5hH
/Zh/6LZSAf9GuiF4wJYrf4q18rAti9QzyqALl10lLtYhxGTQGrRjwCbaSMhmwt2A
MX4b5k0xZ8Y1gBI5vCz2CHfG/mdo8u004UYqQCl9FTdxOYKpGTip/sg0T08nGPlF
BJqFfRMYGrqgKP+T3udYFjHTzR9iFzF3vBrAfjmlhYF/owiMWrnF0kJ8cOK5mMic
`protect END_PROTECTED
