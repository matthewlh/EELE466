`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Zq1Hk9aOaspfPHxcfzJly1Wv49F6koSgjSLNY5OeF5EhZc0bLlBR/Kr+Hko83ejo
j8LzyUxTN+0Rv+gmnKDde2VX06W8JH7hfJq7ZGqfaYP8MxCTlEnCYqfnv0WuYFbX
pp/cfSI8Dyf2a33q0rRomuzc+XO3GJdzcAL4i+qMLr1lhS4yTIJwZr0KwLaqAVJ/
1yiqCmTw+PoMzRvlbhXA6n2WwCyZ4wMmNPh8edwE4gy+oB6Wfu1d2ZgOL77YI1Ic
H60De2aX7czwxOrB2Q4pNcSdljwJIeLBZrPMz2+pJpSUMSAmBNR6h/1LlyuUn+4a
7arx8WoTHCqcWGyRzTDKJ36EZ4TzHJ8U1uF64myZU/lmmVqG3+fTYDwB5XDZaiof
byo7bc8mQJvOOL205nWzHDI0I/VCVhm8tySD5DMTHI5WEpxaNGX7AgyIegwT5AX7
WEow8u8vFHAgpwCtcEaIzWeN39c+RuMknSUDkasQKaWE+EISpg/UnG+NjbCguQtg
FJ72eJryr4p8JfKyJGU3C2k4Uk7oQngr8T3gbe3CKrDdn2U/WyRmCU4uhyGESkCl
9vsCssd4JO+k1wZTIpzkkkBQ7CADvn0ewWuMm8PdgQ+FkP2ezBP3AoeJQ/mmeXrv
OG9c8wKqF+hUFMDWzKou4G8StL2UszoNr/rRmbxMxxUh0ZFqzX2Iij0AtiZrZUea
p7HKeyAALEuVEN/JitPva9Wa2j5DIr8ctV7h9P99+dSar4RX/yP4IBXzCUO0Ux7y
gNjkppW59eUMyy3kiiryYlDsH826MWp9on5Tzm6sbuUMvOhzE8V4KenBgVHfcdsh
xmmhZ1TEatPZUw91m6oeuaC5xOvyHEP6Qv365CL5UEU4gCNNPBmn1jQcexTp2tO5
dzlURmNxCV0CXjn5yQCijqSZQmsKxFt3ReuS7+VxY+wCd/8NhI7XwA4EK5X6DGFO
PsGu48s+PhZ3tWTmtdA6rt8fRSdp6UfrUqLW7Hr/tamLHVK5tFeuBlZfJr/LHx2z
SivMwcG7kpvy5t5bKshPPbPMAORE8T5dts0ofvqFBYn71vH3lRbw+3SBz8YGMBTp
8XDhJOK5b2WUWB1573QUunsndqLqEMtfiXRCSbgZIS52wYDGS+0bucwHXjvG++ZH
ZBJV27t1SWwJKKXhNCaxvzDhwZyJ7P1WiBJEL37i1nUamw0lRYNxEsfsrrnC0INn
3Dj/B5SADdRnjP7hXFv/421JejGI9pBUwiwyXa6TOw8cTj5bWWSFpD6lA7rUyUDn
IsBscjQl6qZMBiAFguRJsBZ7atShpUxKc+U3Pl/mfpxsimeaJKljGY0Xoe4/gWXx
pGT7n55upXecFJjmw1uJdY/unQHpBmBCBbqmphbX7ZSD7A+OtA1EIUUykyn9pNEC
GrnmoiKe0/5VeiqGNlS3HD1V5yo5iclxvZoxLxzSm55w19YQ8eu1bLSyEDGxrEFN
8SX3YH0FtTA0J7rFoQWL0Pv/xuvuWQ4F0swFr0SdeOLASZNn4HuGSbcdvdBzECRd
q0FGKNkDEA5A1owUK+HC6CDTzhWXkP+TRX+cViF0C8TbAyWOabaThnzbgqwSqyA4
CrffDb4tbgQClhGqWfSOdCYorAjRX8mdKV9UO7QuUNeIoHz5nqoWMoYJYel6HPhw
ACeS2WRD3QqTyDqtoWM4NXKKUXk95IpcrADHnMLHoxuhZLv1V9QWUnm4aoloffIW
yrw4/t0Oq522KvtI2UdknujyFBPilW1dejCL+Xvsq2GCMrmVLY1ghZQ0y17NI8Qp
Yx8ch4v4ixygqEpgEYYyLckZIqka/fznNsGDYUpWncb45PjYxobSSeenKRO/+pm3
gQGyciGz7NO0mvpASsDbUCsa2hcK7E47egtLlLmoHsUjxBM795QUSdWxiUfcb20X
P0KEbpwVDQp3da+B4qRn1efvl5LKsteCyaKuiIyJdY3654L+35eUh48ibR0wbRCO
RkvN/PeO7v+ir1sVRYydVh55eo08w1XgTy4//Ve/2o0/LOyWNOgexYMBonL/lZZz
GC4sOlpLsFebD0eg6goH9vc79vgBUXvG46W6NT57a0JN6HC+5QLZoKM0ap6n7dEg
m5am9sJyPRj/XhVFg1eLEhCqxLyGWxyqN1DAunWyDcRTXTTbHQHQoNWK6qO5X7Gl
bg3boiWo64MBo2AjLTPtnNiLfMUhVUjmUok3fiOUnTcDwCoiDXCeqdtZglUChIs0
yYSoiOLgyDuB4wF6sFsn/chxUANJIXUNkOG3m3owFuhd0jFBuRFL06jpWxvOS2CA
Ez000yaH8qSOq4SDOcCiWtgxdCl2lwUh48zMVE0fhoiSbRoFhibMWRq4bbYta0YJ
RBXPxjNTUimOKvCZk+FFWdo9hdwvHZ+4WdRaY2F7COKdthVgqzflXcOH8dAAlIT9
GoQtdtTv3b9m4pSDw4LflDRzoD1MugzelRcLmtwroDh6vb9493v6zGexPZbGBqO4
ltfLXQ3lapVfTADozw+usGZY1a2/8+x1v4jIU5KbzgwJBwhPmEVvQB9g0FOLSO5h
J2FznwaPTQb62qmPyDF6zbbcdXJd256JHqoMkNwIWZOHZIM9PXb8/fXLqaVNouKI
4Kn3wgUU0Q+/LL0FRADp9gQz+AVSkAl4mQaag7fPZ1NcD9z8G2phtD01b2tKNkIS
R1uYHXLl+3MS8Y0vdF/IK+RPRhHsYZZaGXQXxlIw5/mZrL/AGIGABC1dYgch+UGF
TUVAnr0nr/B9opsSy/qOxgkZzbkNCsUQwvN2qWdYjV5ghDHBIaeuJJhet5EVavIn
Zwot+pBSD5HBpn5jzhHlQZvZa7GN5GmJdoc0dogUiReKcBPQ8r6uI2ctchxgWPPL
chI5CACOP7Vul2fZ8Cr7mbe3uYTR9zgB/08bfTa2JCD9Nx6iCxTJ/pJ5VEcg1KJH
O7gETXJx7FVgp/o6ZV7T55KinCqgmv5Z59MAd4HdG9ZP+a21A1ApbcjzH60FivTN
Q9j17Vcon8yfN89Tm2PZbGIsoETERTheeu4smZI8rG+K5fEgWgmh/At5QV+lPb/X
b4uUtMs8dBsNIFM5Sd4XftU3gARSOafTzxuijsY4vrceWx+QOveZ4G2Pj8nS8YH6
318IcLyfDCRaimIzSp6Nr+OotKnoCPjfKngigIeUL8JJ1jA3EAsV7O4BKITdJpiB
ILtlKwJA3Maj94pG58+eUqJkCNmoSkd1vHz4SRtgqa306tdexPYrVQGD30Fiao+B
BsKdzFAR0qfXBDLTK8s0IaJnSS/OKs1ZC8cqy9W3KxdwRiQSs1oguhQN3PnSBrGZ
LvvzVwksTGszCz2H1hBeAY8SUP/kdZ13bIb3boP5KZOWQdBw926/SdNWVzh1MhZp
o83v74KtciTmoVpxuxN+DBAJNRUa0B6FPeE7i8sQ79k6Hhm5+ZLdz1JsjjDUUFsg
rhJwqO7zZEFRRSp6QQbAx2hTzv57hgx46e7Hx+W5BPx0BuSIGJa/c9hHJnpeNHgV
TuZ7tnowAmocyEfecWJVT22/gzSBdbtKMUsAG7c4TzLG7YgEZkPiFy6/nHGoHgXU
fOBnLJU4DIbKHKoytSctI/3Cvmi/wdIvab0jVTQ+Wb4f2k70xQkpxCbWWkrfYAJN
o1BnvJbgvnjOj3B14PvFnGNdAOT0ypnqsStK6h16Q7s3ooStad+cvMV1rLo6jQDe
lSjvknYKyYmgWaIYuy/sJO0q3sOzquyXUSuIpfO2RfK+Z6sFLmHfIPBoFSIOsVUq
EcitUQJoRwDQZcg82ZPropmMb8mFrpQpCLasx3W0XdvuHwnNX8XVxI5RRCpTrPby
CCfTT/GyT05s3L/qy/nrl9X+y08caluru+cd/ZGciIMHKGPn/icsML8iDXXPcqQ8
Lqa9Cm4U1dHTG/KbQmkUSyaMlBz5KhPrs9FwD7FdIzsLcCk1yJRudp2dzyymxnjP
5i7HNKDTd71djTtnUdPTd8jCdcrj4CTNkjTPmgZbTY8qSdRCYrT3XP3yEVZSLKAq
f1KHFZ0zwWwjsDX0UoWvmCHLmhTfAy20k6tpIHlns0FScttlIDSstq46HLmGVWmu
mK0j3l+HcUCJNR+aQFLBUbuqkM5pwvwQLIhp9GLAc5IMyRHs67sd2hCfN9Lo6pHy
sn7ryxXCP2BmtwaJf112xkJNzpX/fNTOpzJz+Sm3lHfnjsVWO/WNHuaMcb2BjD1x
HyVL5Ii1aX/xuddluT6pbf/QlRHuYxBACgILYMd8Ub3NCcNJEsBhHfiM1QJz8c3c
FEE9xebP0OBAvSFXyOvlLr0JPYZZxNwQvVV09U81CO59tQa0a8IHQOea/5pIWPHa
4ruc9I2W6t+HeyOWwH/FAbgHrRZ5cFuM+LDw8A5XOOoNLt+i9pqYdZnh+hq19Rqy
SGWgz8jzZiS2dUoDz0oYXVpb6pvQzHNdQ/x2LraEzi7652iCRxR2GZLMfwAsPTBI
cf5KjAYtQYKe2Amjo5elihqqwF7vveRANhW154MJXNEl0dIo0jg+TW/j7OFKLjqp
1Xo+xPnI13SqaQnyAPXyjo71j7CQIugEuoSrhwkVLTEtJaCt99IX7cmIM2Fw0FWt
Y2NHthl0jTdQ/87YkaqKwjNCWUd5mcQiKN7lC/rQqakT2Dac1lZ30xvy08ShXY6G
bBRCTyntYBzfg6YqgGw+2d4DBBSEz+JblxPc2D1SsNC5pj+tkzZgYZb2ZnYVqluW
mzl13VjXh21yIEvblHP5mpRFjJHwitpxytGlRhOeviwIigcGzlymPFpbW9cAfFwG
TXRIXjfRiR2YH6lTPz6kDJ4jsTBrMPHoeMw+iRR++BDlrftvS2KGldrjcTqy5OKb
OTS1AsogbuSa1kGnW3O7RL8IAQMC3dltSzvTeTmr/C2mVsSSK/q3f2JAVde90BTr
B+UzdgjjPWUHicle5q3/5mGqBWfZuEtqTXfiZ5nEQpfIxBdPv15w1F8oqYHzJsgy
1b9CiKCs/sr8MJvxSpf+S05zatlVj4hGlLLegmB65KayUQUiKxU5z+nElwFWo1d6
z3L4Ih1qHYF18rjxhlo/K5UYs+gmtXnnH+ptootQk1H5eWR1IIImcUyjsN7TJI7E
toxqjMTnpOBVy9ZYq6E7MO2U9RhizumU953QH3EzHaawlbieNCxqKGtkFDVaILi6
7MTKyA/ZGINLTSMP3U+0xi12xFj37k2QGB03KjZQVnuRRBYXp9eA6qP0M0R7orxK
PViY6mcg/n6KTSetlPu8tb0fI7eG3PWb8fbQyYCbQ06cmuqNmNWohSxAccYeO95V
UIXVSmrxA4CF6zsSdbCf/OA6niR+7Q99PKVY2oqZ5jMDJyPmrUoHIAjDLr62wSUv
niSGD3S6P1VROACIAcOFJz+S0DjbHtZ2wCHupzBHwd6qM8n3i5eLktCmOpiWVu6d
KcKizr7E/5t6MxTPDSFiohU3IG1IzbwXdd6fIBhhzKe82/Hsk52bVvS+VLMpiR/k
AKEutTVodeqstIq7fWqza3mFNiNkVwOoxK/3yeksRmZYYXeB2EechibZR9S4iP1A
d0c/ehsA+uX8CMN477ZFy4ALMM3sqXddcJFa65iCmvDa62CeeyED12SEttoe/leC
cZDpW2plWkNSDFz3kLtrbvdvnYXVfVhK60gGS1DTwlknwTAARpaPsU9mHawFqvFJ
Uy7fR6umjX6eAVc7uKYGSgbVW5zRrwdSQGxJt+DlO84C5XNK7sQBNb5rwCRHcayM
I6jCTnw/P6zSv00kP19oCNDkOJf/ZqfV2ias9I/RkVZXbIsqjnOXvlSE/zYjunEw
kTVvNe9EPG7HTiLHh1dZp7i8Wb2pRZkofM/sLQCjVsG64dt+1XTWie6fiXwuUMCi
aGw0C6eIlKOZ3fMNMl/kjySskXGgjVDt2rNIe4hbAcW1Xd1kGNdR1sAIi3CRVida
Zdz0gJwZNCAZilTSqSA9lDATH+sQ2N91q7aHasLoFJSHQY4iZ3Avc99h4B7QctLm
2ZbyI5CQHifQklettvyeKYi8UB3Qd8GCMGBOHkrf93mjGYh5wPtBYz7Eqr5wqA6L
7ua4qFHGe1SeDe3fVyW0dDKUeuMB1XX1GWt0wlKK3UU7Yvx7t8GcmsOPmK4GwQZg
/fIdZiPBgQ6ntvs4J+1pxs3bVJ0iaJ4DjSTQ2BfjdM3qWWYXR1A3RbD7NoYstvT6
VXgXr4vpoGOHF/kpWtuGIf+gdnTaiLKsVCYnD3jGuUlATy98g6tjN7JLQPM7hny8
PjcYQdEndlCceYhm67gfe2YWHP/qKUf08bxqUMmPkm/sffiL6qETEP1DtyJ53KLR
M27gD79gjpdXetMzR1oD5DoB0Gy2nj8rL6mjxSXB6DjHv+paG1i5b4DhTAbXxAit
eX2imUnfEF/nYRc9ijhDtVYkf4mLAUndKo0Cp+0+KGC7WkYTK8wRDJ2x+hq8JErV
y2iD+qf46R9dNryC07sXnYr98YhAy0nbelJbqq2Tqre+nGWaG5BJ0/UvTuNLqIbO
axVaGRUb7+RvpqdHTDg1Ld2FJTSBxakIW+a0MUyE6Qx2hB6D/IKoMLs0N30G2n9Y
2/3iQtTlENB3+aCFfaByid0darVTi5tgxm1wa1zcbUEjE7Dt0qhKJ7/aSXTZrm9h
s0TYkBoC3nNozsHnEhTsKofBs1dkINbOTczuJSbgtmkB59eLARQOIHa8uW8q8sIM
HrRmELUOaPbP9eNkplIxQwOxEVZ5hE00Hd9V3IZ8M7DbFbPKYUi3Ueb3j0r63O5/
x63b+uI6Qa7a0SsBYsneZOAm1zuxYJeOqOgwcrsladrqLL9/iG9qtEqrMv98MHW3
edBsceGlZELRvEfQ2fAP9r1dnw9GmCXXrk2hb0pQ+N2qBgNzN5necnpu66FWcjdm
n7OEL/N09IA8huIKWpJHyBTfqgtnElk3XQvYMCaSb3zCkhSZsqNcFhDhTdB+iySJ
mosGeZ6Po3uKmAh6xi93tWrPV8X2Twk7Wh93qaGg13nQ0O5MBhvt3oUED7nJojeO
/Aoao5Ty/Iq4wcoHM1SLjSo8sxo7v6PwYhy18/rU0OzRo7gf2znyK0mkkf1ToGNX
dIehdg3YbSGrMWUaeQrIpmYdF9pT89jGiGgh3jB1arib/DsTdl33UrWeKCRb+07P
JG6iokH/cszIvQ2+3EZU5HOhOTmg3xGToD9HM/r1xyqTth3083Xz/76UqPPg++Pr
oM0UB+1f9HIc8SKrZtW6y3W+gQhlZfxApNbWGRypr2KcXem2/YbQT919hj6xkDtN
dsn/mh530IqpW3dRF8uEn3KI5fMMy/ttzSS4foxeOM8OnhSwC0cSnELwkwHzfDy3
8Cvh7f03jzdBorwSavDFt4PiJgs5If2ZvhJAZfG92oToAhmAYXX2Nxoz9MQN59hk
/2vqIHOhjObX8zTjAmCoKLkme2v1CtvMtsNoKD9xz4FtDptpv5BUE61kY2tmE0Ed
cMk6mLDfz8zJKHtZFjo/XRmpwO9v42DO+VRCIoYXQ9ycuqT1gOcvp33gf8OWb15g
zfJizk6wwuBjyGDHlcQ1h2li2Yds1Z+GWDKmp8/AyChks7eqz9D5OSX+lnaITr8+
7dQR4z8cQpy5BqJpwVY+EzHMe8Omtu5Ac6ot4cfOIf6SsMScH+82x0GQ7KHgKZF1
S8+TZwzbR40PNOQetMwvDkN5VkUTkMdRFoP4cwqwsCx0s70iHdrsJVxrSDjCshbx
lYdB3P1orj0RKgCYxB0V6X939XvwTBycLaNzO3Lk1Eii/qX4HP80UwLZBXXtq2Ug
Z2Rdf3Iv5S6r44BSV5g3xuolm4NrDAEb1L6JDMjsNYddTE0AkndTg904pkFhsyR3
XxZGSRRSTcGsOiLR2NQ2JFd8RBgi1fciDTWSzZaG93/oIwxwEgTF2au7f04+DFbN
ayZuwu4aJqqRcg1AYBGdh8FN7Mb9xx2LRIsslW+so0cBTXoKKlQog/FmhyGNOlyH
lMj+zRvOaLQE6hoXgejECqnCiaZXz1WilTzjlTFYiuTUDHf+bKpIKsgQz398SvPW
5W/V5U5heglhDddQ8lQHrbQyYO5kkLrXxHkk2sX5mew=
`protect END_PROTECTED
