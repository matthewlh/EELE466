`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vw4r07f4yUEzfpV88sQrUP7wKEtx3SSRQIH+dhUmtg9RVtaLp6BPMdPglltZFJyS
Z0c17f1k3PcXk0HJYbtG7GHgSs5F7iik6X89/CUn+yCebk2lMo7zl6MpHCMpPqUo
xkF/2eVb29l240iQH+QnLr+8Rw1moLJJaZnnWFkXkXiOFYkcwrcGu3nNA8l+uCIj
9HGbYSs5YO7AcFWslVsmulydwM7qbW4lRpGNyA+/QX8tqPMeK+M34IrKpArnTp4Q
C3gdtNAd+8G4Hh0R4XRInO2nCwMaTBnOn3p4mS9PSzi/RVod2Va/d2ykx79z4ink
QcYVgRfhVm6RcH3ndU+RGPBzFWF0+HtfOvjnBqT5vBXZaC0NnjSDpyZsOZ5HgrwY
gUbCTRbDEB+FDjAUOZu8fIPY+M1pv+kj7h0/DreA1cCOa/9tmqXWCRhbGRYLdNhJ
+yIeBYW4Vq+1rL3w9MZrXUAn+4dt1hlNGkmUgv6Xw/zMrknMF+obBg1HjEo3IG5E
OmAQ6KZm/TOsA5iI7l/q+J0hzHbmphOCBtu3HeKd6aPz/azgv/dNjD5lOi0jd5RJ
f+eBXTkqWTIfqx4Yr5Hfj025sOIRwm8QKJwIGK9cWBeyGj5q77f7cmkifaiyvKRu
w3lHT9lniNa+j1iscqbPsu2se5qwGJoaFrc0lVrwkc1mjlGMhuuQnvxBSrLBioNX
FK6PvPpt5AjNU5r8QRpQ2j2DgSoRslq0pCF7iIHOaNCjlNRORSUy+n2m40YeG6SH
WNip21erDz7YCJIxCQUeV6eztdCY+MYaaYq0Wo6y7J1eahro+aKkOswt0xAtwik+
6hZIm8tzjiB8AB55shye2mJD4fiaa03nd/026JkwbQYgRVtF6lGh9hCdY28qiMte
PqmmkALuxmBHXX8RT9h7MglVo5LGEjoIoDJMhgksyImD+KL/lGq5WRYcJInklDIT
ltzZbH3+wAw2r5rkwHyukkTVRv/titeDrzQiSj0oNmRDcrl8bPKL5KwNPtf/Rric
1CWRwqg27HpUYxbNBFpyR9p4+qQYo766XTi8ZpRgI2OdQRXrYC00TuYDj9QE0xNk
wsnz286QZRrwQS1JGNmJAs0l9dd3kNxc8vUM7pwd9GOtpl/d4v6N2WzQmVyDKDO2
GKtb6kx5N2/ueWgp/0Pnk4vied1Bn9S1C2v3lGi2kUrSwHHK3IvaQody1ni9nhx7
QnRRvZyKZzju2ypxSI0p2+ADRFrFL6XCDw68bJgSBhGxa0eH834Kwqq+LVvz8bNX
5Lre9bZbro+NoOQJuyKi7ilV9XezFozOpBMRDCrL99Yn1hbcicYC+TzKRTM/GIG2
TVhnQmd7KjuVsfc/pGazLUMY0zjp5jUoD8X9LmC4wPJjka4e/ilDJumXbk+b+Zjc
o+Kpg7Rq0051gW35h18wH6VMNCZv4+ljH5kPqG6OEWJv1zrukaaJZ5+bKJPCCySg
8qR/V2uAPN9LT1g3pBNthOI1c5TjfUpBkTRBwgEJU0EAEeafrmqzDCRlGZex5NfL
xAdFR2KU3OW0H3lbMgAdFu4tj0ZM0HEeoEKCzLOgzJ1ylRq1QTVWeH84qd8Hgalw
jnS9wYIhFVJPA4noNB64to/hM/vgDbrwXDWZFeOlGL61c++oSPxE90JDgNYcSxHN
necqln7p/OO1BSqTF2wxoNxKoDaDSWwgMfrcwktI3ItCwfYLcUxwUzNroOuOdJ0W
cSOqQoIXSgAa6OlHpMQl9ZN/dd009DY11bhGwJ9fbd7UVORnD81gnIEP+C9swvw4
WT9izGeANWEI0XXoXyuX9diJNsD4elEd6DqRsUs4P6Tn311AaNca2/0gcRFlCVIO
LB/pc+lEo7xxlJzJn7RaJH2Px9l2iHHAPDvQXv/U97IdFb8CQjdb6c1kHGAktJRk
OV1X14aQvflp2gtNdoiankyFaNjbKRIgXu6wEBOjO9GiwbRi2vmCO9YVW2rkj4/d
tsjMpF0OGWgJWRxYgNEqpMpmhkajZo25JdhYRnhV+YVg/F7Z9BZKZ3FwBAQYpmeJ
vU6wRAPEQoEvz7pALxkcvZQlKsqavrjbvVZQnAdHMtx8wuR2zf9HTtBNHgkelXV5
ielL4KBjoEC1dds8UW1zUtpnKrKsNtgxnpLESXxoxDjySjgBLsH55+iBVzY12RlZ
AJtFfSkqukMf9WB+HBXmpXXUFHVhARIL+yVvZcnUf1iW0YUoITpc+VJrfxcyrfUh
i7sDusReNDkClUdQW6yUvAhTdHN5/IN0FgQUQ227lnyAefCUrUv2n7H/Soo0BaPG
CdaMpzeX1E4MkfXL1Ouqt6TKvZPoifOA3CbZ/lCX88NQbKDYlj+o5FBkjQb9BHdC
N9JLh5ItnLg3FERru8JS3hR9hODC4JtyNXTcGlbQSOWVQojt/d81O7jaNwQkCM0y
K+dPgLIzzv+Q4MDT+2nVp3MGMwN4bn9kVrpAvwrtrOtbPfAJxX2MtxUy0hflNuzk
shTxTU95cIk9RIOdAPiUgpnn4EUiS9abSWe0hNGwlXyjiF67T/sc79JX+cnfGEn+
7O/yDdBXsiPxtHcpE6D6s7WqcgGpyA9BdzUuka8IdyjxagAzLH+fOXBZ247EUQ35
VzEfrsXb8jES8kCrEFyaXQvBom761hIYOcWdyk6RaLepgyjRTa+WySIfq4RWdq6C
b5WyI7KsVtpaiqBvoJ5d2FlHixUp3Lv3XVmivkIndTHfOgZGT1dd8l7JSB4dblkQ
HTqXepdZVJaEhS/bB0jnUwx568zmn7NEcME+g1juMt25+kXtCdhig4eqFwGDmH3P
Mni9o0L7T6gCb8Ird/kLKsBZeikno7+5AWChdq2yRDmVYYDAP5+II3esiXdU4cKm
UfDmvWs83Oq3CkLXvl+8jnr9rjSRr3DZGlJ7hRIl4uoP4RqXRQo5hElvj2U0aB+n
0Vt2gZ57kCQq6VJLKLV+cJE10qqlmuez6zAT3pRdNsN+geFcNBC++PLXSO/m7nu6
AroN3/rsEcyaZAW6BPVXT6mzgirC0e603u3OD0kBO4JD31nVgebb87FV9H8ekH9k
6hDZwYyRNu6IWXjUetQ598fAcMqF8GR7+4jr1UQzCFAASvtWWPJ9QqYK21iXWTke
q7DRJGx1DY+TrM5DkCbggX4sbBHgMUtYpttwMLQ4VDvcTwbWQy0lUlSrMZN15Nvk
986XLARNDeDmRyX6QoQ22Se2Np8lNMbNjlx6YL8nQXkAtY/Zz/Y4woJy6BxwkN2Y
a0V8lQykYHnaGcm70ueikD1LZYxEmV/sR0+mCqyH2GZlIqZvY/lP/uygGEK7XQgp
xXJ/85HLqXJPoZRVqJt3sswYTbhjo72IPCm4M5jtfYmsRPH+Q5etHc6KnIs9Axy5
dwlOkTJrY1W4yur1LTDBDq4qY3OUjNeuVhD1Rx0qobJFUrssovp/X3j8/pTDe2hy
5uasVHhelYDu5iNjzxfmv4vY6u9prB2B3uaArQ2ItBtSpluSw+6dEo94XO23tU66
goLsAAHVcxhXxmFlziZI4Ir9NWwcrFm1GUp4uFZ4FAGmld2g9V4u1yrvv4qcmbA5
r4cXaYW5V1d0FWwZZVImzL+UMyjOPi6SrLNYp+JTWvmVJXZ/5VTh/Q93XS0v6F5h
IlGXIWoiVHwvizmv5c8xeDR+4H5T57NvDZHq4LGcoBu/bXoHXSl/Lfekv4qVKZDX
AW1llMWLPGhltAe0Fm9BEuAM/6ebRTkA0cEltOqr8Bb23n9IMWYOKRzxG3HF+an4
Ub5W0u0tOVK42oxki5J8ChWVFb6FjeoV58HVBB/fxhGRvjmBHoI2SylPiHUIiQGl
RacXl/fRBz+gRYS+fypk4VlsvwsMLjHdgvY62yneP8BthXwsfgbEW+A3tauPMPMu
PQpwgVtLjHF1OFghTGwsN3LECD5Zh8sLIBFjWJAnt7WASLlXpO2yGALG4hEMMbsg
Vd8Nn5KOaVeojg2oavsbO5dkiAEyjN/aLyXoX77533t0J/lBc/qhsjaQki+NtEqY
x4D3p5Jhtl2ulmmSnfAj0qz7GG1xmSGrLVg+g3E1iCm5fPP5RGANCvrVp5hPwJAj
eW61Gzx9or/JPRDQH6uBmfdYUMs4mXPtGWFcKanG90THFp2DxULUKTLJYT3MZc+J
YgIumk7yZh4oRIz51XilQDYZQGdOPZHH/2U2OE7rbuPK4z/bBsqEoPsS39J7v/dc
DtGLs/MxgDF1Te3tUUz/hAqwFsGJc7VeQnV2buYPD2Fb+Ojax4lsLMeh6VK22Cea
WnWLACCFxz+4ix5ODm52ON75U2Jv9tOJl0hWR+A04nNhRK8AaHGI6+y6kTpt1Efc
fNFEiAq32ZT41NslDcRDNRJMrllcO1j9jDVxAkBsX21mpo7YGAwGywMWO/NSzrFt
s4JF7kE5cSSbIibY5XMRchdlUWJ78YEg1CfHZeMCZwlikcZprZYBFMx4iAA8bVPW
3N2Agr7g4xnNMtJ5UCbRX4mDsLSu/bm/xyD5DtZCDZR34s/TaGLyj2aN7b2pkCp0
3qtBDas8KefNzEFGecMsJvumQlB6++ktyNr0cCsKBhjMXIPt8DzVkSEYtRkGKXMD
vBOVIR4OUgpy6FU0O/Arti62IMB417A1HY/jFbyucC8249xiOZSGuCEwA4K419BE
kF55/2mawa3J21RZeVR0/bxA257Lt8dTMEMQHMqtZ8OdTGjrQNWdym+2AovEWU8l
O7pxn347/1RBIz8yzsxanrrZnlyEKkFNwhVMddsXYyRDPpgz761eNb07bwZzP4no
KfY5WRqlotkJ4++XuWqDu98on7+1ei9dS9KdCo0QaTZ3bRsoTJXWTergNB4ljzH9
+4RT0Nozd2GmcC8WohNfdXFdM4lOaUJWyYIdx3cKAnpufNX4WsXu32LOosLubChA
9g+GVba4jr1Dtg4yV24ZRsgvv2O2Sl0AMKZswBVsvdwt/ymKgzljwi7le3iw2SC4
CeANSN4RAdKZ6PdDbycU56lHgtxH4eThcAq0C9U1u/5L/uJ1cz1Oel56/y8HRsEu
DUFefPcmwr47Hn/XV0/nSav26fnC5D9muyxxJK1LxgBiN6WB0iK9qRcqmNGhaSH0
Pfvb8N1fM31fFsB0dgA5Udy7BJOzoY7hm2YgCM9sYZeD1sdpQ0MfAx0ljZpkw4My
9O9xz19Ryt23u1AinRJYpiEt/VMYgtn+y4ateFcDHHWTeJqGRDogvOvdSKarDrG2
AoOtzVc9e9meIOrZN2gRpoKJwoPWZWUlfFOY+3lAyYSrmz7+3rJIYHaY3J3RioBJ
4zzVkcSYx2+SPb0IfZbD63slcvh+UDUd7w9UwBCper8BKUTJwbRdFBEqpaf1kgty
wVfeR/+Ai89DTt4JjDsaV7ekYgNjd5c0k8/f2xPffLqN5s4dXDg4HycBUws8W5CK
W/PA3Jgl5qJnhBLmXGncxgnhUpFHDwMzuOVvxMxH8IXTKfRHeKQTOoZ0tnfNmC01
g1r02Y+bzL6jGTUOejlVuLoP94aB8PvLM0wD8zkSPX35i/F4My0P0MTNKRAoDzn2
waCmRSVa71wLjGLe4rTUSPZhtKJp1FXRcdQoTnjad7ux2SjbIiN+IbZ6Bl9JiaFI
z0QT+n7w3kmW1MZdJ1wg48EBWhTnQjC/YRuyGKlzL7JwaBAuatenZjJyZIDdZqHl
ZMdmnTrkAPQ1LKFmQGCjrZ78TipPD0tEW+OFCGL+aj9jRKCupElJ1+Zs48X9xsDC
c7YnLjfx5ih/a6CgQs5GVDUyjX7fREI5lz9JEF994L6hnDPqXjg5Akuap19J8Mac
C+ycyhmOzaOOwHiLr0R+BRD7q/L4IrP/EeMbzHSUBw4E3mPwN7qvVeDX5GMmbklH
3zZanD8Mg8lhdONBXxIIqY93qkVra7TsL6wqdtHFQ54rb6O1CJOWNWV9l4GhoHd5
Tpwhwj2fsRJFsmoCU9DLdxTDM1fkYuYBFu3uaEPxF1HBWVuDKyHkdG9LuO8JeOJ8
xXa7JBpYMMQsrFOdyu8jW4Wb/XcVlDV+3JrWNkjoJL+cdMG4f0XFW50mHhsBqc/k
J214J/05E7kWxPol8zyv5uO532e4xhVbPuSdDCmTHKkaIg+YxIUOQRDZJamWc1pE
Srqp1vQ97d0ybUvWCDEH9L2e2QIr3YNQIzF4ZevVUJyu9XNLLmUCQThFTfaWy0Wx
nXt9AKUXchOQcZcOT5duyWPNS72a13Yl832CcYeQLXjaONg5JjVyZeHV+9wfJDGI
OeN+KIWU9qOdkBSxGeel7/wU+M4D9LSOYboUYXDauSrlCLiW3uR5EpLJbyAO6pzW
RmPPoP1CpoHUXa5No0X7OXkHZ7VSdyaWFUQZCbvt3urAm8gf49zylKTnB4FzHgHi
wf0w8/mVY1Dx3573XuTwGO2wH2/zT2yoVwccJOW1eXxC/n7XSdctWmNTpDKZj2wd
5ZofHPM3+LE0h53/tyHr4kuk9Pp2RfJ8lx8TyLg3pPMvoYa8Ll/U2LaiG3fHFI0W
ZgwJu7fvsuIihcNtCtukAiMPHKNbb4LAKFq94Atcrf0cKHecaobW7sMmefOMkoim
2XX7120ouIiYxy0AzhCFni6rWyTTi1bql+hV2w5206Lj4mCoxvlGnSZjimcH6+fX
uozYoT2pqsX2DK7xIK8MiqzyFYXWs34PWgbxzxno5sixrtoRuEfJEDLWM5wNOa4f
Csj/DwopApxKRXIkOa1HWHcXWmk9e/HqtR7AqlcnUYPy44k9rszxymVUhRHFZcp3
cEuqCaVLDVCLowN4Nt30r+/hZjIpD5LwxZvEIG/uhqPuVxFlI6Xxy91LvNTlIQ2l
b2if4qukdj5hvS7kiTwju2x2Bgw35d7X6hjepfiJUbSX7oVdEXvsWsGUlVuKHzla
6vnGSfRVhyQSaO3Xk+i2dFgGSfGJj2wejtSLQ6PMwCohEGN/4k6tWQKWDHTRznGj
+hakG4Sgf7rfcWdRQM0tCzkB/zw6j3DQKd57bLnj4vRRA1bVukVor1AhoYC0F45P
cODjXpRjubFeD1coI4quKpKXJjGb5meKBacgyBHkFdiMrIpCcuVAuKHBD5J8Ue54
IZxqEUKKhMoLVaEO+zZLjTPNl6sze+PaAhZ2kyHPLdg/r78C8L0kvSL8sq4CR3KJ
jyEAPCnpZaMh8M0s6XkQ2mcOK0x38NFgwxKeWH/u02vT24EUraFlSaZwcnrZ84en
h4yIHjp1TpbKdnnYC+zm3Bw1kl1Cs40Kk/eNJNpu24AZLHKb++4XEUhK9dgKpe39
uK87gNE9Z1p4sq/c7V2PgF3DYR9+/rm2wZXzB7gXNuUfVZ2DZsJyQshUgVY+JIJh
qreUkJUDZIbVQYufdzrmhHcVBJFbv/gFW6cepzs7uOsZ/qw6cT+Pr3MS5zNp7Fuo
D72WW+Rx7BhN/U8lhF8xQ9dZ90erN2GkuYGHotmXSCvkpku2BUk29IuC5VE1lihi
F7EzCjbc896IGYvVbtxFlu5fB6DaTN272ZpujA5FlyO7fIDdK+CHdkQFlm9TZR9a
GKo57aY71Bdr9veqizpC5sIZqnd1ynPk3qkx0xa1Lh6bnwHG+c9tFERRsAoPFAiX
lzBzV9jX5ItZiQU+52acxC3XEeYePHy9flsy3fHgiFe86qS0Muv07RRZ3x7rYMGN
9oQoBriEl4CY+gjw9X74oz+BdklzLAmXdvd0SWQN1M/3nEaTUZ5yUqIMY+bDZC0W
xb+j4gIw9AktAvIxbkhmckeD8GqoIVX6Qo5ItO5InMr4kcSt/idvv2KibaI9/BQB
Epyxzrw2/hxxmL+soZChPk+3qb6qrprybqTN0SfEG51StuMonc0h6O/pVXwQ2/t+
lMnMBKyxNLtbTgZTCOOseCpsqmt5DAOkr2FTf/emFoGwObEDAtlwE7aNeQl/s6Ey
yZWm6djq2hIKpRRB6NCyIPUrFXJLq3+c+IOVVrkDLatHmkQBDdHjMV7yl9ctiAXz
quoDUgOb9LJhb8QaO/Z1++ELlQznHrynrrG5ziThwN7BgNc5UvG98WtRnC/GU9H1
GUlftuJBkBTATYxsUelwKxZA3ef3S3MSwGNMmTV5TNjq2zVQgQBwBMTB7zQPghdg
1azDB+QLqy9S7OTmJ4kK1L0fGL4E//H2OnpoB6M2KYery9xuFndKXUa/pZaYnFAp
O1MeiCvc9YWq8/ZQyO521aOIEvDTJlZaZU5SDFR0y0BbGlgdTuqVrqjR/4CeoXjY
HJI9k0fM82ZynH9E0oOpkaTJPCfcEStzRVVFJJHYEAuvO0NAaYDnpaWi7l5fQ3uG
QojQ8kdN8jI7bKh6fy2pSU350CmsYDFZg7c9GkFVw/BccqB941Ix77WlH80CO89o
lxfRmbM47gNTiQPETOIkH0y0emJ/aZzzT+m5ITTRdFPE32lNxYl5O2WsfCAKdaAC
QrIdiYpgxmTwBTfpVaOcvcQkNgFOORoVbgRazNis3Usk0KakrBBtsWNqCSZIbXqS
ng/ShTbz+GUcomYOal5mHsDr3FNLpQM8HUq9IzbiS+Ck+23qvnIBg+Tf5I8RHG+8
ToR9XsM5VAUHK3Cyhv2Ymnvi/Z+jjoQTgzro/bJL3aMsX7PLUISxOo5QuIIhjHcW
XS+O2lM/tITzvl21LelH+hj3KcnWWxa8gNi5zs56d2HDUnw/iWix6u+8NUHMOq8d
WLeKlIn3j+I/3C+2GpwWXAfiIzUsGRtvkjhnwq1mH8X562ACy58850jwLoo+Ndcf
0LUiiTXN6BpgUSIYVRSq3dtvCpxkPiCBy8QQVCq3G4qApTwaAHVo1Nq78mWwCmO5
QxbCiafst5u4eFXf4cy/3OlismszI6iWNhGlMSNCyVx/7ypKnXjngBiinHCM2d6O
bUllSrI3/u8+JH/BQZYJQGIRl8uCsvjWRB+LldYi4t0U1A6/WVPXTXkbHJkpbakx
mqhJWNAzj6NJkCrPYxNFv+9uQFG5nOgxHfBHSG6/qSzP3KqXx7wZqgEoJRdiVCdX
fDx6yjCG+wihVmyYCGqJVJCV3GXhBhAHEs2G1rJQgEnWWVwDE/mElXb0WRcBVIie
8q/lBeL9EeoSaz5NeHI1NZooTEFw5Rpo864WFxO6VV/+g2j+Ig7Rsd4oMLay69bM
JU8gw4TL99sSZDiENMY/UcgPhE/BtTdXEaob8AHqxd7FxCvzL4kuKOx+rqFTB+qw
ZetUguuGUfBmepwVAX3aE0NwZjm7yNk3fq8GgY+oeUJgFFFzXZGDm8WS4ArZUvDK
ZYU7ImA8Y7G6O/xkomTVHvVBsN6ExMpdORhdXR31fTOphgp65IQtVbt/PDourbZd
PXNsH/H4tpEtwcnLotDGgLJei+gRQljC0LWglN0qgRE4qqzL/3Zfn4a2NNvKvlT/
HMdVEc5evGOeTx8X9jq6nbCot9dd6cKT775oYjH5vw6AsCbVsPtGeDIGBrQERFu9
3dKCGlCqVj9ZQVmoDJVwqnHLVUYdGgrlJdKbKDQDa+bUfX8+dnxLWWKMQH5NFeDW
XZgqK9Lg3TO1OwBRb/ZT7cMnq/fk1FgNQ6EiOM9otteM+jQTdgMmlVnPGxJYAz2X
K/nwPCe2/Zl/79g81YfGsNN3E9Cdkkav0VFxUJz6RRkiqEXimOTxFMr13TwYluXi
7dL6wwXo9+cSuKVAfIowB+9im//gbIghZmfBrbMHgKNzOxXJhAlqxt9Kyhouhdyp
fVdIUAW+x35wUtYz5hT241rS2VlLmLhEVpRcy22wmabWCIKJHJEwKu4dSylCnImJ
Ij27phKca0BLKb0um9bHQj3RRC6MEDbX/MB2r88fUFdjN1N8FOJMACZ3RAPuwKf8
A0cD+EILCMBARPq0QPe472xs1ZuL6D3OpzG9h2rDWeK8GcyUJcQBZ0ZPItYnGvWn
ikuG6qDsPCNGRjallKGhKTKsWlc4NawZoXTUXaZsGfD/F6Kxp490nog9eW/H4VB7
vP17x6Vh3JMocpEtQhfkD5BZpBOE4ZX5HRPpsnWHGMZ21lfibENoO4Ti1Dx5QAf/
DewuY5p1ewIOy4d+7DrFphgWeq0OdAyGfwV4QFmhQgrPATGG7UK3h6kfkkOOtQht
Qj1mv9R556U/d11ZE6NQLvMzgJIjnpbcRfBFvMl0/s3ucbG5tPvffBlM2Fe4UJEE
hF8dR7ozWfL4+GGKRe9nulN4RiL5XaSPtBb9GK9tBcQn4mJvnyI0fXCmW8r/snlF
KRca++cSwPGOtxAU9xQB26UxrJU8TnJU8fyfP1xIzvDk66rgykUN0sdL1bBsRpPq
5s0fhq4p6IG6wxBYiRUA7XNvj43ggrq5csR+7dbzATSclYQ/fOpkdsBWviPRqCkx
J54uHnF7drnI0m2t4OrclUtOjTrvZYTiGa1YzRW/OzWdEpkLKhfPYc5sfV2uyL54
8MO/DzwT+UoWmLMwolHKO0pBH0YpyuXx/kTay0lna0+7CNrk1IUWud96ZQiZ+YZ2
++yDw4Jph3pV1Up22rMioURxsKMgGb4Z7vGD/TaH+IcJxd16wvJWgNqX6CltdCfs
buefcynJKh3ExmUHn5hVMZI52TrxjTAA1I8zQs0yUOJWiyoZcifnJR9Ar9MQD9yT
BRKJWIEHQ90eCVJvLNCEML/JTghSRwuYbnfEsu59m0PUMALNVgEnapW17f2XyhN1
ZGMfv+TAubX4lcQ6sRAmVjM8PFfkLbJ/Ra0MEWURbUkgSPcWkBLEED0TgG9/IG8+
JCjhaoysOFhTRxKkxvfm+Waz6RZcXkAqqC/Xwvl2AEGI5wwIaZK5vrSNMzAe6I/S
MG9hT0VzOVTAg+nKCuubUG7IsAJLE+tcPEM22rAz9tfkYJTrHTG6RMtCGQ60+MHu
+VMqGF2EIrUxJBJaIB5t03TrCdNFHA1expo+YuqKPqLe8+WlX5Fca/KwkyQNGNO/
LJP7DBjpkFsmYEh0V2IAyxtEo+WI41tZ+RNBZ9udkx0Wv3S+JMOYJbevyPdGZf3e
04DfcR0wqAvXClN2HGHzjgGM/1439GgEXiuNodD3a4bktF84+yqz9zFNJkv7lkbu
Ak4nkxFV9DYRPaUihxq+nrqMm992oWH8/+0JaKGcHuLFKoRR+D3kCjAO6AWNKMP+
p4SwLAO1QxocqzB57f2SkEVBG8/rI0Lp5gnIgcNZhYBuP5uJueSlOq5BVLMBWU18
XLtcqKy5gLh6ePzSV1jgLYGWs5oImtyGSYBiLFyp1y5ETX0mpF/D9Sa6zJxtC39R
ndHW26SWuWQmj4Bw/wx5Du8tfCmL5jZrJRXnJV6j88iKadJ05gDDGfUgdUpwzJL8
0xcuyOgMxBASejrgasQtpdfakWUykE7pp6BS8CVT2Ic786B2q44YnXrUb5RahNWo
khcnnbky6ejT80JWMVmwWuIUt9EoeBWt+yvc4MNB3380LIniRkSSrrBK4h0jNddV
MLGNKrdQWWl+10RbVCeIYVb/OL/DMh5AGv4B0rSMVdoUAkB0GyPrBFRLVl8FKmOz
Y7GDA4spxpmA6kVFPq6aTBQbJPNV7MQ+xdkCXY5cba/rHBqaaHIDS5O0VoTwS0nh
09slUAUD62SIrBIYKsSanhAPV7Z5yU/WPXgUXR39saXGT6thZYoUME0fdeAuOZia
0bkbodzYEWC0fvNxlty1bzWixepyIyZ/DEUMrYsLBzpguJoF9Ecjc8hugZcUgBHd
kI+r073YFRnR+8aJ3DaxJFTvzdc/ewRsEXK8b/dxnwuPEG/LCfh7Q0S3fmU9wzAo
ap+MX8pj8EmHdXjAzDLr+MM4FDDN98Gf9qrblWd8/vFL4abngxrTXQvsI+nqkSO6
MdmeaxSGPYiMFudyz5QNcbH+NcYHeSzS7d8b7UdCwO2KFYzB8u8UBZmeRrmnURi0
9rBdanqhPVzhEKlicf9r7LDvWGAWAUd/zA5R7NvzTVNBkHYp4Pt5GKeGlg+ZrMfz
nfnjzDdLRhjE+7iZqDEykQ6DpFQ9wTxqnHKdcQui743eL+RjLhcR1Jq+wbDFOu+F
kZqh2yWK/qneyIbuNk77QE4QHz0MiIc6PlYCOFCB9Z93QqP2xjB7QJnwR7d2JYxZ
Z2LUslCOChFOZdxxoYoyG11Wrq2jUaNr/2Uc8FRChJiB/CxOQ5HxBUrIIF/H2VGJ
8AJhBSl/CsPo3z8uNX6ybACnazeKxRMlYMZ7MEm/3PHZGCjdODCJdYaM0npUJFrJ
FFq6r19iI4OkbuQjrotIikvPJo+/U2F8XFKWp1PUOC4UkLQRXr/sq+WnpO1ptanv
/i3FM+PcaAJ+zR3rYQfu+eeRkTUpfxPIiMoRIZiVCQ6rtiinL4OEYE75KTokxWtm
GlAL4rjnoIHSLv+/e8jl9mxocH3j2HmswcbZKecbPPAZY5ZK/NvYZCbuWDV8u/sd
J3c1tAivM0fuCgfrmPgNJIVBtzlElJmLuTudk8ygXcP3yDs6HKriBXKUe2iwDPt7
6v2FUR3xXv7RHcSoiI+puNsc7PpAhRr9XD64IaDRndGrSMjT+84tvhmw/IHxYeTN
a1JG6xd2s3wvXLScKwi/EEyMV774rzISY/Pg9rr2cPQCX59So8YxtqDJecZOhsD5
DZcmLzqSmi6Mh/ReSpYfyNbsKdCFfp3HJVZY391k/3rKJFojIuS0zr1Oo2LIYybW
PVSUrjhZE437blwI5taH/bN2tmRFUCkpo6x9cS7ciNC+uR33K/Yny/cf9MiV+Aek
ey2OJEC35FXvLUaHSZbftThEVG4Xb51P6tkev9R+xSbHIY6vJbBtVXBeQkAFHJd1
KI5Pwg4EEKaPOIdAgwSUsIpQXOTle50tko4vrC3Op1oLME06m1RBeyzoTnqIw2ax
dQssEr8oR/mnANpb+HVCSd/VK/ovbjevFehP08CZ5TkUZJNw04Nn2b7mCOlwSJa7
VXerWRY6uYA1V4XLpEnvNE7KibJxvyL9WQFOvZbYcz5k04uvL68hzLk2v3KnRMjc
4oIiGTqLM9Cy2iR3LVwpg2zjFhT2YkE0LmRDq/MVs18YkOXjoSYrQIctRXE6DUuF
Ly8tELnxqL6CqRx1LchK/osyod1fbIWHyxxLuZNQ3D8jDJwCYoQdw20+5wQwyK5N
FiShSfiIS66AQj5xoAkADufsNw15CY9FsVqcCXsjpLKRR/VfKNklpoBwemkM9gE/
+WZexnV4ISTlXQ/3HKOCug1Yle4dGZI/Wb0wdk8nrlYG9ITBHmCrv06AQc8flJtj
EnPslRl8UVH+gFLsGcQlSd9aAgWrqidNyFhE8Ugs/+zaIaw+8QDKkhnLTRRu0+rL
FYPzRNxpbYKrTCjAqSzGDKtBzkmdSyX4F2nKst02yVSDJwF2hxu2FnT9NkzzlthE
hqpAFe5VQIrxuERXUcozNSiWIjNSaW4j4tSerDHhLEtVk/9Cf2KjiZ/DtnUewzM3
cf59ahlP9W4I1ePhHqi+LrfJH67QRqJYgFfTkYn4r7/eczwiyi4RwFuuGmPHOAXc
lxwhPhrvrj+BeB1nyDs1XHnR7BNfWNss25KjZE76j7tvMJt79xQBCMqGS3KrxbHH
q/1X7+xrlE9Y0sR9KoVo5B9tgeSO4nYRnlKtW4fCNi7tJynkvmVg3UofHWgYAyxU
uSifUqzViufxami1axI30/L0MHruAgvJAf+RmcjSsZrWHzbkuV1Burzi1X6r7ZI4
u0ux098rxE3VbkDdsqOTt2fdpBFcgt/3T//eryImI1h9QlTBUkhg6u+l/fjGPSiO
8rf60nFxyYIXFA0IgL+khG1IvXDD4jSBneBJUKgVoKBa1MuGWHXTC+n3VMV1TeiF
jVxv1t4tjhrDT0njY0/sbZsVBAnmv4fPMIvhA56e3f5Q7YdaTd/l/7Z6MR6RGsXw
h+YtOFTm1SzP3v3fRvyUYem1pAXy5oAYLfyQNep5QD7Fbt7wF5FzK049DCDyU6MU
ixBclLaUpQ7VJnXNLmZKUoOZ65zYOPYyTwgeg5+gtrxL0MCG8dz5v/MIoLQp9ak+
anCjvfSJTC2Hjmf98trAASuaJmI2P1uq12QHUaee9I3CbgkIGcxXZTXgplOmtMPO
LgcIZH8X1hDmJwl+WdH4aEQRo3tumD9PTmj3lDyg2eBIKxQnTtQS1tsfCRJYw+kT
By2EWRrRiiF1TCQwquO8p6Ve2zzFvJyybMCAe2fNwhk6GwOM5PzWgAV2PSPGzYAw
19iw/Iejs1B0KCFime9qZpgZi9sshdjzjJ9nbrOHNOrtQcWJJfq2j53maktfTGrD
/WggR2aQA9B/KADRwePtccriWYTmGUYjiBHwfZMzsJreyVpA3AeqS/qKlAUFxl20
5xyQJaKobHu2U2DUP046xwwmPut2Crs+3y4Ue5D8X8+MDkzXsbu7R++KEm2Ti6c7
2chTVUa+e025KZmGXJUY/E6fWUDY+uWxN2OKkhx5fZ/XgQUfXgcb+aWCuJam65vY
wMHNvM60R++1ZDe3BSceUSMKCz/aXXeJv2s/0+SSvlAilMzubEKiO1stZeut8gcg
fhPFEDK08h4SaESSQ9ZXPRt6hXXhX7fi4J3hpCRIfdeEc6Qmz+ojqsguYl/htDsp
uwrtSATaBYn983aTzOK4FRzaPNXTX9gcr22ZiB/IIghQ7k8N+Y5lCedfRQcVWAlt
6Enm1baUmjgCbQfVYsUspwahxspk0njrc4bd/sYhpf9r36IG4dlfyGD4Xk1a99Nn
jCgKP51HFO1ZK6xF93yhG2rM5375TmfT/WDUl5k0thhxbZxhnvEvxltnIezGcKc+
EYb2YL6sX+PWOA7iKM/d29R6O7yAw74Dl+hDugBk0ApzB+GazPIwi7QNIHXxLP1r
9pYuRaMQGbg2Hebsx/WksBdqGLRImUatUk9GTGwINSOC9QLTuVaDdrYk9yvQg+Rr
DpiwIfpFrfR5X2GP4hc1JWtGOoCYmg4bEz2fsBWBd4ZyZsHcg2k7ydFiL2NvAQzu
BaL4LwHv2FCwEgLoHRAGGb86XLDh5dG7tpTin4si57E1enobUUU3sqRLiIAV50sV
Rb683B0y1dai1yScCL0aEte9S/HbSH8JWHeMJvEdr6PYSs7cpSm6BJ0XL/bcmCmQ
FD+l7ZCb03ViTmj428fP9Y0A0MY6y1I1blOb59Hgx3RI8qWdwxKPV7NITAjmoJJL
VkHuWDSoldPWD6+SyKOA0uU44Yv5r5RlWod3t4mu/af9Jwv1T2qUkRdD7hBNxG3S
4Jw1iEVr3XMFyA9YMnVvlOAmJbkcxShQjZVB9+6t+M4967S+JdcKFaRuANPZnWqp
38rVW0BKX+P9SDfniizGOBY4fGVdm44kTplTZxd7dS0PZffOWoeqDt2JaqeB9kLO
DuBpgr2WdxWdLZk3NYplI3O8xenxsYZPvoY8UBRm6AJNezwaGDwS6A0vUBOShHev
+NoLuqisHatbC/Qg3dXHZGUgM7Qo8JxnyQhSUahzCIPddiWtpUF3+5o5UrS5cH9C
/tvfyLKOFsRGbmNDIclEPldBSVrxr6jHWRi98qECxkbq1i7COhASLMuzTRs14Nvt
ybb/ML2qJVfMhYdB+ngbtr1SvuqSKSoIpa3HUzIwYO/dkHPxIXna5+fxpHUKUlVm
dMFlnZJkrHwczCyFpqYB4cW6aKih4AXPxBDzDg6qJm7PZGxnWogQ3A3mBkITlEL/
Oqg47D1hp4Dm09rDXYK6YbVVlCCDrlQQk47KZjkXhSk6d3pTiCnnOX7PrvOXzdrb
g6zbUEFA9SBKCXxLuB6mwS7HHj6BytmgReCrHtsPKCPS9gvDPyWI3hMLgp4A0cri
PhONpoDpyIaCS8UWIRpAMcY+mvljlkYkQ/CMniQPm1zD67FTaS2zKjOCt6D8DpNK
e5O/WIaxmFa73x+1Q6hnIadBGCQwDlmUNgcv6ghM8qROzRwUHAmQc167zD5km7lo
ncROc0cItvtIXYfxPRtupnozM8Na/NjTer2woPts4M8HZlqEPloDHw8zpmePFa9S
8Ot+OkG/mT81HeI7XKmV+9mQLyqN/8B7tyjj71SpubTbl4X/qkga07XjhykmPPjt
x5sbZPt9od/6GOlNI7OPLCsUy8eOm1DzxV8C1ZrwV2RBcIrfgXpZEbsbt3eiOUhf
bPnQzxsqd5jFM4pWY5JrNP9ypXB5veZT9ocwXRJoo4z+yV4r0I0lDQpNKA7b0F/1
aIo3ue0wiZfsw1Ndb0+cT21/IvtjSJSaDQsRZRcA+STuKcBnVZwhAafh0iUUxAeC
DthXVTi0TPSROOyiAuSWxjJOTijCn+pHqSf5IIqjwif7QaAkPzPTJi1+l59bb59A
HJ1XqbOi05YUkYSZL8WbbzUcmfhoNzdYypKRWoaAm+cHyegE1RgiMvP2f7moT32F
5zRd6L+u+3FPZje26iCrQj6ApNi5G9WHUsu1rojkI+Rx+aEIbfwNwb88zNFReqoR
hI9HUU7I6C+SmYwvNyY+AEvTWB9DPMS0oAKp+vVPogVwKs4In+5qCsv5pJG9SAut
Smxw99hzmx3LHCcQgXqeX5zmcOefvuTyn/hqkWFr0JgHI/GU1XBvnqmIvLC/dCeQ
Stj8CX3L92HYkigqZK7g500I23bUikmWq0jvYi9buYLvm2fJjDxE+M2+25lqnvNH
c5/2rVCuGV4S/1f+G9WrFTSc0Ou7tyDHR1TP6k1oQ0DpYu/nrAQJ3k/3p2PIhmRG
hR7WAvnuvvwgvQ9b+EtLYT7frACbJsZgovpHY9jH2O+X0TRESsi6NmxAvXpU0wmn
t0XMadoBytQ552sUApDE7zEXxHNXTU3w0gcfw4274nW2wG/Pyu6ahXgf6Aqm0Y1j
haxIi3zNwffWwyMF6wEqBmP2v1VczVdNSQhkGi44fjyXRTR7uOV+X5/LWSh+eRi6
G4TxFmilfcJHuoE+ht2gZZmF7xrEVCQ/qOQm2toz/WyCCtHBuBxBYhMCzBmS9qBt
ytFdmGU+5iCUkxCWvY4aUvNwurEqSfZXVUMKPRzv7SX5L9zjl5dj7EaCkS8uWCSl
Huq0IDvULdC3pzeoR19x98lm9jr0JnAKOGcgr3+lJLdnXfPPUSSr9pcuqnm2ioaD
AbjTM7sWWiNtYQviK75SCYq6hJ+1lU5qWN787uXUzeI9hC2chm03Mh89k68KspCv
jfefnw+g8HH4Dq2X11eo4GxuoY8MfP8jRtBy9XclbXgzIbCGF2xhN4+h/PZsRrE8
yrCVOU+eOox8W70XRV7ISM+CNO2bPBjoykzCfMHRxPd0L2nLtA8op0JWIcW4q9G6
YPINGiVGyFOH6dwfr7ga5QikPCk1uuAaKOdUfZbGJLcDx1PD04JEAEByK6p4WVRP
qOeBL/BL+bDIv9rQFnUrUWEybwStVUbAvrYF1GdmeHTKv+Ueb6Jf2YJRNUSgwLCu
GlFQqlJiDuAv9/ucZe/U2chCKReD6cIsIBa+GLnGexweGSjvcDpWsNLUO8GvmHJf
1uxJhWab4trg/CO7ogoX0lDjpNTZ59F+GP8M/Lcd2BlqZuUZiZ/CbXhOxUXUmd78
FSalicEmAFAEaNRyne67wuHjpdpdCrEmmEQu9ZxZ7S3kUU0MKDJyk+DIBeHdYzLx
UxWWM/RKuMwUoxX2tMx6tRJf+YH0g0q+gHO0dr39RNQNHO+LAFA+v6NWKTDyM6Br
nrII6HECtTcSAKF8sxKtGpdBMjDpCTXofYiLwfRJZyyrZZ/o4Sdy1bd4yl/xL7M0
OIprEfbFpEZbpUKHq2H4sxZxNtOgRo4ExgHD3iJk8i5tBVfAw/DnTnJAVqOTboOF
YOncg2HIHZ+bniILxBK3HhQlk5oODe12Ll1SzNzROD3ORSkVV5LGELG8nwuTIdIV
Tij0t30e1wGj8qXPEUghJsmrLou+aGE39Wta1I8f5PbxIjCjJB4yMu0/pQEwyUdA
vVt9OoBkfKOLwWFdwINOF9SZQXJR2xHFC8DCoxuJ+xmSXpt2JZMvUiB6pJJAYsnL
S+OiGEbdtXokkXbGr5Sl7sFDRqaNlOSTk+5cZ7FB2TOdHqQP3SgLk+f88J7CAoKI
RWTpgtD9fRA8Io1WdQn8E95rZcwljwrPr+XFxK3FvExPEY/YE8AUnSWIZYmVENtF
GyFE3p+H7KDrXtT3jDDr+FBRrDaR1ixYVt8QkxqejancTTTEsoyPWzgH362ypIUs
dd2cLocDN0iDqAqn5vPuwhIHeE7dgYRbJ2Y4jYNXd2MvJi/LAy1v7ErDK1Z2riFT
VTsqV9vayB3DqwlKtchp9tZBC64DUsCrIhnO+etCmNC7D7P04Q9rdREKVuyqMZRK
n9kcncIHD2Ipsa+cKLJCbeU/sANMr716Ip8x91e07FV0msxEDobNKNfYV4qRd/Mw
UFRqffEBeID3PqgO8MEyjw7Mw71ObqiP7FyS0rEkcLnSKu92qgQlv/GB7fIuKomy
Jt8Lt1DkWF0/tGAcgC5GYinjb1U1L3RDU611hJvM3nV5QVZMDbWivE0oZSGPk+iO
lvxSDPaKwhrThhVZMUOsKvRxP8TO/MnS6PejlXeLywrqgXZa8bRug1tpbb58c0ok
4hwBBAh45NUev8iP+w0hzMQ3rZPqZqvuh48OoEOHw3LmoqYTP5IBYzrNlPr2UTUF
WbjmrOi/1frItvlnVhWObi2+ZgkQ1tLaTHK2IMF0Bb/iEqDdeiUMnfdYHrJjko7E
xkbg2BXWgJ9Ugl9Nl3S5/n9xpYwK3kBdrWNhZRjYIFji5Ey+7F67h2cbx4r0j799
+Wm/TnqV3rehYK5Elc4B++/CV7TX10hStGxbkWbqwBioMLrkHJ47hCaGqZrK4fCP
EYzCZvqMEM88hgczHvk/BNPqI4iE7+Aqu6KyYHV/0h2N1QpAwGWJunkBCRgpitcg
XZFYdiEVLYqa5jpZ+wY6AaTtVgaam6R4dMN/zlksbE/pEch1iQJltX3hSHLggV4H
HFwio1K7gsYUrIKSX7eFTVROUF3YhM7zY7LGyIz++XxGso3q7maPnYc4SNdEBxbS
QcLZoOCwL+h9rP+CCp9233tp/fcLivyeLEXW7Uqjnq5xnqQKRwLLBLvT6nKI2Usd
mym4O4WsuRtCao2vamsn2ttzCORFkG9GVIHioRcI/Sk+V8XQyF0LsVV3+DQwdfGu
RDjjODKSRQCvBuy70WnX0w6iV7T+tqUyqju3pYRd/rEgCeSoKpWWWuzo1L6dWbO6
vOUc6qR2FwaPVfaoQ0hlbfbhA980Bh1D3p0Avq4Ua/iqKpvE8Pxg1qSi/OESn/b8
w9umq2XEAwFNdPbnk3WEKrcyuozj/aOYYVbr8EA2T8dFLBT0q8DSHGxkTQ9sAyFJ
FDZ7Z6Yr/AovgDLxLKuOqeZcJST2OErpNUAWzNZIr5y2Sg3YJRVHqgzP/V3vEqGe
VzYlrSiFuvlpD7PCGaeDhsuMWPWnSCT6PsEIQ52JwhZFID3I49XQfzNFNT+p8i6H
Jhx6A5P8k/B5kudVB9RI6nCtSijqiqGefPdS5o35+YVgomZK0sh2Fw2dNniIMI+9
hOdmEZlgbGqza00M3EljwqFKarqKFrfQst/u3wJVD15MG+j0KgrhU5GLr6tFpYJ/
F/tBCPV723/S3ejVMNbc8GxZECmjxSYxzmKP0B7chhaw+YoGBdYwL3d1jNyB+Hdh
wt2hPgZItT+3uoWNO6Ef/if6YHlkqacIDQRZSIUqmnRNYIHtPxcfTe6cuHHpBFsO
Qu2nxlr6VpDmsSjhNAC+MkY5cS8mziwUYhwxuK5nxp58B7oJ2WXY5jmXrAyoG8RJ
bJL6pUCBBuD38UsqfA924iU4k+K8GClPBZRMjpH6ztizRSalQvTWtHpnNaEHWQzD
YYMB7sdA+SunOIOeH5LXjJ9uAmnvj5bArbwB3JegvUn8NRLqlf4aeQ6t9wMWt5W5
5MPqrVct6DScl/6iFzGW3z5pxitFKgQw3ZtG+tvIyOprgAWOrTovMy5DjjFudkJs
gR9YXNe+lPyLrZNgb9zUU152F60MUrVd01yWzF8zgk+JsHsv+93ZastMqbunV0m6
b/nBaYy0+LxeE/Pb9rIgy7A3HoKjzOjtNl2Bwp0uIeTCrZdqh5nrlx2FSQlm26hc
/kiPa5CGJC8uDEbU8mvwB8PZuBctowux5JBhek7cK6ZhFwtu6LDFgdprm44G6gmj
DyQuMu57hQng2uqge4/JgCDMDg/W1PHNAsecVbZmXOFMaKUyd/KKVA/7LySmz4Ft
E2YCn3FETsU2vGBUbB7PaNRyw0/KFKwE+wJpcYX2W26fQw5lv46XNV3y/otjdFNp
pxy3pKiGi5JjUnI584O3ubiZe8z/7x4K91UtbiaMhmtAmqe7muDDs7XybtUUaah1
ZLxnzRcTAOV4f81biCN+BRfLpaqF6dKrXzIndkpShWZUgPRx/nS9NKRelulXzMSD
yB78VkUwRX4n+Qyb3FpXvshym5vKN1Gi440GF7aLnxfYkzxmRMQRcGaPN8ce2MBp
YGv/Mva/skN36Y/4i8Amv8l85LT44K4AYKKLcF3UVXnauKXPvYDgB+fAzDPM+ZWl
kG4hT9tWOIryw1/FGSjm4abwbJvxNg11756l89ViTI7EeNvhHx27wplAtL9MKjj2
LL87TS/lN3rOIqv6WhyO5nwNuzGlUyznWJVtnul6D7vA+4fpbFCRIg9PlNoy6yU3
DZ3Txz0XMCj4GvPNLX0p+aCegfUbSZFw1jG8uTPowEfG4DDfyR7rQqn9TrLgNhE4
F4vbCTJ+jMwvokPbrIXS/MQKcpChvz/oapHkf8d56bLHsP4pLTvbElAHb3z0fYK8
Y2lPTmdrVkPKrBvDU8kWsDKGa9j0LHd2VTvhOHlz2TbeXRXxKoLSjxywiToKu7Cj
NsI55TPk7JFgCImRXujTrfNE25Ehl+B6PEpo22Nj5z9KdWBHvUC0l8yxqwAWVDkL
VypYvjHPaXeiTfF5/CsOWNLoQ/YWtAaKfAUR8ER5hgTIMs/VhNg6GMnYwN6tnvaE
0cCMfbokoo3iIal4BCdrBTpUKTzCh1BFPLkkx3OOJ68Ha6bcNvl11HOT2/Sy5WDX
BN0lo6HXqR88tc/sabARtCCmLESC+C3rOUjPznCG6JhHG2CRU19lqYl5UyQMAv5r
gNDL39/nwe9WmtM43RnOYCxO++7wd1BnoUbyksTu2nWe9HFu2tll2ccBa25b92p6
O/2QaG8HfejS4J+++VzPhVL0ARcksX0vYGyyneskzcdA2nuszfpqV7ubYgbIx/ED
qY9e9jhSDCPFm/d+Fe0qy63OD4q55WB7MnEphdf1Gzzl46bJnstcVDkjl0Qk+9Do
d8EjleTYK9QfscU9YN3NwpfoX7aH1OHwleimH67O9CWDxzPcX+/o51V22TRJxZrq
6zqP9N5w0fLTg1WvSBKsfzPf7pWPvW5R+wUI8RaEMROM41rUxlFIZuIo62iHGhE1
fancVathc/YQA3qTQ0wCtt/q+ppkaoO1D/GYJJRczWzaNflD5FmGKPfKKt+wimak
tBFy9/1lJ53EjdoRD+ii8M8K6uZl1dEcke8gZKN+3r5ms1/VV+UxCTczX8gza2Pt
JYUJ41H1KUoF5L3JgMPz0a9IsEiGDjI14RXJk/MD2c/OeQ4oyAvZ5MeYWioxAOmu
v0lz+Uks3Ohl0YEM3a25Sh79o9w9tVcdlLE6+z1aGZCb6ydSw/q+nCZxXtfhYSQb
UHOXnnp1R2aKBekgSIDeO1MR4GzKvRv2wTy9wQmUHt2llGfDdqCAZB2SkOEueSeG
NdwMOD2x6i21w4Acjh5EG00kSXHr39sUUM3H3FnkPQx9R/4ios2sSPzyjfGWVmMD
cze56Pnb0sziBx/wKPhWF+ZU/JpsS9dF81tVSh7dm4jUFpBSieJnhAcYsF5FmDHO
XHEVbwH9Rmlq3kxxDEI3Qk8hocY+bpjk52oeyv1ntmKP+iio9AF2HhOI+caebviX
FG2vWAUltbMk1qZG6u1rSZTybA4MdDoLaxOi5MUD8lyJS0Q0bxm8PLly/UwbU6ae
ujaXA0SWRYayLkGQ02id4yKO2X7q2kL4YHyTcspf4n4vOwKbcJA6tW5FYqZXrzX/
Vdk5NVCoC6G3+u26N9Z8+exYc+dA7DztqEdY8MQJWU7nTZldcidCgFebC3bIZitv
4YvToqa7dftwvruSjIY5REHufocxTBs4ENbvX8ESDZUWk70SMHVBmykQdqhuBBaK
6scK9IYGY81ICPvcKp2KqY+vkSALAs0ukJAKQ4lP7troEQtdgFn3ykOnRatqYeF2
8PvW/BV+Uv8J49qxr4NlyHHpGICYWwCNLoeheCB/qiCCRVN9CJyGdZi9jTRjpAuc
3LKyO9dknSjYdOadJ0dNxz7aGWGL+xuL7vDfW9AI4WUKvq9UNODY+Z7PoRPkwgg+
fzwIvXkaLqXeyWXMXh5NeVubHjpBCxpmtDdPRAeyX7OPpJptrvCrdYEqDWjSUQFV
acbolk8QDYMWQr6Uryeknzxj//WwTaVQmWxdJhkRCaETYVNf3MsG6eqggMAcW8Dj
PErBL2XC3fFA/N87a7FAt5VY/0mfuPZbziYJfUzzjTILD+mgRTYMTnottkZ0a8ua
hgeDWv5f7J4IqDi5NYC2+gGsVxA2eqqVauqBrjTh81QwZ2+b7fHZlLzJQ9aJz/f5
PlgeTDo1CBBbOhZtPTQbFEMDpyYgEBT+70h/fcP2T4HQmlCe9rJ0TmOdwYugfIjN
0Xg+98FGfmoQZdu2bTgINkQJ2n0uHKcRd42f932to5iRGHtpyjTbTnDfGCXspj31
HJC53GyZenAC98NxqgMNN+GzMhbc9/+5jzE2qc5v3gjHjvLlUngcC5wUQ7v4veth
4jkAC3TPOT/+E965scG8XYeac6fyOCMTd78KzguCuGaHPJ5Z/hRV0QDYQ0T6CnqO
Ha/rj3vC4DSy6G39GNUsVdweN3j7PUjNf2BVUB8rdQbvRwzaVBvfR6Bcjok1vwvt
WmGXmVbQQW9XPYhaeetYCPVQAZyPtQGkxxp1MOaXkeu2bDj9KGtAQZ49Km4y6wPz
nemK2y+VmyOyq7v4FJKkOg694x0AaUXuuTU44UA4iO8463pHCOPsiiFHfYRyc1EG
3tplwa6l/zZaillxh4ffcZUzfnaacT1r+SWqg/ZfgNOKDn1o0cAWMOyOBx6J6UQ9
sTpB+/E+qFcsQ6B0P/F7hLTFg4X6+erpHE55jPggPR3sQ/voOd52eWdWuA7hPej5
Ybn4p7JbdAn2B8O+eNK+k6eGfVMUNA91VJ9wLz5eyuFVbMCtIDhWkuVE0jANEkCQ
GQan15NmnHbJi3/wUwPSGJG7JBBREsnlLZP0TM+kCPlwnWqoKuly1kSvJWKTgFhB
ZvMKW27kQHbxK6RIqcE3p1/Iw/rndfCZ3b4ck66/cuRbmJNL0qpjDWqED3Dy6j2v
zxAlSp0dzAVQ/X8cK5pXK3eIiTWT/Zabs27M5VZcDhv21cEQiK8/+Lw7t6Uw60a6
N23eDXgHSwNCEcOkJ5zVbCJo4t0KaQmaosOuY7rgIxx+J2MMLBsAfGxDq2rFLR44
DF3Ajj3SdesCRj8PppuD3O4qG5r/5WvH/VT5Brn2RQFvp9zSrW23RlFLdKQY8inI
AGlrsenIqfYi7MmWk2kdsXdJAZQK0Me1uZf4G6bNk4LkOLnCVczi3LOBQZ9NtHIJ
AgZ7aCelmYOzzwFzl35SLOoNOOVwazmI3J27SxZiwBXXCBD3FhXC+djdTE5B/Pwp
7HKXCGIxeVIMHYMBY+wJqSwDQ0+oZw2kDzSn/3bPDJuamr2fyPUZAWsULR6SJJEB
WZ/URBGSyboEdLYDWV8DXn0hdLrs3McVzf74lkV9R8sbNXbd0Ip53FDDW3PPlh5j
+khz01HQGnPT5OpNMLJ7oe2b5FJLSq/egjJSqo+7nm445KjCVJrud6KALYecqIWC
IT89/vRv5X3D3sJECWFctk8jDHQZUg/JU4J4A1DAcD5nwONEDA0OtgYdSBDkg71o
g2CWFhKu/+ASAdJBkZBp275nPP+U0bZAx/V9b90rt7dfai67tRVYlpH0x27iKvdp
M2L/BWpNNw96b02w9IDMitZQ6+lIfZE9E33d5ac9l7Jsl+PU8hMKrwglZaUV705w
nwboGqs3I6QDbqmhbeg+8EB0cWqy6iBg8XiQNkfFFq7SUmpI9/bnUUGm2wAmmsnc
Ih3Vz8gupHDBnsP1gLx3iCoo7VvXCIHvxuqMUi67ourV7mGCCZBp74fYx3+r0FM3
ovHA4bqGRJMGv5Xe5w+jOEP3ti/PAwq+yGk274y89q7rfQUiRFlZqOCLnI9X6zlJ
1u01fp3t7RoZco1mOjbcmd2keYMDHokOtL6QrNcFv/S37qy9xZE4sUidS08/vk5H
WLgzO9kFT0ALK4AnvF63r2efOEjoypN5G5r94e9cfSHgfFMxJeilSWPBOsC04pH5
8e951uf5XEnQvn9wcwM5Lcy1dMQ4qMTWo1+1G++YMZHfL1+nYI+RMvJcqxChsDpZ
FZuAZScMp69DhDu2RCAu7FIEEZJuQhdVJ2EBQ9+iUfuNZZSSWlniL0HqfVf+86Lw
9C4vxZ9Vb+3wc9OyhjaY8utUcY7MHEC3c4Uo1xaAic9+Nq1mvv4iScB/xNvvII5A
JDw8Z5yMLfaTUhit2Qg1uWdkesRN/+AGbUNxWTVL12ba9NNfREgkB6TPzEt0d0n0
owTu5+xObpzLLX/YHNo+vXX+sDJCyV1g/SPTetLjA5plK8lCT7J+E0uAxfjf1mgA
QO7XXEq5HXjgcXmhZtdLfG8xVj6meeEtEbIH1G4zxiU+/UyGOKhkdy6JmxF5wRWh
nPb9TDgnxJVufLiWsk9JIsUdfqYqWb2rKDbA2D4aRVj0rpU8s5AhgyBdXkACugZ1
hCU6/3SCIDJ+WBNTj5hZxe7VgaKAs6gNuPcZSNb0Yb9jvvP8gpjoVuYGVr++t7tQ
hdUpHuJg/XyX2qumzUxfNjviHoOiPOqsobt78kr0/IzzVud9QRRcjFdkUzuUn4gC
RFCQ/TQt5NCb5/RUbhXJk/rvVTG48nLHs3MrkvPJiBZDk9Peb5hVMkRZLTMDm3bO
NzIoCzdVcTvwWDG6QKzLivoNTHe0S4bRWjF596wkZ//sUeNp/qNquPG+0hhKK1PF
i5cVkzwq/vgDAYLiJeAwqysuS0hbN78Uaemols90hfAOa399bsgeHMMuQOqxVdME
OydUBahDylVeS5Y1qErsNtNf/5UaUcSxNS4rK1AFbtUvasluhwP/WmwHtFyzPM8X
cNkI6q+z3If5fFDXBAGi5igKhb/IyXzJhebFsVLdAOe9HiRD+e2jKJ7EKERA80RT
XKrg3OcmjJCv3OGHmgzlj+A/0TAxj7x2OUSF0tSul4iTZVVi7lwqb/4ZzSIc8AWT
CkSMFcT3VDEcrkcJDTzGZIv+R0OF9NrT8a4os3yDpPv/VxLj0DJfDfXWXXMlQ9Uq
TxhxZyeDuWBN39oQNDDXe7QjCSkSEP3U/ChWJCDa/ufkMFqQ1b+VoKN1pB6MAFow
Uhl4+otEj2CLT8Ikag1qcnCm6VhoaDEB6Xae8VX47mryVg1uzL3ImHkuz9S+f1js
WASUY7bnhuK372ivqwpkMjFmuJU0ZhFcrcCeBUX6hv3h0/r2PnXG9osj0k1uNW+4
/imLVIE3XNl+tgBkiIfVxk/vz0vcSMnCSlN0mm5/JVz7FTsS8F3o3nvw97mbvpiM
l6Y52VNH1cKgSU41BsTmKV97BKhdn8nsjHBzajnv1RBrmnzLsewa4X3/VTCWOPZV
QowghDbkNZaqhQ5vcFMI0wyz2tEL/QDLuC3UQHZLeyaqIZKnENwii3F+f6OE/KUG
5zzIcfNpK//DJjs+AFMYK5KXFzxnqnefQ1kHVUR4fIyiV5fFNeTgB7ThisnIoFsy
gxk1iIjn59CqxDZ9AX10cooXBX8zvXHfakQrS+bcXCnTh5c898YP4bagoqWXOAd+
ipwU+p/u/Tis0P2lR/nwKNXZN/tylDTeZxNbmoX+KwlRxpYCT8c6hPcRzEM/3EO1
sqlcVFNTspK4qCb6kjpBQk4SLcAvfGwTPmR0wutZwVNMv7xKNV6WmgY0OyhpVSgK
/eJWV8l46TmF+cp+zoZi+jZ9LMTQyrm1g+Ns5G7Oy3CLkQBtzYBkZIAUg0YhZdkb
lVe+PztZGxNUgBq+8kl8ZabF0CK9we2lUOd/WevSxzJ+TzcskH5FmOiBm9rHg8Fn
Rm4kDoHvQ25S6byGdlTYb7rKTaLVMS5/x4lWIXgIGl7XHBt6Xi7mZiw6HpN69crB
S6WjsmCtG/kw5FoY7Mpbj3OC5nCEMeRoZuP9ZV80HESRVVhoCN9pim72oWwimuD+
WHSsJkYb0zO8lsvF7DTnnS8D+uW2tJztnlCsz8vz2p1x46ucLj3RD1fJpH0//WaD
6HHPZVxB3trUJcP+dFQ5kdS0oFO4JUYLgO5Ec9m1yvv9HOWv3jK6aOkSLwNVMm5B
q51PwyrBay9d+aBNRVjJjvLCMEFXQytmopcblalF07VPGpTlpbTRS8zAFAJq285m
LL9P6E9tnR3qPl3xRiVF0VVxsPGtkXl3WtcDtF8e1RNJbGKof/7ZO3lugw26LYZr
SJp/k2yLaNx807yxVW2fxSaVXyqA+2YSFG6mLnKgxWWcWL7559ex1kJRP6kbm7o6
c09Qga69IfwRxSrMXqvkOCh+s64O30ZnMdJhuaxQv6kt6+YUQhO83YLkq9DP4Zmx
VO1E+XQAPN6uQiB6Gg6pej9LWJIqno35A/gVd5JrOdZfZrJcHLOq4Qejnj0COrVr
1rgk3+PsiNdozciZkY6SXwEuDPsgbL+vXBHCFPXPf6MQq+MDtJMH5t3JqDdhhApr
DjUlhMuCeHKMY7/7oJ61aEDE72iStkvigu35ojsFnv0XtiR3zluqyDqY0zzE5+8g
RqySIvz+Gcq2JQYBIOhrCbLpwLapAvaY4NzVLezVZQPlR4du1HfIF0CBvCN9g3t0
+R04y2/0VYzEAJLkUivSEjEFmCPLvJJB8DAoD58JQYuwR+HHFy024VQrBTNPh9nP
44mkx8M6ButbiXI0BDfnHei0kKpKxqKe5eB/TskpWgzFrWO6fuhCoDAem0096T0U
9HlYiSb9DUKeIyqP+2vA3uKUBGc+6ZEi6gp4cvHQLyyFgfaA5ireIffEtXc2v4yd
sMotvdktUuqNIzB9J+VO7wr5/gK5OB/zoIQLqb8Iqu5IjtydqbNzPoq/E+E4sSLR
Z5PQ1h+s4ElwTAQiolWlzrnKHGRghgUdT9JprsAEOznxGDQoms+mDDbDQ3IFNlTR
kdXcLJ5rDXsjBTnFiEqyefgH7S2jBRS8Ss7z8roGbOeOKVBmO3oj+OqWRp5VOOhp
RppkfIow8w/FDL9LNhoKih1Y9OemMGh/mJYKgBMndmnN5CxbG25f8ZWuBcc4NNUG
jcVTlBkrlydOWeyfLxRG+c+e445pQfHuonl95aw7tnv6TkPjcKalJ1GCs4ieoSco
C1oooEe7N67F+ipzc5+G8fcxuWf3AzHkR0qxj9EeYNc3osyUtx0zeDKmPf/pvI0M
x6P2pottM+2csgwweUyClbxu2MzsIL/wUIfT09GwGvl+TUqJPSNG7zpYYLlovVfL
VKpCvEMA2TL+jO7TIlSiTCpWYqd/EiWNctS5gWTc+V0qqZDoKn33J7WTLGC3wMDn
p+JnL429KAnJ1eFAbDyiMwKb7pCijBDue/4wbN/K5+e7SxTLFOH3hEDw8Du8dQ7D
yCZ0hGpLO83mYH+u4gX0bxn0HMYeXUsgPfSSjEwoP6m0Yem/juc/5RbppnCPvn8p
TVebtneuNjqb+ROBoP5PODV8G9/P2G11r0g7nb7/NUcJC37/EWGfvf+fWbLLvfpR
P4bGw1pYA6ACUJLboNpKA/mFRvtOM7CJg3gvR0pVR5iwMGnPsWOMAuAo+R92LEVL
KH3t8PrqEiM2Qo7g/HTNvl7QWFatJQZSfC98Sy/SByzbrETf7a6+eCZxhg0HJiJo
pNskIVSyvMv/gwmszKArJQFTrr7aUG3biL5Mn3k6LK3rh3mKyTctd9jsq1UT4chN
2oIZQgj1OnOosrkGGSIDXRFFZL0+hpAeeaHyCBF3KEgDNAhgbkpJf3iIDxOcgsgO
1gAePErt1VuLXimbOWZs75hsJJd5gE2+yQah/pEbPmgG+bcwN3gXrEoVFBbON4Bo
vPb54Ob2z5jwp2Jg+SLMYjrI5rjxkBO0Thkb23yUYnpHmqG8uirm1LyLUESKXDwf
oAkrZkk2vyTVTrvs5lR9A5nw6wLYGnKdraZK34UVxt/k5jn+zYx3xzOl7fK9gRbv
rkCtjJGYoPfM5gxnfGEoWEGtzUdgxUt/8xKvh+BcwbhLaIRmedY4G6aKcwNSOgbf
7karxVVtkhlSPCClu8v8UziBWcjq7o4BDL8vEOh8mkk11r7E/h3+D8KQ4fT3wHmq
O0QW1mnofAxv9z1lDYjONbtC+MKgoWED2nGjz+mOT8rS9ObXpCfEeEJ9rEEFDW0l
NwWCchJmMIVbTtTNYHmDhB4RjC8dBGygmjj+KDp5hXzKUgqiRq+dIJPqzvsW4Clq
MW1EfQ+ysN/+vbY+R+Qb96hROeotgpmPoBJab/3/iK3VmVLq4iCnYjVJ02JlMJ6i
iv7Duj5RcjOGf0d16XUSFVyasKP6ECjL+hV9c958Tr/adbYKPlGXCht7JB0G/XiT
JaGH7UBU1ulmo8hyKx1wVuUkJ62Ss07ZAhZJixXKaRx78PERV+Bn6i1C/dX+AnSb
NS+cRKwB2HMJmCLQrXFz7DVt+9Qld3njZTHOonHVS3cvqFX+LNITD6WLYJUalCLp
Zztlov/+7GTQ6UK02NGG6cyFUkq7SZHhAKRTGZXgS/uB+VQJWr0kfZyp71ykJaK5
siMt+lu9hE6Ct+nq4zShP454BZXkDqIoDiyjEevV+H1Mfho2FFpdQvKUyJ1bIVc2
sBvMhs8womOQekTsswt8ppxq2dOIwq1TuQa4zgQ1LkceG19bH+M9kN7J8GcMF03J
GqSakLuPsfZ+XUv0SdkSN6TgUjoLAwlQ6K6tuBIu12pBoIftTA85NGx784Q5v006
qTi0ZADI/vLepwO+9nTX/1Xk3r6hv0pssEQ/1XOW3BZYznnk/eW/DJ6J9aTyLNES
Ar5MiUg8tM8iuLMv2gWCwOqYtX9Rh/Hkg4Sqau+OadNWCKqFJK/QiuMVqGXH3Ai0
mbRk5OxOPbgNHveHfk6ECUu5tJV2O4MIJEfAG8tpvZt54UVZznTOaQMDt1AmIvlJ
9ZPgGjL9W+pN2vTss+SMegp5vcMLQ/B9A1WAA5ThvPWR1zlXbsrwVJ4rcUYu8ghS
nSh9gYP1HL5jrGI2KnbJ4SagTiO/dUiQ5/t2FHmKXrrAZQy9y0TjkKjlkU140yw6
44Y5fxoPqGvwnPRdIhHVitH3HOXbvvGo7iIgqa+0ycCupQ+udGUENVROTgoA4gLJ
CLNOuajiNd4j5Ug5F0pS0bKKhIA0zpMkb39R8jhq3Kp1l9wUDLow6BK4Vo7lsbvt
5F9PVc64v/Vzzz+g/O0fZvqwbTwx6rsaJhAoVhcnETMHxId9bGyljILTWVLl7377
udl1eBKQu0X0Lv/cA+CUJlMdsKSssbVjVC8JP3vQy+AEsUAFbbWZAg1CSaze6+jr
IN9WAEbApDDRzIhzdf5PfGCgnpu7yi2oN0SG3oEmDoen9i3RfZuEuHdctAWYO80t
BNoKXOvNfw8fwmtmXCmD7q/MB07BOfIuumWw5n1MAnwtP8nJ8zEU4P5l3J9AiLjZ
I1IPm2XN1vFpGO4d8tQ1pS+CEsTKmGMDZDtbyJhjjG2bIjDwK4X+e9ncXKPpO7SX
U5z2e63HO1ZHeGv7GrWkzZh0vc9ZSA3e3gY2+o/U4Sn6vyd/4z7+dqip1UGiGiSE
uoJ6YMhOntOBUqM4purQGsebh86LvZdTBJqF6/QYdI8hR7vQTL4oKO2sd24syRFd
YQkcVSjiQMbttmXkPDKFi5mtqXTMWn5NiuzTiaq4TS7izJ1HeulsqhT91AcVLzpm
oziN9I2F40jVsW61Tww93DVPdH0gK8g0lPyB16MGB11CH1N5N+G0hMfLRFCjoNPz
DRCV1HAglnzRuUrqKvca88f2MF54sU4YxN9Zb4OG1dnlxo7VE2L1UxCJfU7fwUJp
erUPzjNujitUSSpLZeTLuFpZTVXvHIBN5dlBCyrE0FSB0udZ65Na51xby8fLWF1i
+gxq1HVnKfMqEdPd1+9tA8wvMvrGYvIFiRV6ccze5cJsz88G/ljCiku3gZv0YDC3
LCjQSAkeXNVsJankj445jubPaXBLRoK38rK51eMUjuEvY2U2lmOTvjEwTUKSxDuK
ycnZTgo5vXEEAY4Ouzd0TJVAMU5fNNdKI74CmIUaN5ya7c7xdsIenjhq1Mbtm0wV
EtwluY7/4A1vylMEaXmwa/O0WqxWiABP3spPXZF1xrgyBEUVfgvzJrA+I+7qrZHX
5Z8LdgwdVctwIsIKzJulOuZnS4KgbccmNSwP8njV+dibMukInwoAv8QrcZF8zPPp
L9ftUliZ8cm1a/asie0b3pOo6H/P83zYOVZJCM30MZafLhh4uX5icQBybwKjYyaq
e/ddSHjHx0r7g1oBXdvoXVK+A2aJywneIPtupKRZnqdwwg/Hq4WR0Qd1TnlPdBZD
yaCdkrvbLk5ZCk5DWslJriEX7PyC1y+IKABHaoyQkKVbratwi/E+ICDRRFh3ntt8
Il1H2KxzrluktpJ77fMz2SzORgKyUHj46/9ucFaLpqQ74KxINlEB/TZjW6s+8UvE
O79IoUjjNBCMOtXtfdC/gh+aIwj062ROUfU18GQqwAGYrA/n3pacRNdN1i8NM6Ui
xiTofYWAet+WH/rWxLCfrslaD4YcyMMf1VdtrTNkdtOGa+guFCVEqjwxAy3Yq/a0
X+O7yDxW0x4+YnMDJTbEUsBWSUUJeJVQd2/qiaFb9U6m2rlrBRH+2NXoIrOHCq5P
tT1+TKN+/U/z8wfZusGyZE8uOOWHtUzI4gBWrV9OHfd3KPXs4oLalCSXQ+9gtJlr
4UBdCB2/fG7n1ANLPqubM0NBdiYtUpiymMMEV2I760MvV2o9Ty84iyNyBAYRXrPW
0qD25p3MchN/W6MU0/FgbkKppw98LWuZwYq1LTg6wPbuAV49Y7x4oa/eSTl55Dfq
0Sh7ZH/leO3q3vEI2G1ZynQi+aNlAPAN5VodgIU0hRBS7dOoV+pxTDCpmyGOgj16
U4tz2c3zorbBCg9pjeFSf4ABZSrqdkUFktgbABcBcXhbZa4o2jq+W/Su6yH9/c06
ASh8OO5/XC8KGLey1ZodP+hN+kShuIgI0Jn2ZlJGKSymnjj1PcYSUbipUvTA/3mS
3fEAf9BgPeLz2WjVddVEuFi0iUSDdQ4kRpyEHfB8gNZx/k5MFdmhQIg3ehC4GDn/
uu5bZP8EztclZ542go/Twl9yijKLgEqNiTHe9hpmGdtdX7lrj+CI7kPuoJ39cFN1
95FEda0tUzmhgsvGoVTaJ2FAXRo4zFu7+20fN7BRw8LVXkjCi6RP9ncWcBIV7FPg
T0KS4t4n5cj2932Sim9F1Z3ovOtYCHDgwz3XFbQ15uN+fcqYLnO1kF9ZSlIQWty0
3Em6fjVHHj0dz6N9GXUyc/aaDq2DgsSjVJuL0E6h99FD4nFHOlfak7CGiRQJPFep
7t+PbO3pmMQUWXhLdUCtCV3lclb444AocuWF/GTiIu7V1HykplWII58lklR18QUb
Hwq88nXTD0GX1xZFKOjAoAriMEaPHzzDvQsoEesHQicoU2hStFQBfB3UE6ddGDao
eV3T+dMVtvZwEbVbkK09lyxgsBRsbdOg69mrUVDTCYDYDA63EQW+UXVEUUl6R6C0
Ocpz/DCesmW4BxDyG/09VwhKlCvzQCAcC8xGbH0dB1ZnD4gDn8OC6LwNC2mfeZrM
7FQPJzAbBC2iFBoZ8eUUYaH2E8fPwx/UFkZUiyxzPGl8Hn/rFX/nLknmmIpTpiXt
fee1M92sBKnHKSBNPJouh+kcjyX52F/+5/crvVOuLYNzi/sVs066otMshIpugS2M
hmCeov82KK+6jVJduLNfkrayu2/n1YDcovK0OotNN9nvX5QUGo0QOnjNUnDov+88
00ghWqPQeaks9ijUE4az1ywYH196rENKfyFZE+li+73+Brvw9TX6mo2/+yALZTAU
wEb6sxa5LHlhIVJgBfdEl+Si1RqNxh6h+zjJQkrOR4s82id0whNJkddLv7aX0YAa
2qtcsxaKM6m6VeEpeb1b6z2g5tgRn8vH2NRXWXKGCzu1BQmO/3X5+xzf2IxjpHB0
C41rwRe7ImEX08ubuMJx7TMEPSKvf8Zw6+Sh1JeL90EV1hST6xRYH7d4Ze4pPDM3
Ay5Hs69L+1bRJJKfdRlo+WvGO6NWsaxaFA3rJeM1Ew5vtFq9c2BVWuIkcj7mPhYj
lqlTL7DSrWhWV2PzZCyzAaOblDiwgwnifKwDguYVyukLiA44h8HWRBLALe8PmI2T
DQdJHI4yeuT5f7aAL3b6RVWj0CMMkLsAYDvOETKLotFpEWQCeBkKFCWZAOaEGPil
GwmkTjdtk3l8V1066T5ym/7/8za4+socJ/zPKEJAfqliA2CQgh2B6jiVEDM6H1cH
Ea5SokKqxDb/oD8qe3w5+zPrDsMletM+BHpsnf6ru9n4oZc3Z8tBz842uWcUfu44
kyPyt277nlItIi2X+1RLm8aMpMvyWaQ0/f1yts/D3A3qAbALiCN2sD5gchUp7H3J
tUI4GsEQwNLvEwH20cbgVyr9sNbwreua+2e7+LcrCCtSUt+iVhJKgyLYIOKMziag
Z/4y8kE4/oqfEAc0baPrkB4dMGDjdpqRiR6arjuMt9tc32KPhkwsNy7hbX35hC0O
0OSaT6261DffVBWeOHvE7jrgmQBJaGsX17hDoX2bU/uAF+QDAP2lEPy9OybXbBZY
BkrNRGzNfZBpAnYadNDDxf35JqFWpbfRO/IZncRtd3UG499vbbAUWUkjsyDOjULP
EjuatU6D9u9lMKW0TSLE9O4cnEXjFmnZZDtTbMtLKGE9dmdFwfJWgzr3ydcr83ua
IUwWGpctGzj2Z5kXyJVWjFE7ilaFu4hkkLUojVbXzZGfQzY2Mhl6R1Y+Lv/prb0O
Fn+55mDmzQ9RAGcemwb90QJfOa7pg4wT89R9AR8Kb6lwvDHBUGm34nkOcKvSeQFW
p7ck9cZNjMgIVEWsQqitwjkxu1d08HTw20RQg3RM13/VwWbPKJJzJpxA2QoTB4V4
/OqUWVI8HNVXAE714NJEEln9ijCebNvl7Xjo7ASAjTyTgy1hyR529X+ivnnM4xeo
k+fjFuHxj1XHl+999VQHKQbWIZS2HinNFdJD/z66dLVW+IttaD1tFq3mLKxhOrET
ur2eFJ9Zr2UL+dRmJRt3as3sWrIEVDCDH72QpPPOk9ahXDlfTdYDX/AyNWRWWP40
v5r62Z5KLpsIquC27AfrJExjZ9qR3buCY7b6APr0kYk/vhrHsBFmXjgPXh+q+hns
Ur6EEhgfO9N21FWqNro8lZrrY64+QUwe59ya6r0jGNOE3kOfJGz1crFi3Iv89SWq
SbTYdXAMHBThv/h3c+8Gn3i4gTfQsb3hzsVbS2RrwSXB3gIIxx/rVb5+BrxHDCjS
PILe8oxV9ZKWU7LOjPY6Of3ncT4+TXVBjJ+tBjcbsiIAQqbRYGQUuaZc5HPjjL8r
dWnkKrZGuq+PuIa/wTLKwjH4Q9ux5JxJnf1iBBZPY6NfY8YZ7M8SNIM7V2WqkIVV
h07BivN6oMXG/J7OqbN6fz2Fn6G+xZiUu4m+yDxjfx1b8QV4soucoXaE2Mg0bhYJ
mOyUjTIRzYr8su0FOfdXr/TiRVWW5+NPloGi89UtS4jJleNI2A6sqnZTXStPcT1g
J9ps+VsZ2ajKAYdU0WNo1eYYpEUdMVPRrPGW+ane8sj8LPRMsKLGvbWdt+du7eyY
Oy4b/yqBPsjZ3IGE4umDM7+Af1ycpw9qvjSKUOogdjr+kwi0zo1X6nCertiqiJy8
tJOks4xpe2ukMRaSvXa8CMVgR7+RakZlXBaJBMHmGyGPcYMIK0qfykxxjJPp6D5a
QNc0Bh9M/JR8pMxTSam50U/3WoxRPkzMalERUoO6taNZ9twDS+ZGF6gi9rv8p/Np
AWABAoiWQpbg+6QkCyq4znDjVg9cBBYwZ1QsXCoPDJpyr0ZjlM5AkGAkvuazgkK3
5x7PuRXMqhCwnhygoUu55NOYzpnWLQw7Apr6nroVHKldxeuNouBsmyioylA3Njt3
gGlctoUNfnLFEWDqmO3f7ubcrNVezZlrHR39ROp1NUkKQtyHo05LQ62O7eDh6/Ga
FS8jEZdjeEDYW7XBZyPC48OOFK0Pa8/KWHdHROKHLNUYZVPjwHpph8rbC0eECnJl
iUwN6e34Ra9Qw/5iK+x8ui9i5F+OUqSQog0eqk31nZJ7bDXW/PCglyX6QcW0neDO
3kR50wQGalmiS4Cs8gZJZf1QVXCPDODDnxCHdHvb/FU3YSLIlpgzfE60JUKjtUjw
lSVUWOhFEK/7VoQ/zjdcde/OqxQX3Je3z6RqGcsvKk0Q6h6cq3O7b4FOcm/QUmCG
N5roF0OP7T6ueQzHvyTPYt6BSl6qh/NqltnPi3VsBRBH3gMetHP9s8RsoGOh6cFT
3zgu/OboBlSJNKUgGtZx/J37LQLqLKz/BBqopZKAV6q0mDuqgOD8ufAjdpDmiy01
93xoRlw0ytgnpTzdY8DizFaxRojRwkv3zT1v8lYEss2BQ8PzGvSRoV8ZbACfZm6f
W32LsFzTYQ8ziwaUHzVal5Kl/ghNwDxrIHQ33ixJBjbFOqaxoC+JdUAkhz0+p/cS
7FjJrgyuUYWW639EkzIG/1z60Txd7Wl3r8ebIVcxyujadW67Gy11PymXW/Dh6Z1q
swYeXuByI7wvRzyfgtWfIWU4+pDnv3d6AT0dDjdy0rHj6Vu5c+EJ81pzxq0Ib0+V
NJcNOYgM8TivPfJmtqkMtOEcfdI0NbBshkS1oPFRHgMbpzloU4mUn5XSVisZ2pyJ
XKlCJbVkY8aC6Qh1PGU6UgxP4Cs9JspbckUqT7eTddqevaghLNY6YCpO3Jvzyz0X
tN7LgjfOnvjOEOkVrcTitLbpF5fzgP8UBP6m8HdQf6SQ+D5XwuuLsVr4oDjfRT07
80tiYCFA742/emgmMpERyJ2ObRzAEA3irz0qVxLU60kIRrrrWHKuMcrEKpjtuHdC
tHBiHK9J985saBV4IFFL6HdRfsvHYHSmh2bGZRQ9Zd4hwUiGAJozpS+fZlp2uszh
AP4dBbi0Bne10jOT+KX3RF5rZuA6kDMpe2bilbxM1NBQbOTxYJ7c2wxUcarcdcSX
mdENh2DBTJFAIvZxOQEENPl+QSgpjkPk/CkLUf13DOBS8yazR15hbn/goPAtZy2N
x8SG8ewWdp/NEO0vXStZ173sRSD0DOWA3MwNE45vi2jbg8aSQz+Nsf0izMt/Vvoo
HFOb/+A7036vhAWQF3GpJpYrKXQdTmdLcQg8X5Fuzfi/Y+/EZ0R9ZKwcAYfZgmZc
R+ntIh0n6Fx+mwKP9TpucVNEcg1Ndf7QOt3vkHSuwLl1/Kw1uUZNN3eLXGu28M8i
TssD9lCO1y71Ej6eNJY+x7gZM2ewnMCq2HVe6i03bJAcM1H9OukSFIyOM/Ne7bQw
e2LDnGs0LzsOeF7eaA2OWeb97UszXk4gGkfbbxrUweSoMerGjaiJ4j3XONJIiWps
+GCZWBcwzM6Ms9IAsOKUJgM+n8YWoChwa981v9eFwUHn/liG6avvjYlN7t3DOSgx
/1yRunzbaJCclKplfsS2eYcCzhvZ8rkiLssdv19MC8gJr3xVk7PHmA1tl1uOtqrf
G3Hlt28RK26DaNtxeKEL3QT+QY5y2riZutI9y2b/hVM13pt7u/hgClQ2RGBAKUY6
PQZOK1fpxZh5gV/BhPMR6lxrd4nMe8K6pZxa70XWYjCXmECKWVNBzjZi0CLca1Hm
0btrIzpOWKCD/R2YKmzNMKxzQoKtqVOptQ478KN+Oj3DHa6FnSl0I0uALJ7S/xIb
xbygbCOehRYP/i0y6guxeqbRIojfWKXLtluCwqeGIBPB1gO85auOoiafiuKiiewI
5b8hcvW8tNmlv/Hqdci+52lNjzkOnWYQKYPouF9yqCj61WGyMISzeLRk22Ehmyd2
z7H7xPbWeb+Hgg2B0kanDybhc7KIkV5YGlhVF/2ffcmWBf6+BxHtNA5vRHNLQTUY
ZOtQygdhIEGJ8u1/FEMnnMQIzg/9afsAWsrIXyMO606dTawD/MLbsJ54v7BkG1f1
ireLHy/A7pORms6zYAUlEy8vsDU9q5+xufTu8sFnn8dVTXXs0GAi2JTpvqSAyWpn
471dMMjs6N/e3aLhNRB0n2OGs7dc4hP5BkRS3TPAS4J+lTcMLUwbVdwQAesuHuw5
Viw/Rw3b56p82ypkQKzvBTvSMidZ4PNrepFLH1JL70ZUN7vfMg+bAx2memiyBGDu
Nipo2obZsP7u8+2S36ALnIavYl00Emiz1lQusSFtFvgSBJimyXWrhEu2JtKzqPlo
thXv8w/jzavPQFCZjqQHD0SjBkq4j/HMpM6siAZoMNVHDBX8EB8qXayolZbP6CXV
PbK4EcL0Q5FL/yL34UgmIuivM4Y5DV1eUsYwgxnolBUtFvtJ2ruI1/mmm2CIxxoo
mEXGUO3gH/18Bf+5eJmqCDUOom4p4+0I2258YAty9d8MUux7D0VUGo2COEWY2jxY
0ihT6xaMd2sivXCO5+E4Z11f60H5tZRz+w5QFBPAa0zJmNzsD5A9GflJxYeKFtRK
+N45P7QmpE91L6XY3RhHQXqBuOHmTeWwmSuQiCmD03oaPHdPK/9Z5qzRj5q9DJnh
IufUSXFBnLFVyEuvGpqKrQNS45USDB+4Lav+RZWQCb2tmdRC0pmD50jZbwKBl23G
bPZsifPhw6Z8Lv5vIiW+LbSKecymmrg/VonbHvBINEZrRHXVgjD2hXrmdn29o77+
FuYzGkoxHiYDYDxQH5u3a9ilwzoumF87k1OoLmS/jjw8Vbnpmu2qFG6qQR8rqrxx
VAaVCb5w7gZyuXsE2NZ6E+ZoU1pDd1uSR66jt8Ftq+ObWfXtf8SMvWRn9cnPt/ry
D7UTG7cbw9BCNJ2q/JwNmZXHxr93NKk4i2QTrxShJFgADKd43tv/BKFpHstgS/a7
PCXqSZB3+0JCAc+LjT8YDEEVUGKVapYGEwU9S5OutPNS8Uom600TooKT3QFOEpxN
ZhKANCiTRWartz/VYivVdXRwlIaMLispx6wloYqk4Ad8qaHAWF+qcrt7DVALxdcH
HNqaFcLO5ELUy3XvrEeXfAvKDjc1q5y4YC/OcVA+RM7uIz98qGWkHX593VVCtA+m
rXmMoZfI/DzN4+AxlYtnSsmaydBaZgKJtskSTxo3TRescIrK+jMsj5CMPRu2l8sH
BFPFoEpNmqi1mWGwFHnfLfp5LBaGNP9JPEi2mh15g3Z93PT552+AzpjkWilyhinH
Q1ywEssst0eeQJ2CiMMHYSUOw7+zT/VjfBTbAVHhdtY+LEL/kC3Wp6EmxMLOCWLm
+45ascpxJoAc2zoLfw/6ObbtfqFe1gGLr6lzOTivkgIMwiPJG4hnQwYhp5OUV9ay
m31WB1+/Ry+IUh8ROhyYnHoK+Tm7NHK8YXSoY0ijsXxVUxtHZZsDAKN/VlDtrOCW
+WnuniIdBiaVurspuYV5JOkkb/N1SKNKoP1/j6GE/Bc70RQmTeLwxrRO6zSCXlXc
mO99NyjXSxot/LNlMOvHcWx/g4xCdwjkIX/c3TY+BlouKNHjd0omVoe4XluOF+Gk
EXtsMP7t5fNhygmHx4h0b4r+Xo9XjQe+VgPlmt2Gl2gAp6QQnFECX/m1Nxoq/Ttf
gcrZK98KppzFT4wyZ7WEF73XiLU6q4rRLBnkfP5Dy2VAPNtY9PnjaQRVuyOXLghy
THGAwR/2D4WJvynb+nviYVtb7zsEZWq0vVvaTRym6YCvWNs9XShinaRHcDOhfo5Q
uumunrR2PmaFyadFAAg4YKyioJ0ah32oXrocnjnk+zVD2U5fWEj4vleTpu2XWmS7
BEOiThKn1N3klH+SpFqQWsrK3ii19mffn9HuEX/nXoeecfiX6Of3XBPpKsYUkJx+
KyfNf9cyGNPX8b9H8kf8tDrcOE//4QSnAPs7IdkcXMTFb0M91duJs5xed2qB03v2
4V1Nn2lQuc5hqNklcbyvI8NfXe8PVAzHtaNhRJlCc4SU4pMy2deeJTFp6/HyZMVm
gf/5AjWcEGJ+3Edg3rATmED9yeG5L6XxlR0I+1jGgWoPnkJPYJniNogYvhJ7CGyu
qG8YbTczASxwHsoeTdaHxpTNZWbQrZyiNACYx+s4vA0im4lyAo27VPYr3Xtt/aAC
ZQ5BZyoNOh4Gs+sr/8oJNpJcvbsEp85JqOYoqjAVW7g+J+HwL/KzWyZ5CbjB7+Tg
xRzYMkOJhBNS3F0qEy2OhrCau744OLaiGuoX6aGo26Jjw7jjcoldsgaIhhR0diPD
+j0O65HBusUEy5VZ17SdRHO/+fvqDKwUwZjy/kpN1ZgtDrc6mI0+YhexTnW/gFgm
DeSWKRHHJyiLVDO4YlsMdfg+gAZeFvhTghlDkqNGhhyJ/VnrRiO9wOnrLBaNg30w
R/A0AHN3n+n/8pDVcaaXtSCQdBZnuKO8tkkKML3oD25Paz1VNX28rxmFPgHhQY/W
ZK/X9hVFH826CYxmaJqTqwDpq33LMtM2ekAKmaNYKiTmhz/wXYcGMzCio2Cnf84x
FMoVs4gkCjeYYFBRe4QFoWdChGADYMmOra4x5PlrHceoUAayHTfh1yJt9He9+dB7
5aVQFhYo/JNdQkDjqEEPG1ppGkJqJK3aLw6ja2NUyOnx7Et6ZiL7gzvndaMysNw1
BB1/iFzRsTKFVi9U6OodhdPhMIreI9iVRMvb7BHXG3B+lZUQbs2klS27yF3z3cqw
LslFHvTLHbwmkMJ6CgtJtyvKTPwuX5YS0FgJoWjaRoK7w0JkXjvJuhgdtfUQwB5z
SEyhLImYEXxd0cLfzl2XzpRXNmx9Svkqpf6a/KGeuGf9kUeuPRciDR8c8CLKgaoi
U25Hn2cNvzEJWvFz0rT9g3ADWZ4GCxYu4XbSjVXzBV2tDxt8tASZ7cjlrm79E+q0
17KlaI+naQSwrlIJjvEjo+FVyY0zc5MaBiCNpmNvVNSV2QQEPaak/kby01cIwmZi
kw1QWw70foRMkCR1KdsSY76msFzY/wfG2BoMAvKb9o5pYvlWaGCUt3OSBOIEKcjd
bySD6DiwIs447+VmFmRHQ963Rz1b+8M2+SBg0/wcgofsMrhGKb8LErznWpbWiLnF
mlp1rv3epg8zaNpUwyEW+HHH1xRqzwt4YXRP7jV4jYYRatl+z9WQZkKYXcavk2YX
r8zZbd6wUDExlPS5oEUs81zPIB7pKoJk3Iw+uROR2jNnQ8SJRmmgqzr8ItGjz8ua
xQ/QinDAAmPlK0fJD/kce3eY+NYkKd44JCjntjuD9U514E+mqdu7k5cEZQwMGQ3V
0LnXRBEA2a8DH01lRLxhgXoxHkYtfMFbpSNgdfXpzGdAVjQY1VZSmsvNCkMVLwr6
sm5Zwj8d2rEZgoc1PcsiRizQxrPlHX4uJrfgEovnxtSjM1+uiBnoot/LZg6/nbS4
NVssB3nl0sq1amFAbDLrQk93px8Fhbp4dYr5DcPgbsphMHwMWYZd3fkA/Pd12SAI
XLPRIa70yweA1/qnLf9J8pe0XZZS09OIkbx1LWmoPVLkOU5hBYH7bTxrLyNrz3V+
uM/UzPqqBWBzVpByCfwScdLaLXZO7N/xnZDOhCBjRLkQlLsxOjoDoAwmxNFNmw6F
H3//GPMDpdQbW6mzgbg8gRaqkq7hwOR5MLoYNxoy2rcDtz7fD7+N7U1g5K09/7qe
7xE8maddrozlw8whXQFuV779nzr1le4qFv1pY9NdLnQi/Oqab3ZATGPWVD1jYvCU
M6UTWJKxyG3r8U4720lGeAG6QXuwCeUQ+krRjM6NT/ifuKVlMx4c/0J8jem88zfq
pOvdH1txF2uB3y2w7etEgfONWH75Y0QO21C0WtsT5c8QZDupENLNT/EfYT/L2sYa
yQyaf7/EG2I/VwjKifMr6HYS9mpTAUf5mTtU5Eogyykvt7K7QQGHPGHYnM4rLy2p
iOHzcl6U9WTVMrTbDaxKiZrqlEMZJpl6aUsZIXC4zWlatzcOGc2QpZUNzj3mlN+5
lwgBvZ8O1roON1Bb5ioWj6sIary0nWPyoMKnEAhS9uzJoST6xBDF+xhULChwXmdS
TFZUAA9q2XHgN/v83fiGcyz/nW05CBYMcweb8atlgmqcvYvt7pCMaNydTJEOdC8I
UEFvsFSgYo9gf/u8vijWMbnmUwoqdBO5E8N35FJCAQFg43odBCC0OlL6FESpyU+7
P8IeolWD2iZmt8jsb5+DrBJujhFFxPZ6xrZ/mGX5HF4wAzzf3IUCJIPEmq+qh4lg
uZCm8Fw9Z+oBkMIXma9GuMKYAimjkRjFml04vmSjgNhXWJXtpd6HiDS4wB4wQ8UK
c4s+Nnq8mnjwjT/5ckEabvemRyZdVF1MEYF3riCKxk2YYFLxerzI9caJyJcYBawB
yW3ofprsWN4+h85a5ESKeaOajDnBaPgIc3Rha1HnPO0tcdY2cG4QdspJOKa03aUm
PCZFmTBPVo8o2NXu0vLUl14wRhveMbOsmXVZObuFxJd88fkFeYz2OXMz/Nu6mE0+
3J/QcmW9unNhbf9RnFBpsGlvRbdCxgroPq374af8gcr1WjH8m67W8GkFpqNbbXEM
KfpMyoks56eSO/SMgr+fgiLnPvVEpAOm7bKA3dq6ZLUxa8ccwSHm4HFblRO0fxtU
SMOQ4TBezCNerpnJzbgUEXzbumqvfQaLwKMEdgVTKjyCSvZJFloDU7LNbNKLJ82C
3CsmVYaWqYsZEhdR4Zj8N2oa0wjEZ9A21FtFYJG0CT+X/1iF2yKcEBTqsmNBaYQh
7z0OcnaMORufRuxMfx3vwU+Nb38kwBSLFBot53pH7XW1zfyu9wa8UYWRvLJXwCFI
NIM9hclJ7ySsUbPI0ADP+DpX6XPefDPBJCXt1oZSBlwe4puOI1UMPiNJm+8MqkCO
jYjMSeYsXZCxml0RQM2uTYPZQqnWk444CJ38BdCPryPo+lr0NEoEuDYq7hXMJ5X9
YgGohVw9HHCpbP5xC+4PjPo2odwWNKhPCOKYPPobQA5n34ltNbHcPD5SsiJzCnZT
25qYbDEPC5d/aRNPbzBHOsNhr3ppYcJBVaqEjXBPjN5vWBXtO3ktQ1bGNz7Q5a5Q
LgjokYUKjijMLlGX+AbC6VabEULIxH/ITWM2qZYOmJC6sQi+oY1o9nXrMk8vXV0A
32RVUeMs73kfoGKUy00pFXSweLKrnYkX90qEzzLwE4R0piNvPYT78jYSQcZN49My
tomIIA4yrCV6H8W3wbXoBfp55QodWYuBeCpofIKuyc37eFBulTSuwdPP3+i0UjFY
6lprv4Jurl/pqv5FP5c6nlsymI9vTDqBsdh7iKM80jDquJpFDP0IuGNddUeiKJxW
vNH0P/O8kPkb95VB9k9DrCpNkMdH+OTdL74Xt5AzNpFYpLHZeVZCHAx1qK/el30/
JqDZ4NQ4uN9TZwZR3fnHbway64mj/BIX1hoWZ5pRGu24WMbaBDT2gR6Qc5A5OEfo
O2h+LiJfcQFzb563Y1SxIWhfTl2GXSQp2HGGI7NGzlkNWU//nJ9U66tK9Ha7VAPh
nFTS2gIWf1P9WRezJrMmnb2PpqDCJFkKb5jNWtg4aGgZquOdrK6cQU8ZHZsUaFRo
ezjDjfyPudPrIvxldstnvtfjEHVqOw2js0Z8O0a9y/skPeeh7s/ZYytrjKy8AVqP
wHVPZSrQ1OnEExTWGvZlqUNIDdn59k8j+wRq9q6549KT6DyHvTZZJ69u1O5rWKIR
aDQzVfVuI756mijoI/pHCIDpg5VZyynYA3GwW840chJW8GSbySM0Rm7TUTmLkFlF
FDVSzVnY74EgDeMFcgPIKk0VrlBsYbAQG9cxulFnblhwWUSMY/R7SjwRG+Fdgb24
kS3/FFAq84NEh0gLFwj+c4J2ypFOaV95E+jSPbYlMe/MPXvZP6tH9sXPJRUtpdVW
bl7gX7sVPBte1FlGChwaguZU6VvvHhkXARdayP2ZcVrLYa558FivgAZZtUD2TONB
js663W7jecOfNdQ6XHvfQElQVm6IjZm3v+OyMf1NCVjwRt5FYnS6a8Yoki4RHgoQ
W2eG7u74+vk1ewJUPxxfW3Dj56BGuucMWSVNXCCDYczOF0H3yGvtAvEXXsd0FCoS
Jlu+aVPnD2ws+7pbWMk3RbjwRctUazueKeO/hoPNE+p7xtA8WGCfbhcyJHkkQdQn
hNDbfi5ALf6GRWd7O9PUSsQUUktS6AwMFjDTA1FCXIqKYeUPc3FFu1AQVSek2O8r
JTvzTUpD094tVmYoxVDhL5bMLoLAHJ93Rz7zjtxHVI6ez0kDBhsNVx2GuhUqX1kM
IxPlLfPgOU+GAkGLoQY3c7QxutTiOHRYhontfpXE7v9+RXaH8BkeDMB/5tj2wqEq
p28PlV1hB1IHvVkRdMgzwQZ6vX6ZaYm0hhWUvRQp+h+vmiZZhj0bODBJXb/WgPKc
K10Q41gYRLM0bsj2TVMitz8S5RkfsamrOWuXdaH1A51jt2sCx8lrWxk2M7I90xno
nwpEOtV+5AFt+fv+6ZK83bAA7tvvmSg6JxFIf/UAg5Xtx9g/+hDTRhyaxPxtnk16
dcJJ6FF+f1B0Fm/Lk1VEhte2G6MGRQ/nUnnKJf5FSu30MohCVkbFcG57jHL32kqT
wpD+tQdfjEFNPolVUU60GFxPok0D8sybObVYBqc0gryhKWwcH2P1h36Fwd/r3/l8
Gg2i8EZqHhS7QtYtnQKRjowowjiUZLdzSrm6zhs579rRnjlbwNYualz8xzDr0s5C
ohHtzaMSEpDzY6/09DeVzeIzG4v1+FMPbGvuihUPMYojzg2AyE99gTNRoO/w+Zm3
++zd6OdK2FZ7X4NdXjF21Q3hXYH4YKYE5hpdNyb8CqGpKcyjuAh/LaarPglkOgfo
sjWpaKxtCxT6tDdLv7th4p3byRe3yFplWmZf4xUipmM1SwpQbvEAB1rt074ZBuJ9
UxsC9+JC34+r8H1ZcAwaCBZGZV7XZzZQhy3eN2eolVDxTU0WJDfhiQG81YQZMCp+
RFpAHkIv8BVfSMkZbilnH/OTNb96nmupYKkOPiWA6zxoY9xs9ZWN61VWVS0S5LPY
MLzUPO5QvIXB4jKPTKBYjxXAzg1oFB/5scNbimtVbA6E8oADOFw2aQ1Yw/dOXdJF
MJ9o1197/q47NE7r5fcAb0o0Ni7jKpctN2Uyoc4P9IpbW2uZW2hEl1uhfY5fWPbO
eZS7xQyOHn7bwXHDGxa8TS9wqV2VmNnrWbGhH1CWMKxFKHTblUS+gB9rlh9pydjB
e3QGgTrejYSfD03xUD6aVWiV/fhSJN25NyzoL89tfPVHCBmZ2wlks4bb19+5iV7r
xzLLuOLoeHCyrNplH/bOUO2S+qM6CjWVLkEwXQXLx0Gyfrjv3hjBs1sSRnRPVfKj
2TfuEy7B27dL14dADsDqM95C+kr2oNoXJKuon9qJ3+25dT7iYg1uOVXjLnhFwNcC
/SJtaU4RnXJ0jEHINPAs5i6HNClgtyryvl4MMHhWAl40ob8NUniEUj9SR0MJQe9i
acq7aU9JNTooWjV7X7tNz0Y/95drfciaPLiz/xWDWJDD9PwbesWHe+zDHT2jry+m
otDs2KpvGm9H592Q8yC8LL2q4GNnTgrgm/ZZ4YnGFhyLMUcqZ3Ba1AvcPrE1EgMU
D0UJRp5xSNbLc6QfQCn35+jIDTiXWxt+ZvzZNhNtBe6p1lqIW6e/gGs/GLpnsPmn
IKChPV5ZV8VUILsjywDIYIarqcJ+K+/BPRTvncqB4ywAeyX0AQhvPxMxDllSR9hs
Td1ejE5vzHxcgICl0AMRA8DIB5K4cxLbN3VOzc3AR4xRFsOhxP7XCsUoIeQnDLyU
PwHlhLcLaiH+XlkZ3J98F6JyNRDlc3CUKbpIBWc3M0Y/zhGPhJeco9c6gBO/eG+j
ZSxPdQJivclBJT7hVjC4xgz13hpWM86654+WHV3cdQUFiJWu2td6vGr+wEpJeImx
vamPLSXUnyWL9cSn632b6k+cZoOsRWp3hrdQr3FvMmLeJ2GPveK98ctrU3YeJ2N8
jufNa9YdnDOVL/0RbqrhfUUNMvzxmQnS17HqTSsGj3+INyfLEZT4OQFI0fWuXTqa
HsObyrgvV0Ap7WOtU3HMdSVjNCmPzGV0QQ6YUiUwUUkHmzT2MERIkOTbJhUW67+8
Lp9vwJ/FV4XpCSOA71xPsQt0torzP4SbsiNiBcHX/peKAaoY7n0ODyInSC/Yrpo/
c9mF/zWPjtDYgsZxFpmCU8X/0d8hO7rriwcHRbcYO4ACSHC3kzrMhWUSa+4t8GFZ
JX1Gk3k9ZL85sKhQAkmmstn/xFrKrrunllmR53NQXy9zvd9iUZxUL0sKfxiwWEvS
8jxyzS9/rAZEH8KTbvcvhpMT0XACsCuHTRZmHQc4wgjgbPsDIyIQbFFAYX9crHMm
gBDdDd0swyUFUksrNMGIHY007IIA0kh96N28A734Pj/sxPqg3syj2fxl5FzUoTgC
R7d4uCxzKW5CFn/NTr/mtGWffC4Z5d/qramWjcScA8bnTWmLOHk0LmkIFF2pGPxU
DRp2cn4fJ2mmS3WNOi4QkeGyXSBsnLIGVjwHQO5BU2rm9MItw2JkIBW7x2FAm1dz
LBvqh20wtml3eHKl7tcI8FqfL6pCZfvu2wE4VKRPn3WDfuImttUgfx57+4hXC1Lc
7N0Dnn2djPJMZ5m7JTryvPFP3n7GU/h1fZizmifJHCV+UNZUNOTXaDu1/yjWSfIs
KDuxv0Si4f3NYBDEIBX6ZtuyajKxZG0roPfXBw0aZ+xsww+mlPhXlDAjA9v8PD2L
KFbq9onyp6DeeVwXJ28PzGB1h3cKx1CiPbbmutydo/QK1bp7V2AssRXY6nn9ugPZ
n3S5iIMJ+8UOGFsemPxrC71Kopg1fTSTfi9PsQVGKw43SemuxJA4x5qS7o8UbM+U
xsbkSLlBuzJWnEhdiYRLDPrTM2iDsrcNr1Rl4O583J035cHiZjKFfxwkxRtOV1kM
dnz7NKo6xxIKkKEG7tkrg1OdPPmv29Ka+CwPDdcfeBKyEuQupbuZAmMvXOpt7T4F
ea6HrYlLraJ45DXwiyHp+EEHwHHsk0HMb6BYRZ9cnnuA+w742lifJuNxDUAvMqe9
dDfbzmtff/ZKg8o5nTFaU4KLxQ0wQzS6ANNRXO+dJZk9ejt8rDvblOsaywtaVu59
tLIRl/GeHzrUOYlgowQDYCcxfOMA6D410bq6Eo2ryHbF/A6jkovE5LmYWJf8kTTs
faeZ85G3tsh5g4ixWxsb/ykg/IK8i2Aqoh6hgr8VWGt1byEx2iwbiUgRzJwY+Jcl
WclEMfa6thTPrVqt5f2M2B+cBk+Z+XJO255pzNQu6Gxs6iivCuy45dSQ+DpRx8CL
FrG143qwoIhDcKyTUK/lXGKEdqV46ziz9TI+81nHHih8M1quU8ke/161oZG0R/+h
22bVB/O6AkEr43/npsPsRYINB574k6aUyZYFMZpSpuswOUl40ztxMEJpM60P8dBf
vKr1D7ZTCvdusm2qXDWEZ5xFrNL/Eufv2qVED0moo5WNSvUU35/3BdzuNof8OKry
OK4WtaWHz4B+BVS5eJRdCC1Xc5PCsv0Ag1CasnL12e5iNoUaZQ7zba9YAE7WhboN
qd9PcLS1nYJUwofKQACyrkGWSvzrr7XxHoHaE2a9AVbO48LivtYlEr+3eXol9YIs
D5Vj7jXo0aWLGaputLwOsD7CjmW2KXiN9B6skmZy9lYlSQpQDookH6E11+khsD9c
OqAG3K6iTAlgqrz5524dS3Q9W19gTaFHrbQQ+rEykMc/mq1O3F9yVSuv7m5mQzcD
Sq/VxIlftOwh0Hi4qk6f1wnmV4Q2wt20SkKmt3mJWXFmSeQuAslJ48kS42OGx28m
5/4HA+j95Fqob1X1WcLIFfUtgyBZCrieRyP0HTHKpy+/IcQN9y6hGXu7GqCFClC6
iFDdcak7ow9YGAZj4SveH1QOzdB4WIy8z2pgpYQ9KX3jCE0ggxMfdnKEALRxrh+w
u/bddjM1tA6ftw2Kc6v8Zu+7dPuaClkcxtnZ0/k5vGUyLJvt9nx1kOrU9mdBpsMT
xAkuJXGzpmxzDom126WLHHHa5nP43wLv83Mm6+XGMkobaLo7gwVmuZRy69CbbM5l
R0j+vOhYiMQUwvrtIdXZezToS/ZsoNvnnb72NTGpVvQ8V3hoOvzihHeookF1QUiC
JCDrTKmmz8LAiwQwK82AVhlik/ef+Mw+cjHAgM70+AYO2WHlIfqNkdMEkJOWOOQC
AORFBHVJwwhcrN0H8fbVzKw2MOo1Hi8JyaWs3p86fLtmWDpSspQ1AaF29XUI4Hmi
X1TkketUPkxPT9UjiHXwnguDNtCLF+fr6D3iMh7kVcrlVKONYstoiJ84G5SKOvV6
jGOTHM1uA8eLjQ7aIzb3Y0/Nn9Dpb6kX6WwUQP5uydjwNLaDzAetZJZ4oUoSCFKi
CchFXrnFCi0lFLFXNgDGr9qzVwIn13ssQRrSu35L8ehUv4YXhiuf4Suzwxgty720
Lqme7SyuSiEKjJ//WdlYygWjJHqb7lW5eNe1Re6j3x/qwKcSK8s/Esl2UgubPNnN
45yEj0OFVGfxAUo5nGWmw9oE6cpGkm+koUDRo+ySDJtWVsMbLlh488q5wjRP5c3m
2vVfgXdhL/1IQaczojKoDoCThAyEvCuVN6evcgbfevAysdiOVeNDbIHvYNehOtX/
y+hHl89OcVVb1SO4Ifbtd4JLpwpqnF1Q1NJi4fb0k/fwkDr2RqeAt2yiUixEooIq
XWJNh5ljlwrxZ0dmTrTJwClvJUazz+P94Ic7oq4D3WjlsjGrMWCsIMoTz/oluxrZ
E4dP8JjH0V+EpFCoWNBVA+JKhA28R2QQW41JVsK1Tvr0wNP7ekZUCG/GKRjMVTtB
kXWpxY0CMYrlwM6kt5njRDgfEUbhzdKuytHBgPQsQgV6QJHWhlxg/NlXPnE8RvUy
B0ARTEGZa+DewK7d4g2bd91OIUJqK+JMP5dZmi+UIXGF0cfpf3a5VY/jxkc5TzKo
78AYfSK5mzTLNjhRt3Wnd7z3K7eur3spziZLt8zahe6caDT3hxUYQ4KfBUo3N2dL
Aw5JJrppHisP+ft/tCmut7f+FKlx5BjMkAprnYP3uJmhQFtCp19Md48kKjdy99Gm
tYsXGKDafH6yDHipAh5TrPYbP0VH2DFnLKEzVfeKrl8p5BMESaqmARlKIKJOnPS/
y8pej3S2tMtwzzbj2mx61aJrwRYjafdPT2hSpSnjUDZx96IsoCEvU008oiUCo2JM
zeOo/5j1sIlQDNejV8NMSRzgzVkBil8HBasQ6Pb9fHZPCV7OnWrEcHeeiOLhnZ4v
ygpTQKjzqXo3/YPrd+AXin/kYzRqvARzm0zZ9iebas2iXLqxYu0QOY22YEtHDpBj
9twercdoCnYJXWUfLmQ6kKgjgKKS0Gtyuoe/kGKUrBhzs+Whjoy/bFshtq70w9yC
8+KD/fJKcdU0PCZrfZGmC+CyMYQGCwMlf9h/JSKSI3EdsUiaASzfMsiJ1eqNdyJZ
Zs8taKWP4YCBgQ225+X7MBB7D3eL6WEsduuh8H1LtrlI6LLnzLqkF2U0X63blr7C
AozzGxvQ98vLqFrfgROQ0lSkm92fl2H+sb9jZy7fT184QIyZG7H+BoYNM3CJ0SJ+
w59qNSsODPIIySZi3Yg2aZIPqZE7EujAg4FvBpD18b/Bee4xBv0jfa2riCBWbr1e
4MaujS6WDkpXHrG8nG29AQAApK/LO6WOlVcg262lUiZZBFxRpq2HdpLcf8KY5UFB
4p43s6dZdPkrzvaCwz0oLsexCMz3Iyl3JQO8Fhdga/wrOkMQvrCK7uu4i015FLKP
IyLuD4iFvJn+hxiwnSjL+TEhYDz3A6JFwgc1Fr0xK54WFhPjymHQIFdp6OyuiZT5
KIZKK50Gb8M43cuP6mu2otHALKmoGDN5wne9JmffJibbgO1uNefeL2OVYjZ3k3Rt
KBC34EnGA1y2mg+VR02gSI77CB9AzrfkHowJvoUxN0XhoSU+UkJEjQoqUygbkaeG
feZcM++l1XRqF3PsWe/PuzjQ9j/c5BL+gYAwaRSWRctOZpFLvPnYqD49lbeburla
cTnRSkgTtVS/xmaj9g4m1pGmTgncPtUrHpCFfZI0xyJ0PupXpZIuvlZuNcGPJckw
8//S59UN1qE7Od1uB6CFCFVTQOUpvrWjO1bOXTFcZYwEJSU7kCRYWpDXWekEx+Lc
71hMCVqlLrxpC6xQ/dh5a1OxFElBGlJoD8CTgY0b1k5BMOBp4n7CkuOba44H5Go6
9HNknmrvcaHGaTKzRKNIWGvgAZNEW00I2fC2q/7uAlJ1YwF4kr+SVzjltkNfC/WK
+4GSpD2vNgcVCdBfOI3+8OhlLglNWZtJK6DT+oBbooVL9v+Ii2yumD8nM6deaPFS
F6BnVZhkrEL1x1+AsKvZ83Yl4Q2uxmYfU2zfTd9LEfsjdqI/pndT4SWRiNfOb4c5
hxlt2rAbeWKG3a45VClshRd0onHz/XKvEV2cAZyT7zI1nHOgCXS2kmjp05XHwuNd
9Fc8BGH9lXzz4oapAlCPOLn9VmY3bDB3tOjh264yFhSxKkFEHE9WUqVI5LEvLmLJ
IY/YZGrNLKgjgo8nTGwopCnQbJ07KBrEEAdTLRT7NotM/bw8tzjOCYzqs9ToPoGv
O9wMIMruq+jcEjub3s1tBr+QcLs2ktixK0G9ZHjBQ/FFitC5KIm2mXo3YLXXOv05
ukpP34DLCwT4dt2W0mfmeIRezZ5tT1LBu8R8bFx+urmAeu48IySAD6FGn5GJvyJI
RSxEBTYxi/nLq/dkiRNlibfUUyfeWT2ln9XFv2NedQMP4NG82Du7FXgl57WFGVpR
DDxBnCkIP8eBdEASCSO2VGr8rtvGaPEKsGJJjy/nsthO0fmNutbvQXxKQdU30WoY
ipT3gqp9weo+eB8ANgIsY8DfcHgo5WtwcGMfnKpgaxnhhsxOVs711TKLsB21MBRu
8PoPcn+hT3UEGxKNeMUJuF8Oqd0Gx2pIMK3Ll8VgJRlt8Cn7117RJVrZonSfOAov
bFviJ/Y5FyWc6KRDo0wTFdOBVI2DK0MWbCHJGmRSmNmP65Fgc4DN+xdNpCBWzA5p
tEWacbxigwe6eC/mxuI+Y2MQeEfK0n/ACi7sYD82nPpJM2pO3t8B1FdSVf8Gyqoz
FWkRDKVUrymXef/6lWK+JQ5ljOyIIO2RLRaIw7HcLqMo2n7lcA+XYVcFdNOUeWuk
+YaSkMihfUnyIWYXOUwLHZ4NCtrNqwycChEDw9TosSaf5BoKyKwxrp2EJHoA49NM
TBF6PhpSBaNjCZ5FQMVgalvD9jjyhguDBLQ+C24d3iKBEJbEGLKnuZ9k+XRrJtli
IYxK2NiVjVo6uy4kWNIl1ehnX6b3/PpXA9e01Ror8Zl3eD3fhlS9R2YnsqwnG0ma
FZSTDROxTTRKOEU7eFjY1Ol1aT+PadcqRzX5W7qF4U5NFUXT2aHtEYrC8kH1+U1h
8xlZRGA+II96Z8raGcCsi+KsDrfEu5x2RUTYM3tsjGLHg1JJ4Zj3y6akKs5vip0Y
v8dRjvlz1AoIMhKdsHQNoxnuw4NDHJBvyTSPvVq9ba9zoVZbNd1HQeU4wFOrXSGX
DXPhQi6sJUOYm4zvQXqrrbBOFfESYqYRv5lxrxJ8BlbSmNJUlwb07BT151FOZGSa
hYLmP8y+T4gE5sH5E62VFbqng/0Fkp+Ydd0PJZUgvTElrpW+wxgvWMn3EBZcBBux
5TcwjrTpszDv88WkPHvBkyU3q+TIlaJsznVAi/dO26UifzG/92iuQanyVrhycdfN
1g25+lp0mvQTrY5IWtJbaNEYQjHj+sT5DqdDRFw8tzk4fnBllhDIs5hzKNJRLrD1
m2Ov/8L6WTwoisfLT3yxmcU0CV45ztsiMs7vuV2f0EMTR+mKsE3DcdLAhqP6z3Vn
wtWR4PbP3QIG/H8vm7B+EHvIKaSw1dpGthnpXpNufzJ4i6LEgZt3b4TDQthwfUi3
hQy0waqb9SJiu0KU9MMm7kWMDqyAqHBF+nm1YhCxNzA=
`protect END_PROTECTED
