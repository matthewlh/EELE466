`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ia3yWqtxAIwRt6jSKtGFETwybEQjizJ/1l/yjT8Mi7pV8o8WlqBjzO3o/iJQpCMZ
PJlCkrrsNKijaByIyVkpgYEEayw8Ng6fFLOiC7JOE+ZZJnZ2CorKpY+foHJIM27/
Fc76ByLD3o441cj3ll0kxJHeGIroDo38BMv25gsGDkLpYETx+8z3PXtzaaYEXu4a
XOFw+9NieM8EAG9EdMUEybAUeLZDwrHwqObX5+L1OVkYkLH72QDNpXP+QUDbbZKI
6uW+FmLqJ02U5wXZk6mCIEsouUwOjHQip4D7m0+/iefn1WfDksxqSqP21bLQHm48
ZFkLod8BU7nHml3LcyZeipDMoaQtgd7l2fVpOrkYGbfa8viKT4Wi+0CA/HTyt95B
fvQ+eN3YuqQrKY/LrwF3zQZY7+E0sj7TyCCq0ANpdSkG8+gFLr61HUA3H25wuW/5
f92wQiKn/YdYXoaQoCwDsQJ6Qyxpm1KFvX8gzxe2jSMLaMfFCZr98/67qn+wfydj
J0aEyRLVKqKC9P31TwgPhSSFaAnJZh3XrQh7jWhfYsZ5j0Cp1ugSk0SJbeAfbFV6
Quv0QD65A7Gdrpc4N8s8ZNAirgLjWrFRL4SwF4xTqxksiDTgi68CWfVW7cH/UFcB
ELKfvIkYs98pyKuKUs3IVkpPYFUF0D1o3v39SFE9jOTHnvberFFtdhzVsGz/+1r2
KOakC8VzRb3wb3I3672qpOrE6xlMQzSPeYkiVgLLBBIfRP/IBlLJqs8IMhLgVf5D
iLSkjZQh5bWzwNNYU+6edYPbpm3tSLxeQgIVKqpaS3UHA7V+j4V58p81TqGbtnaq
3NFyGwuI/75U4qgx6NxFolhtcA8sYpYtvM8Hyi+dPJA4PUpq0JDNrgW0REmrfHgH
BsGpuFcQsZy1sRpa/Vt02YbsXBXF0tlWKIW2+ObIsNpuD+/vV/ApdKEf4juzNuBG
5OGF8QdBpKo0FvQMMizQSy2CH4wFgxXSOLSoqPMl79B2OmgKBktEkqn8i0f/CJFP
VFzr4TBonK37DrhZjy/X3jxfXhPvNPGLgRk8WzXFiRIr7JKoYfOnFK1QvgG0RKT7
U5OZ9RbXeq7k4arJZLoEU79d3Xnc5o/6u6LKgMWu8/7Rf+DF1hE8E7ttdgj8MYLY
GCOENqyMTIqpghidQq9Fd5KM6a4TVFtGIXM/zDTfGeAVvZHvs0DiqpLn1Y9t+Wd7
CzElPpLxu3dg1uxDGRWXVAxsla1Mw9/YEiDbQCQn3CRCT102GVSAcrIhS9HC4uTs
8/suZ6eb1yI3VEhIQOCua/GCu/v2iLNtcTXVJnafqjJhaeZwh7vecPKzqy8hGEnR
NHNiGUU+FvNJ8RV2bfBKAMHJaOQnxIQt+R/d7y7umHWcqJdxJLcRk3xMu57jYO96
haZBjvmkC1gmWJrdaLxASRlLabprnPHiFOkGOMOOS7fwgxxdqEXyHcEIPA3Cxges
`protect END_PROTECTED
