`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2BJdsWgC1bGkRlpK24rTqJoHlOsyP+6rGkEZH/GC/0BbdTyAgTc8AkBkasfo8rQ6
iw3xdVodOeLsLrVps48DhKb9QmCiUvFInO2gg9dJ27v3JPWSXeCiIn87m+aEozxi
86tsEhAvoOcFKrC2nCYdXe7YPePYMe4PXpw1t8zW902uJekwcauWTh5nG/WGz/Vm
`protect END_PROTECTED
