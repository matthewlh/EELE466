`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
0YfGYJ8UT7V2QFdJBIEqtyfc4KVaniV3I244cRT+010Sl/uSIC5trhm9lRU2E5w+
19V/KOFeqmVkTFij0oNbh5bZkR/leO89WdszwxQvs6VTZvQhZOdpATU9E239v5eY
yZWLJ8aBLybbmwYpJgGoApQirt5RPku3qSJtWTHxLGwztvSQI2O7mqmMKKz766br
2AWrl30TEtNZatQt3vWU348UzUJiFqn27luGyPzkfi8AVDgYI+x4wUTcT5DDHddy
+BCchcIRjwg8VFLY8dWrMRXNDNc0g3rU537rT4AZQlvjQ+b+L6dtLpnyxGcsiFab
Q1cfZY+nFrHFmsmTrgL5DTyK/e0TT11jmPROnXSjTgev8VIG/YfRZqDICV8ac5bo
n7RKan/ic5gbmFQWGK12/RfQ+zD/aj6CTyGMjaHEsX3jgEBt/S1KdCYj7JprWZyg
XYwCYyq47lZWGm47FuGZdZjRMG6NxkOIINx9z2Fspbd4iyhevDdwkL/YAUMhm6sE
oF4WTMxWcCUto4OsOiIVFdN4F/2roqJOINeSWsThQqZcYXdWkrh3QeCVhdEwfDiw
qUtJfxLtaQBfQtCB6I20qgmUs2K/H1Nt4tBbQvMmvUcMSaREojJ/mwqY9NT3ktVA
WNlDo6pFK4HgoY9BBWYFcD92ffpN4yhp5hw9QEABYbufszRFP49qh/aEtTE8D6uM
qK9c1ixLXOJBRJ3qY5sk3oIfKPZW1RwCGhUXkELUbSMysPFgFkJf9QqdNRfeNkG6
AwIG4WNRUr1IaYVf/0qZlMWGfZjUuA5EueQL+/LxegHXWBhocysaUPc95YkL69NZ
lTAw/hbAKKb5tNB574xd5IalZL5f9xj3fLEfwPhcuaGHkIIoX3FE3bfotByd5xON
ID2CZrTjRXtlY9wZgIwqLQ4I8ClXFVBXtYtNPlY6B9+DIa7hDEUS7loEit+hZ8iX
Be+CnRaPE5xrVhH4kUrTP5jtwjbPoeHC3xlOBUGk97Y6+Es0+Q4YNEpndN4TOrnl
hQVceZLv7YYZVvI0+cqvr+mMXuIlOeOe2uSPv6RkcdjP+T7uVYSZh41HYmyCRLez
9WjRGMIoRdBH9sQuUUgwgPDQkVq0X+wV573IrJMtSqD+qc0OJepACmDSAwo5lXi8
csxJejfYev9Wt+frWZPSsdgG5R1oNlYGRh17WqzyjJwzJJumGhH4LHxpLx9y2j7A
W4BMb6/2ZdPwgH2YfzcRqoi6IbS9iGukp58LMJ5dpSooPHYWDbZzOKTntkuZ1jvR
`protect END_PROTECTED
