`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
raaDIo+AXrAws76IUWQAHt3/QSwNDG0EUgIzF9VLg+hgzn9LBmmRC87XDQVQOYsA
iyzPH9CFNMZraIL86P/m29tfBKXhoS8H7grRwFFVV2vWhfoBUaZZJ0UcFGUld+y/
8jRDo6UbvJ6iXUxqom1hcBG/grtR0RpsnFFHZ8XTUvvqBX1YH4z6h3GfBaidBljp
jL+dD6iIPj2DTBjghWhedqJl/I9L78v6WK3a7+RQZHGUsjy9ZwNG7PDQ42xpbrRv
Lfr5KN3kraVxD3a0BiF8J1PcKqcNdqQVodhH/p91c4gLzlp2dAWT2v8tXYchMSEf
iNP7c0SFej/I9UNd35e5ilipFAv1rLYeM3pMOB53t86GqoUrNWRr0C9G6Ru8uorV
vtJVtxwwPDZ8ZKIkPJ+IzNGGgPApC7YekAzk94zavPlY3VoNN7R7h0/GoQxXJzcc
Y56h60UI37n5QCGkYEYTuHz4r5ZmYOC+9WEf/2Wb2Il9v7KBrHAL6V752W1FyxXB
nYVeluVhpcFBBIZ4Mq9HQtbFCimvEl+FxanwM0yjKZ/HHjr9HGUM8Ssbt9FzNfKS
fv+qJXtAagzHoLkhTpGqfBNyQ5I6ZQeyjG6BcwbXfI/T+vrGxQdRLiYpjy017Txq
paOCsdQQ1ZBiSUBlMFk44M1siQ6AbRw5IYDDhYRy0e1HuQL9ma8n454NGxpyQzMG
vl+XQirl+rgf1JpqTqiu2WCA1xj7eYLsQsX4CgSjez9LSg9GLlcy6YMPU75Py4UV
gjXDX/Dw0CIayYf31cusss8XCX7Pc0+vI2a8lzGoTBQIBpDdDbvMSsJnot3+od9s
z5+cjL2b0i1dkSEV8nBi9urJnDgaBLYr1Q1I2KsbqrMa5rMArlwbjepwGgrtp24I
PcUTgmxKGCNoZBfH5G2GXYlron2HcfdUKQ6Sv81jdtxcK5ZTrMlnjdy7zM2aEB1E
jlDjTIaPl1pTPDZpj4uheqBviD87dL/bTG+mlkgeYGChcBQsfoC1DOpLX3AEWP+E
bYsJjzEd/Cfg6B24J3GFyr/MBbnaqMPlMjr6gW5DO2pHfFP9PK2HuLV2qLUtYkDX
Xt5urXLkAYjHydVT2NtndqJs9wh8B3XS/7OQv1PuKLI1a39t5y8lXU+OYgqzds0r
NrZpzhj3IbwyXE7pdjYCiFYWGeaC2msffLF/OK2+k+IKXjWsIuNZl0X9484JiDgC
Wb8wkx1p5Cg/c2cTyP4haRIj9x5gVTNOVJCIHKoLhezSXoEHRG5SNt4Zi+jQFC0k
jFdMSW1OoFdGqpHpTZ/LVeBOnBLzYsdYrMXSyNtDwF8LCNkOWQwcsn/gllrTAKfQ
M21c2mdwVULG0ZQktTHkYzYqKxT5YmSL9SFNBJM4h1byNsagWXtv/GkAWe5mZH+v
33BCL2q3HURXuAZihh1lcpL9/iC/E67eKMTILHzDLpWKftn/2PNTgD8S/O9ocPfT
mgw6BfkXkhgnG9WlpHDJmDus+KSxcDeu5zlHkOrGPNDvox/fD3NHW1D734SOikFH
Yj6PmjuFkU3PQO5mnMkbk6GN6AwHI+80w7jXT56nksr5Jr+McVojgD4bFr8fP5P1
aK1zS7TVRXpvTKSQ0glTtbpi4T+eLir2OQHGXNNarHSRRbLC0bDa5cX3IhlLcEH/
xd9vOnbBPFt73LXZVJ+CCqi6XmWvPsOXERIIkyxnUiYE/m1oU0gWlZCxOG2kEERb
4dI6OHbYyeLisq/4ZtxuF2M0kQGY4TBGAVBgO3aSvFIMjQtgwwoEDnNOItxcRgoB
YkXgSQd5J/lcB/cqLfgnj0gLfCNd8Vne+OToB6yu7a0/HF5dZhgMKFKIPSyKkvRB
WjMk2WDeYvQ5mpWXxJcU50+N3+elbtY+fswPMAdVJLt7HJ1d42q4PYs9R/2LKbXd
Th45XVf4BiSISM3N4crFqO56ntvkcPeolzm9M86gDTaqFIXYB4StJwQwDy2SvhHO
S+ahRWuj4rBWDR05W0VZ46NiGEprUU2HSk7IydgM314SiZ7BC1R6lKsq5eZDSpu/
LOcrVU7+1DkesjrM3WkvgrwlDwsaWjrpv7QE7ckvGtsdpBWZfi/avqo/M1eV0N3U
IwN7HUjKPJuMX96NGqVV5gectETCWceT9qsDCzdBGuFdYhOi2HwoyVln1h7oPNqM
i9l8b8dbiP6WQ/Pn4hPgxiVChgphfG+AogVA5QXYVOjd3qWhrcMxRCZ2ak1A/vTm
U3eATDYEaTtl3Kl/TiCInOeY62TN/BNAvP+4gwkI0nm4EPrVV17CQvxbgzKzMgqg
GwymoUYbVDko0IX1139XicoYzN/jG4yXg9j777iTxzARZGMZR5i+IMnv7CL8RtnQ
NNsW28fJ92OfY5pX/9sIz5b96sY5woNmxBjiNmIE8drEBGOuaD7p0jQqxXHVHVVt
hpRJVTYblNL1o2xdbYmzdmDDkhADWjxU9Rjm2r0ack5AKsC49pVCxF1ntLTBQIt2
ho8EewX4sH0HJowG8jjaiz9eXcwBZaf9HfzI9a3Cnm64mnO1WVyYMkwcZJr5qMPH
`protect END_PROTECTED
