`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
tVQSwlx6V83WnkFi6KLS+c3ftN3kTF9uHdQf9uqTzPAQlO8xClHD9A2DLXEpXSoP
NRqZXCIIcVVxdvj1f1M4g5sZQw8CgGkUHEdfb2vBKr0lCP7HMeY0eNVuw8cLm2bT
3/LWGi93Xz79J1dSkg3CI2LeSM0Ipp/Voge09qtwi6PvvvHA4BcwlWM3iZfSMlWg
QOOsvpPJmV7E6GshUrEThaGjZKbY1G4/5yr47gKqhI43OIoA+7PQmXsShHV10jPK
dXT2Xrpu2kHaUrfi5yJS6rxSyCg/5XM3sjQz8Mdcs8LRoNBDxYKD0lkVKEUMAtda
JuWXpq6WXNFHYfFtGUEW+I6E4gjb71EeWiRAks1n4dkbIZKQD+hbSq9J2DNSedP+
aHIM9wTnz6ZR5WXtFx0WQrfl6dFwJNcc5jEGGN6td8NSMGdxsUJniSulwxtw0yRI
e6ezOVeLVWQjXFhapBOfSqnVOmDazd3DDAlHJHyrkqw1wkgj7aRvbQ4oWG9WFlvy
424yh7W+5fAQeLX5s98Io4r9WJM27IU6kF16AsLCsC09LgA4Rp2easKukQyARQCy
f/25ux6DUsr5MDtT2XqlfchcWbuSPqFAFU/JyLiU7q9+bPj8GSUNn3XT14YV+KK7
ynXUu4eR7jpnVXWYxjtbH1/qiMDvRP0CucRWAbAX8wftQrmQWuz/CVSUTFI6LCTV
UtqzQTeKGoIA7qJ2igYljzfXxYzTUjXj/dVl0tmy9dFCGUj6OEbVCfaHMgmut7EG
UjNgGJ/0N9sK2nQtu37pSFOUuifYiR12VrLFJVoNokMMr5SLww5oDOlsg5vlznL6
XxKU7iSG55A0+XvUAS/kZkfc3zgn6LwUbu0vJdBvYF5hstSxE0BcUVm38hkpn9vt
nacMhFzz86H+WGRYUvcZGQDhLZwLiZo00d3JfcGlVEO/LKrOohlQnfIUVNz3SGgz
3TEVlsxCDyIDJcla99cbDi8imHDgO9ZJssWq/LCO8M1wwAYcMurKcVt77hXa9PN9
iiXjvzOfwDtWqzD8kQ5Y+Wy+rh1O0+E0K9mRHV6hh6QLgKw2qOtOJyqMJUseI3II
CtVrUnBcngCYcSAPZY+aeBKw413nZAd6ZKKs7nnVPQ8MW54Q5nDQFe1+qTa+0uMT
jWmAAQHm+nrT/wiwVpJ1e6J3LIZpYL7ScucAifqAEJELdzxzgCX9EGkGp9/qliMk
HoyhA2OEJ+94GvReFYhixU6Us/YTkK8xNQUP/4Ta6LdWN3+OA+YowSW4wMZTgBxu
mINX5ClTFWPuBB0MqQhLgr9tTILduc81EQs8PgU8w9mk6rTwM7+fe2PdYE0Aw9Vl
ZOcsauAy7a+5+/ElAtEiPz8UaXK1Ok1MWdfPVXt/Bshiy/ZHCSs535mkgPDlGaCh
yj9rXdwd1J8VN6k6gI1GD8VqqwpKkODhWJSJ4yKO+ZWN8ne0Adv40pu5KEHZilHp
fm4afnsGXq5CRjXIsgdH7BoH4ycGb9VSQRuV2vLa3yftR+VuWD+AyqaOJZv1EDKV
C6xalLFS8FTB0PVqiADYN+KhkW5bu41/64iQ2l5mS5rx8K/lg0hgdW4yc0zh35p9
GsMQUHMhl/Jz81qJa/6plQxRJiGFiR+AIWIHlG6M3pcHAIMMscHixX0yW+RRXeBQ
CbiPiMeIIM9I0dAvafNkkqLhDZIwWy0DfWck5MEbjQAN/ItjVmjH4mLIKlvZNc0C
qiA+2wDwklYadSJK1XYzWyj8Utyi5SFQQ6ACbTt8xiaeOMyoQZo+K0opECOnVTlS
arZEKguoCtQJiQ1srmvjKFNGQa+rK5DodMX2NNnQutuXZjJxRNSzQ5moddFsppRz
SBqY+W1TV6vyOokgDvkcVox/w6qtm2h4bcOkjC/HizVdjhPzmw4ILObRv40919wO
7tEdmL192QNW6/J/naB2O4SXVTNPWcBtKvpJOGATNGpPAw6Y15fH2QUCvTxwvia8
2BmNo9wOYgdwVujCyGryTB4CFuoabAmEGIbiK6R2xDHf0w2ojsxjqkHWM5GEq8eA
PG3OvNRK78fjBRTVseKYBMNksg98GzSLbzhgjIRGhm39AmVa8fxJwaipwBim0b4+
G+vp0V8St3gjWdYnJ7bn+UpEmadu/PLAj7gkLoxTVNmitdPG9k7T9d+uerlcKqyq
bnpB4kXS+5M0jmPnDHvUxQCuUsQPXsQV7skCZkzYMFE=
`protect END_PROTECTED
