`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G/qKWblOL/lQW7fF9LTzeV36d64aqO+RgFsb3Am0znOg1o6SeBV9OSvbAVImXZaJ
PiKEJtXTPRT8UfQzX7wclHKTBYGix+YV1fA5g172qISKedSdSwMwY+7WOmK2rtbA
a5MTiei50+f8xej95HOrIhl4h1UIW4y7BMPy1ZY77549yI3nbX/s7b0LXmk4cXU1
3S66m61mX3vBo6bHUpfqTA4KR46/S7VdeagryvwfYBkTHAOUN1rxg0GSJVorATqm
f2yn0eJofm5ZzGrXurHyEHcVHIQh7e1EF6bF3jpVsqe2Pjt122/vC+8JoD0ljL5U
q/KLFLlMTqmMWdProODHLvUrv2KLD7yMLVWRsF1stmFvWYvy+Se68ya4PsRotCbl
qmwmE33uybY0JQ2PignLqTqGrcluwfgnmb3N7UW81ooc57JvvMtdtBduk1UbwpuQ
/cOah4ZZuqVH82gRqxvXX+MaYdQUB/XaKnnR37sFNETrGcn85bCamr0SXF2zZGyX
VP5+Go1IaTWOus8uY/hMZhvGtJjs1vBTc+2PS3DmOEeG770UQbN+RvMofzPqa38p
ON9lUo2A8yPBqKXYmK/hdkH/rcooHD+Pus4Qo5EV9M2kuRuaF1KmEfHV0UAqbfUR
0AsOak3tAB6lhp3MrNpCZcimrNgnI+96iTNbM3g6MYRkCC7D85gdio+x7DM5V2bT
aOOOpDz8HC8uxK8MupJFFaQlE9bNvtHWJTDKNmAFXwfhGMYsMlDwAnTyA9S8r3aU
CVPewB+zdT/afFSibRbQFHIrgg36JD7G/9ANad5jzGovJzIgGCTBcdsVS/LxSmZc
qghenpBDs5KSjkB7F/s8o64pOpUZGgh64FGCKIEpdtb6B85mjId5Or33hI1iU09w
xVgP5ZaMb00flbOvLPD60sU58UGwIa8G7Wz2tLLOzUufdwvf9x3DwNwV2Nm1ThQh
HRYrNH3AfPthbymusAbMio1/8Ixlxcf4YSImNfcs1y8XLVX9/FLjmYtZaXMYgDi4
SBoFgciKeDP1bBBZBurfD67NNthn/hTiZf2FXIbYTWHWal4bq7VcpHrLOAj/rgQT
q0qgKo1AwWy960j23Ct00uNZEjZTLfV2vJ3y9Zqw2jxxtmeOL2qMjJvyninWQHp4
UvUbobP9iz6MmFkwKQ9GrBvUmfMBSZpwPwbH+lPB2vtkxd/Q/O5lNCQ2ZR5myfNy
gwkEwBGZK+N3YM1JPgBA1vF/mmvKH2eLMnepGDEh6mUv00EEzxvBsm1hEZXXmvAk
heSBOlIPksLFFGnKSN4D2zYhFQc0Mg7WuExWK7DKo22/hGLnWnPy1ZnGF4MoinTe
9HcD+D8d0nBtA1BkMut46kEVfRW6bCkLf0W/SrZWgIolNA4zkos9OQF0e1l0kuQT
vXwREAWiAXSub2c8sre49N/hAYcdo9z5Xu9ZY1eLCW+YyP6QXiNRBN7IA/itch5N
SgitotHRdVUJ63ESOXze5gKY4hkUJpyJ7TFtGTxT33OxqVHxM+DKLhNOcrzUGSw/
UUGPRdEZ6P4lwNyPjyPr4UavzojShl9Gafs4rqYNPdxALe4UDmI6qfzTAI3bhDlF
BL3/PLyLTYE3L07+d2ullhoO+g+kCCdfK0cDJusyyx7geLWQY1b0TKabue/XeUOH
MkXENb9BYom6xY2BHPa298PTTFLwRMDthBHTqaGhx/ktui2th05ImLAVArXimfj2
3xoi0Ome3dQSoIyXCXNkU5Z+OZbSH/KcIAdx3U8nvlVbWvy8KC8Dnkq4gmNGZpG8
XQCXo9rczRHGzBMwrj7LNMIAoxSDs65dkUG9ssp7P7ZvTmzAMS0KYZLHCFdRTtAv
E6QCHKotkKU1Z3JgEU1GDF9qmQ/gYrZkeaoiweoj1Q7EB5Hzd8UPykx1crY6QZ0u
Miyl8JARFbjSJghxhzDn3M6KoFNjo/+jdrG8+Jqni7pNjY0wrFzf/1mmTj8oPiej
7iDYSQHLTGT6oYU5VWI5qBoDAEiZRUh1ixfDuQKh9d1dXC/RHFkrzsIDoUCnDk1/
MMfNaZNk9BjSJqnGRLCDrP4Gu5yQXF0J0b6SI4pe4aNv6Sfpm69Xu2P4cnBtzJZn
AMLZmrxbPJNr7E6r0fMG1Ts/ppngLsuK9SYwi0mYYUA6AHxRHxiC16r3Ygqg1iqO
2rlIgHkBd8jWYwpNPbBhtVzFx0gNOmEfiCpmKlapxVv99+ugu6hnn5rz64fs+KQG
cl5C7T/6+MB4fbOdevdA9424ofRseL5dqMuCaPY4Xp28xI9DlJaSjFxZqVAQD6E2
w9oDfYDAs3wcxIQOPd5QmRkaasbFpmXO7g6vqZsyP9vBNM3XH0fgiKvXrFky+nKJ
n6xN51lvcbFrP2ENMh63aODydeBpIJujEsBNsozH7qfB2tzz/2SvOT1tTbAq3Mw6
ugh9wD7Bb6iOE3alhDx65pZLVVZlKBYa/77c9u6wL7CBmQrSv9DNO9FzR0p/+qdf
eBNbSySV+4tj+Y57visZralfCDLgJ4mx43W7gAsmqOFi7pz1Y4K6AqMC37Qu1QMR
xNA5riyeHdsrFPXy6v9KUTf0rHTU0KV/Odrxfw0jbVtnrztecWjG7kHQ2qqZ0mLg
gvufXzV7efBpNpygVcURHVqz8SH2PI+mTxv0VLgyKMfljFSNRkNgAJixjXZQzCrw
L7llzzHmmYD11vo+crRRV29DAPcHh+REoPjbjugeOCFCENE+mujR6YDnv3gabzik
04mHXuFdy0LEhNIWVcVj/gdqZw+u9cBJ+FAnex1VPApuL9NVkFVVr7nOp5vg2G7v
hgbT0v7QKqIj6N8nDHdQk1jrL/CELaIC+hDAAMSikIll4DLn8uF5ySrqMnPEdUcQ
QJb0GXhXU3H0yT2i0ytzwx48dKk4OxuKF29C9QvHfN7rgxKyiMfADSf+ptfBHr6/
t3Y/czUM14E/NwgOsnKm9gZnLnhi9IgPbE2koKGHf18gfpGcJY+iv7AeDLqYV9ss
EjThUD2ASix11iifgG3VkUfMFYki9B3YHtI4jOKmT1vDEw9mIJ+7EXqp0dTRA04R
nhEqjzTDxK3DGFbupyobpk6QXENCgPe8DrnbFIEfHVIWLtjGYyiVMC2XsedvVv89
SfdwRw85+5QSOa41+crUvFyhOVDgazOajhGmLuvpArqpC05D1l0lvThURKyDesVq
z2NkZTkKc+sEbPei+o/YiXO3o50HkKMkRnj7DAurfTlGsoyF+OGMJQ5S+SBEEvYD
IhF5BheHnwcj3TQDuXrydkLTvsalXTJmiQWohqRtrtB0MRF0hygm19XaUXJLYnOg
M0xjkXZwpcCDyC4qeFvaiNgiqLxLv2JqxTJBHdR0YlVrH8j85mwqW0MMRuc88o94
5c8Zzp2ooJz4pVh5Ib7JJKfqzP8P2foJFh3Y7fjIpBrIExrZccma+YRJ+8+0e71I
foU0EeWRPYOHnDCO4RKEgwxaL+028DyYmXv11g7dDe/GYutsela+2JPuzrJ8c0ek
jvRcCJcskvUr6TEoZRiNOiwyS80w7dr9jqBubSsxMllvTzunq/L//c+WyvMVrMsC
mbfqM/u5WUQX1NGocu6Grymab/XZnNE58D6/Z3Fj55Ve/VqmUKfpWveoLujAN7if
xagdbmidbr+ESHv6m4SjOEknclPDDzRQj6fXAGJ0+kvZSLbw4/P5OKnpmlbDy6O4
qLnFcb9Q+K6gK1a+OU7XL5d8QmXDV+0PAv/GsZR0TydWZ4f68Yf4OEXAH3+pmFBB
Mx+jUPxVg0yEuuQ8r1yjeQx048Iq8jKJIW/180r77b5aw0s7mOXs/7XlZ/Q/1au6
071ZuF2HM6y+on5PoxdihVwWA+JF1fSAppCCW54aaeXaqIcCbM0sVyhniMBehwdR
PFjgqQNZzsyoG3jX6LNB4T9ahHvYx31c7r0YXIVKZbPnWywFaFC58n81sj9/XVGL
VewA1uC+vyxOVkxeFXCvs2FJd0ep6wI0EuKnVDTWHM3pYOWzbe6AfS232cCy74Pz
N8Y2mhL0qBOQ+ZAXZJwbgJA90I+v5ndQ6wmF+G2D7LfVUZMGnOz3ZnNKZbdvOnHC
MRIPCN6Iynp77WuvnfcZF6+OVNhkoabBr8AaV8n3Y1qDPM0vEmEbU9OZT+ZomxYI
cVR1IO3TlWkvdpTmkAEAH4X0UZ4A1Eg836jNlxWq3mK0r2a+7Qa3+YNcKNiomf5v
bhj1gfHzzoPFeB5s98shssQWpPxu6IxWYxLCeetZMOT5Q2HyoIN6p/zqvxC1Lu5G
VBAsbgN3IyTCBVJD8jzvOQftj/NDqlMSeMWgb12MZ3KFd6DFKqSDSAZbSFI1GU1e
xJHmrpM7M+6Y7VleFEbxm9DVvtogpf0g0P2aLfG+j8ZTNEbKVSV0h++Nm/VJ3x4b
tuQbNcLMLQMhPdg+m4YsmgFIUcMG1ioD8nlIhpyB/0/40t9pNVSFPAb03doCNovO
fK35AJ+6ZIlhTVqfQ2m5cW60rpZHqraqFefpoJ5WvKyu7+XmHxreedQgIjwgQBaD
0ZcOhKUYXBsZ7smYW5qTmROoks7QE7tsMhfIrRf5LjE=
`protect END_PROTECTED
