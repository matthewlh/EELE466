`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
mzKhjuOqO1LivUms6Kdxv5YoIH36BHb9tNpEi1hfWuT8AU5eFM0/vSKc6ofp651D
TbbouttqTiCseUszDROitDwkeJyb7WoScxpOhM0+yDHUVV2zDkQj++fSDnZyQutG
wLAdBxoplPvakxUTBT9vztLFm/mX3aPygllJIqeSYytm5Zy0KjlRNxMCDTyfCbuo
gTCcNNmTC7KWLBsu13lj3Z55V/qdQsGSFyZdvtZ4EnR6fya07d0XX2if2mG8Tu6l
qvm07xuRRE1rZJAJuI/6al222o1Q3cbfOl8DB043YM4mj0GwRZQKPRY9u2p+upBA
62DRWsF0e+efi8mnKZFgFDTg7hL5CJBADbeSOHShb5HFMc4Ep/l8dx/3KShfZCX/
GfSe8pE96pBXjfAlupdRbbWrGsRsQM58xJJnsf9T3mI=
`protect END_PROTECTED
