`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
85O+jT/8Tnn246c9i5JGS5t3vAsOxLPcrPZWux8xiq/GlN+ENa3AXMZsrB8YMD21
ejRkPgZ3p/Q8/k6VAQlQznDvsdU2hwP8CnV11fy+OLF5sxre6t3wGgOoRYdaQYL2
7OYQnJCxXbuEpx4ryWWKD2bX2d9JA2MkOe1wu46STXwFtUzKWGC6irtFD2+/f81V
Ass5WtvEcb7ZXEOxFFmzC1RYa7L+/mrPXYsQ/JDymUgDnjlZ0YKzniYFeThMRTPk
CeZiafdlo/m1/2VysKmH5GCcPu5SGXw/hDoegkIADj7Xhk/f8thP0pDzeolHhRD8
U9iQtBaLtgoCFF25UFmn6LJI2HpQ8AFfxfPSsUND++vdQMBQ/S7gB0TgiG5OyG8o
QH9zBjnfNid6eqpDIS8L0C00fSNL7sZzbFSSPZ0LChXnMktLxb8vcT/PweS/f7YL
Cd31uH2+42P4mX+aI3phhW/FLQKHaNUr8mPF5lZOMGmJ4xOHmmV/MwWK6Emz9ARL
7jwxA4dgT6NyUmjHrax4PD1sMeDYJzpmfoH0zsS2N1gW043TNAt+IuRVnDmn01FX
EcEzcLN99bn9lfmP3WvEnjyAOhRVRgo+4kAoUK7lPOhv9NQ1FnSsulRZA85QkcPf
uTQZnliPK/cnjFMpJLthNzKFKjnFprD7b5GW4KMGuRIH6/aJ46Kvyq2ylSTNCmUT
0eG+bADgFGzVGTXmlBVCqv+Oyi3AAgAsg+WBq0dn2otmOajHk6KR9mes57vvfFAC
IHrbnfKPUsIEWRmHhma7aSUmrAlRvwfT/wXzndK46TBHLZFsiS7ZllhkpCaSGPFK
R8GOj4OZayzGUspzwuaUs/wy4eHnn+qXwytHfYNeSAwTVaIHejyseigLtfH2hZ8U
W+yeTEpz/3zkndpzbnZYNGT83uoEg/B3TOTyvhOPVogOzXVTKRWRC0sMEWLCzF/+
JYHMNGXvTgsX+xMz5ytAIRa9gPVALdRjlzHJqwzo7YNRqeQbctcJfLR9NFeSpoXJ
3PGoL3nVbmEqh7nZBZn8LF4uhLndpWHZJK66O97pP28fvELBN2GGthO8ioIVCZPD
YNWDyYLeSHQwN8r8L8R1nxTo0lCgYiaStO0suS0Q6HOAJJ3c8Sja3DSZyQyPtaAX
GWINy60KY/wLdyTxbth7HLqyJWUNFDD2fvR96i11CPBoNlsuniFXbT8YzVjubtHm
Cmug8IUMjowU/OB5WOMKU9nIxFI8HxhhqXSBym8A1yLp0SC6/czcP37wLcRdm/yj
uyaGyW/m1nuCGWpyQ8Bqj1fE9N1kJKwScTouscBRnTyAhmYlnbC7FmYHafAgSbD9
AnLCO6GTrV0FgCELmmA9w1LbrdENrrNvTwhys+md/NgdWzeKBwQodOIZn0fvuqdf
o9Y1l0EiJiW6cUR4GOs49+Ug9y1Fv5DIpl49mADJ9KYdGW9Ss/rTeLb11G0augN9
AmUHtUH49Q5eSyGGWapZE1YPksTnlA0T1F99t4YUexkQdHYwPrBzzXZlMwxdozal
YkaO/QtHB9JBVjeF1Y5/IUrlhDR1g69AWzyjj4fX9tI+pBvLbnuMvc3ABtE1zTCT
5poYgtdXteAwqzFMl4jzqweaallW7IHrwFEqqomaz6Rf2v3St7fxk3c1xS9Bb5jE
6w4VVLwarOpI+r8tlxFd18eTh2OtqooYjJ3z0/D4+USkpMM9Y3K07IkVeD4Wq81R
s2sOYilZ2PSITbAT62Y14bGtFar+D+Ojnag5IwCgogk7Xz1uQ/FSqQUaDNIWrKWW
3ORmqs/CC7qfAv/ffrtmxocnThnjFXwDNMloGuoMvZ2OWg1j4p3pfkWxKI/YsVud
z9iIc0uUIoxjRf9tOpmp/n0HDmlc0dFVKnicDIlFpchIUChWp7OgIK5BytenihC9
GGf7VpKqn78k688E20ZKEq8oWPh1M9f3WiKnOA4r6aFT6Y5jCHrsxg55KT+vhuhf
VwnnCrpsupfpXNzmkj8bE91EqWjUfzG+zzLGoHB4OTTCat6URUUIz6qRGPzXpBbn
/BCKuTunHW2l62gJ7blEqv3gYTDakpvpCBaWIy/jM7KMjB9B7FKQ6wJk4amHU5nf
Ntww3bTYkXXC79/FfMbccSXC7BLThCsBA2iIN6SWy+GjnzWZ2PUTNCc7aPOm0vgS
tuFYdZr13L3d+CqukFjATC3Z6bMBCK0CbqR2i8J/JkAYXwt1VjmDAIAzc+bm1DKO
lTHtZlhF/H4r56WlUooTRSTyeZn6VbcvJDSwFFTnHUoPSdb0AbUDcAZE4Cf4qGzr
5ar3HubZHRvQlf53XPEUYMNuq7gSsl7iRqsgAFnzS1qu7ww8UxJTcEz/sZX5IjbP
624sxN80Fr/W0Xjt0tvUVS6uPY0ZhEXxiLUhSwNo5wQOGl4Kmh3stubXFUnN/y32
pBFd/UBWSwqsvF9IKs8Auofx0Ra4LlSxsQh0AxNYrTHx1y1zCzrxFfmWvHugvkGW
t4hKdrGi3nAVcdnc2N2BdOwjeH6iQxp90GZtMSO3XrqIq8wpDtoA2LNen5fsfONa
4Bl01EMoUyz2JKRTjh/2+c7pNaIGu2V50ISh1h0j4jPaRxwXNsV5zGMTUrZCbB4J
zmzlzkHUei/x1nx0N6sFLB2a+Aq67CCgLgUtiR4YGReSWxhUZrKfIhFJyhj48gp7
IX2+i5+t39AfUQrQfAsLUQJ5rOB03IKp+V0/ViaXn/zoTL3H45qnxcgEQb3MzqnV
DKlXXVI2PNuPFohNjtwYEEM0F5Y+1z1W+/viVLjH/PIQuKY/kYTJaj8CUx3BozRe
cyFsfi/h5rcgi2B/adQbJOfdaRImtKovfvAjPuO2mwFsh/GCTsd76A4/JxaiF35G
pAjvMGZh/3FYzcdlRNhQlI8v4G82KdbaOxnVpQ4psY7YA2gbKkwagm8AiOnSeeLY
+WXwfotGV8xDtbmzbT4UBZP+XW8ttJV18jw8BvcjRLyvHnNbmi9aggEtn3Uy4cYI
5Gysxilf1yM+huPM3WsztrHgkd/dHGOOszxnuVLo8m79cTPkBVuiq3K4sYmx3ccV
0ChvAQz/pKBhR+TNzSXKIUvHmy68Uj7QwtexgSh8aH8z9kvuzp28nk9/dqHc8rdE
MBxSkfxmpz401vNbctvpw8DXUBM5HYaQaELvVaz57ELFXJoik3BjgB/fAbnDHxUl
ChrC10POg+R06qojfBgGG9fljTc9yaDMO5AUYuErBpOXd9qFnsi5Oj4EeJjdH861
kGR4StgNR7emAJzwZRJvCJH4oiXKPqEM3Cpotc4pIY1fW2wp3cfurnBDHIAnqlIo
hAjALZ9z1ISm7+FVAdCIwozg81BLzppwI5xZ8Ki7TvTxnyG5ActnleLFViGmbITk
iRyZToqBe2eJng6jp+F9y5fNSEU+LXb5HqBmi8usQfwIGUKPTGLtZ3WSxF7Qu4aP
DOJMxLqLk02y9akOXf3a5DEkndZakUyPK/cQITYCma1SCWHw/dpKgiScgswouZBJ
dQQltZGQrLprc/sFPBwGUOjQv894MAxsHUvdESSnK5E0QjQ7iePwR6sZfJCNOQ6T
jT6P/pTQPjOAmG0GIvst0+JPWBG402AOBJvXczs+aAP64SXzU76vdcTs/HbHXjsK
gHyk1M4euXsB64XLaRUD1RG12TluaLcKwyMijIUEy38zR5MruKJFs/BlDKD1QUbU
shUHixPsY8PxEzBTSsXqdgDlDrN5OOwPg9eClnV80VBUXXJNUNe1iHrP4ZH9NV+9
g7V6O/zWIWEjLCpJuZ0f66me1qHfCDnvmCSAfRUY4gnRXIjBIM/7/PuRiWrUDiaL
RHAx5NBECX17FmFJsBhSVDxwYxOJoKxRdQZQO6EEfSweTUHO5bHAVbDo+cUjj+0g
dlP4e7ipkQtoqHA5u+wA5tJIuY3YAdxd7GPwfXuy2Z5ak50Ig79Eut0EW2Yu35Ao
79D+Z5pRQdCaSFJJ7qCNfMACMtycfBDJpLZs+sQH2l86kcFROp4sLS2oEqz/8WiG
dFysZ2hd2mFLw0kCRRCmGjbQUG+Okoxny+qpt7h4WIGSTmtj9ocm5mm4IpSGZYVr
eLWLBOZSadpToSrn0/JEvq6WBHMBgNEJWVL6BRZ/G+lqvjSpJhcr76uZP39UeKNW
9MfqPGz2nJiMXkwg8Vq9f+X1AE7z0fUUZbR2rMlcUAODAa0HBIrf0GRbaeyHA+Yp
J4kSmsazAzIIiivQyk8wZNIbJPKCrhBjycOxgXjMRLX/bTSr1nAEddhfBKfUwOkh
zg4ERE3f1Pc9616GGMhI1GDV93cUKe1VIb7RB5YfIBZ/CW8u7f/DCAHEPiw5vKYT
IlE9ho3OjVcyodO3TwYWW0Owsm19MAu4wCMtPI2/eB+E4wOSzkIQDW+MjVOX1AkB
FuzgRROTO7ix648XZhmN61HWjctQEVJP/DbILkr1W921I05i5wxNDlUhVJUncszl
JE0soHFRbgt6O6AWkPawJ3EG8eDpuwCnN9qWtlBTmMqEeHmM1hJjoeC8EJ96pxUq
CxdELyhVap91EWnhXrysJHUnXQv9kP+PZ2qgYlBVNy1u7uuSligFaeOUfS1wAeoi
HCnPgqiF5GEUmwZIzhoeNhR2Dh/doKbJQ4pk8J3yzF40Jr+PVoO7fzIVP2HAbbMp
0/hTx+aIvLOOUHyjLP4tI5zAsyQVdVXVg6Rprll/kLYuW8H4+xHHywbNhzRMMwC3
Y3nxaO+E8w3/MJblb29paXmBeGAg2PiS9E/5MvO4mmMxhuZzMUZ9MEi1ev3Bu+hL
c9ytA/z1mk1OaPgkh42akOd7kXuW8Gmh8p+VJbJfD/vQXhql4Opr4hl5lXv3Hqd7
RKuvHxzG1txzdaxDQwvAlRzrejlPzmIExXG+uwZbMmNyCNe/oCAHgUSUA0bMRtjw
aayBq4l6QVYWnC5mWw/O5a8Ryd4W5yRxswSRXMsAZDcU2+mFcK44EM3RN8kLcrJ2
gb2PVTzfaSO7WGh+3AIRpdR2piSroh4uuUk2JAx1IOrjF1DkQezS4koWfHE2LVqc
Gu0iO9sqJoVGt2RQzfRYi81/l8+pH/LbuH9ph1/5uKcvib0AKxqPOxiq+lO9sIg5
lkM+9BZFLgZKDzNBzwGTFR0H8thTY8ekKYATrRMTd0e5W/xCoLZ2G8ZbiaKOlJb+
wz/f/H+67hEkYT74vzkltR5zkQzfZm/5X+mHcVPy1EZGle8I4R4XPVSEt81BXU6t
jM0KcC2tVRJ3pg5n5lXTZecdQx4iqeAIkjfn+2jlqVA1wJVEWxwdDldLEPTcF0fR
N8PvDRol0m7gPI6G5CAbnR7hBil4IKuKdaU3IuiIqdIPrGdThV1Aud5Ajw+HL6TR
LgCvcK2CEhA4ZrQ34EQD6QjJ4OFxWPHmmzBPhqYRcgj4f69ljukn8ctEblVmTlcp
EmWM8fgAMleND6X5JC3C0K6wBE71rFS4JIRkXs4Zp2OYi9kiLXFO8sLZn40IXfjO
+cpiq2CYlLBcbaNhjcv69mQkErvPdDAWpiWUuzLq8NWnR+D6xiEqAGbSoLcAweHS
Wg07/mZOlkXG+8ZTVjyPNQ2etNsybfqaCkdSC70VHouD98nbFYTNX7xBkDVMMZKH
sQ/gaFUdaG0aI1CANjE4DI5yVEYUQO73tMe2N0bLPBHHkvgeqA7lGcOhGntBhNqq
aQKyGGiN4f8HbDCjPwb5zmsad5+Y4soScomle6I3bTtsFdvmBYmSx3J+RiWc3qFW
jDvSclMwtbbmanZl8gMg7YFrVzC7HXwkXUFem2R/Bm7PUCjGD8Pnq4sS0O3EvplS
yJYjB7YIdmXfBOUOVnPvhC1B50P8N+rU9k4Wmjfojr4Bi5bXEGDxbfYe4jWvCnVx
uKAB9apSIeaO22Uxz0ti987UnRQdoIxxADmxFYDMwrH0JXPuG/ci2CrtcbwbROgV
TqUIhcvGgY+bmTJl9CPNaeZWJbkxv8SLFZVMUZMQ0b+NIwCsCwpR4zYOG46OkvV0
hP3dIBAa/xCxLVOA5ozEMqrs3hH6PySrqv0dr+fHKWbpi59HAcEWG3+5njJKxMRC
COELd0LqoIynNrQLgqswRkfL0PfjxNgWvK+DwX8K07/dUjgSMDssTOS4pdgFck/Y
bl1dp+T+6YK722BofiNB8JBfg6FTuGRibSoO6c0NYNvNNjoardH50hWdQTfNLNwa
eTUpPLK/xXD+WTcuvPRynhH6VrIIkdD25gnJJxUuudhn3DiSjAD0rOs3/GAzPJe7
A54nEwpoD9zIUCbtlahDBn1t+icVWqPyJg2vtxvfDadP/XD7TAIWSbszOklHut6h
Pj3ZpZ1+xQHzM2NPq9E1W6tWP5mQq9gVoNdSwf92gXlEP/Q7INpwqCFfZT+CBU/0
hWz+VQgSDUe/zP/aeJ+gUt0rCogzTbcYqU5XHVZE6EaRXvMSHzGeqgUdnPQNEZEC
qSBzWv2LH/Rgx/omg5pKFdaD01ycBUHGcElNnvc7vVTK1igLOSkq6Nr41+FCuYaX
Hxw0upqkWEpZSGt5JVZdeVftLIBfMPqt5S2HPwVl7j5f205bJrrDd7KOO/mgP2Sk
osZ2Zd4oGrKGH+joiIwPRz0ytHCd909SPObwIrfEc5hkGug8zZgVl94A3XMF9u2G
UiQS4K2M/i2uHG3azyTlgQutZifsZ8RT2t6xI14UJBQTp86j4i3v7FZOPWthhudK
VzqCE1j8Nvgp8h/gEJLS/YSe8rDvH9rn9sLHG4icH/f3SOAOE2O73sYNcZsUpHRP
RAkbCME81MAviU4TLQXPZs0+SnFlV1FQpx0+Bbk8bwDa5jHt3yeSsvnxojFmnK6b
+gJTjxsmHvAwDV2jknFeMDwHyhOi/Dv39cxfuGOZXGQjebIb/3b/SJv5itzNsvO/
M8rapgAlPX2JOCEv4+kqBi72wdCBRV87NBByAeJM+Vu3I2zh+DJD2PTf2MbtuxnB
j4iOTGW8vuDvxVwXEv5XqLnT//YlXyISfty2JfiZfeQgN1ed6ooDetFi4munkcOB
6fCv5IjIFNO+kN3TuuFyB57txMlyXDL04Xca+OmKl41DInX02uKMFrVszjyE7Bk2
NZe3MJy2XQe1PPZtqR3jRg3wwRt3yjEEFPNPe3bBwciyIeoddJLuNqXHJiwR/xto
zcl66ncLwTy23E5L7XiYFOWIEsNUmSwI2Q5nkwnY+Ljg1RpRvIaujozsbSmyt29q
b6lzuH+bcO/BDD+6+mcmbIcJh+1lhDxJe8GyksYWEvFu0B8rCRqxXU9RcH9TILEi
X1CVLtA1P686B0z2h5/VQSEf5+zd1AitJZYOScMieyC2oM2IWwdwKIwPWTEyyuqz
RrEwfwY8QNt2aEyZgvrs4/1m1Ztcrv8p3qjJyE7YDPsJWgSt14ZMYK7hgQaaemdx
4cp2QOpsz7J04mVYXfLX3uESWat6prbahtRNrk/cX2ukeXU9kk3toGx4MASm4whR
kzZMP9RoNrTeg8nh1A2tbHs/vOwbzHg5L+AOlP3YcF4KRoM6vqwR5ksMsbtPsqf2
S3hbqD1Npl3x7MCS/AfX+70JjeIiqGbPIaeQoiDbXZMuqXUNFMHPkEUou1HcxhuF
WQefpXXYwRrX6F2zCxM3JWaGouFK79/8n/080qt0kMq+4n2e5/GW5LxzQbHAeUXZ
AQUVUffaVgBHbWZohQfNhp+qy6BHXhUvsJBZ3KDJsZge+wrUmUlqPER/+3VmQqw9
eR8Ku8Zkv3gALXi4fFLYfHVwkJGiIlGKtYj8zLP/XcxnDo/tPrzKcWsWLbG/9cDN
Ju0QCy2eqRN6f9N21PUTWnfNWhavvy7+pvkfmx1c4VO6Iac+tMdeTlUubfTcRd6P
3pqFXYbpyZ3lwp+dcf1UWTBaGYeYPXlXzBLeFl5iHYm2SpJe8a4HsUSFOf77zxSC
4fhvxg60BzA7DsU7wQbnVDbUTCfZYnGf9JiChdBMh+vQ1+HeA6dGM+dTEwdIe5rU
zhCwMlXF02YUG3H5K04Q3N8pt/C5KqfZZ54Q7UWtKHrfqYy7AHqmYrQSjALqcW5J
MUG2OOrei2A65N8oUbZ71v4GEljoz0oK6QPyR9mnuFxINTenOPNeL/zSYoo+qbmn
hQobwMntWZzfcc3kGiUil6et2bocpcmTRGBl5myr0eF9LuV6p35UoimzuRXkNqTD
qE5UQej/3k8G0v2c5jYYA7bRZP2SG8nya6AIc/ao1Rw1MxVZDicc51qGAX7EnR2q
HBMs598fdkYwLOdzFfAqZUmdbCuUHBTfbYclrdcuy+mDUWvcHnv+Nn0i7xML57+S
HFP/K1vGSAn4tEpC1ahw1L0oPhKvQq1WmyvhWER+53DNakz3NIPFQGEfBdulLGVe
8ZGy4QxH6+xd9dPTcoE/44YW+aR6spGZ5Ibi+F5y0SzRuwVEI+2gqTRoHbwRbwvW
YknWXFm6XDiY7sqCVhxEvTkPiXo/tjKNHxvKg0AOwLrpFjCZkR/4O8buDFCPVOjp
tQwzB1FEnOkLUYPN/+T/YcBvCpAl+S4pvwVp76Y8lHHl3AkstA9vmwfEIn448VMJ
kiaGicRAoNVQNR574zyfnaCvSgjM3Y8SlYUSBp35IzGbaMXb48CoGDi6tzpRlxGN
fP+tRQh53eZ2xekG1x1ZoX3a1BZq00JUiY+p8+bkZ7J7BbmUs70q8iYJ3XunRXFi
LTPe1/N3up9wkHeOmVToSaXpNtwGkvr/lvDSoP6D5XBdYylfWcKzaESwPdJCbgdj
1zuLqpl20VoO2fMs30saqSGXXlMNJXyoQelEjKFrJ403eUnklSJpvyY8c+yfNPV3
0d3Sum9TSWPIvhdjtwNuF0ug8ESrVcR3RGjdjxc8gHjfdI+nqBhUcAXWop2GKCJy
KswMuAD4qQW9muyWRQhiXtiGNtxdwYPVAvLxH8ZFK3+97m3OJBEInwhvlSCQoNuq
KEV75u1Nr56k+8IuuPYHEIvLe2/0z4HV2qgivMQHXusJc74qWUa1DFMedJ1lsDyI
1/pguLJ+vUgWnb/Nrn9gG7bD1x+GeKBm5j8mETyjI8UGT1YYEN9rn3vSwZNoAofU
P0uGohwG+RyvIgVwecwwHNdhiQxhk8vHVqxvJr7UT8FNlu+NhB8tfhtlgTG8jppR
DY5uNveGYVPKvIiO65wfsouPgvtAGSnKWI88S7p2yXr4xxdhoYYDBbavFVgRAmFI
NxRcD19SCc06iKvDK+UVS7BeCyY5dYVhwnN85JaI9dldL84INIDnn4EsP7NKFufH
MieZjqbGRN6GuZKrT2BqqGcAGGwaoYR2rxcNUYdr6+Hs9tL2r+F3fERj93uF8BWi
aMjpAPNPstQNKl80PBLLHH3ldG6I6nZop0d5XlX9oOkH194UZhk5GO9Q14TNJrRO
vqPpEVlZ6g/h4dekmh53S6zRtB5nftz3hbd+zcBLvILtflka5aI4ii6IEsrtDHkF
EXaY9MBizhaDwuda5pibrAHzrBLAQHAHAPnjxTDDzIE693TnhIJPN4Lvn0w4CwIe
x4qN/arbY7PTkCCw3pwHq6bw/EnW9NjYZYc7h4IHLezIUsNffutfW7ghXdNAnt+b
9ZfIqiOqAlTn49UWwXQzf3PPspvPYwCUCI8pqZJVH10kiN4iTavrS4tQSY7YRiBB
aM3uRWwzBEHjDVGN+EEn5Aba0MGzkzX9rVNNwyqiBYKVZNKIfx+VPqyvDPjbckvs
/WY/6NmSbEU5DnI9E3wDjNHlWEXdz/WqtbhLsrHUugDAyBgrqzungq8eooYaHLrv
k++WJRnC2aBlqMlI652gbE/nDoLElFV4K/usvpRW2PwjvysR+zNWVqs4B1I0ZPDT
r4Ugd6au62g9JC5yz7+SeV/IbG4qQzm1iecmuC1HDpskssqyAZsy84VqRbhQbLu3
3/XOlIb38ynaaA3lE66H3mxrTjVYZ+XUHUDU5oFMyruIOCy95nxhKLjLpm1f+NRy
anLMn45zIYosGyh/aG+F4IgLt5OIK0mJAw1s9Pei5llh39TZXr7FRlRoTS3BFq6A
k6H1MC/Jdci9L//2Awwf9tpY9xZd4VvqAEItvcP0w3v2Obcp8/tPvBGl+U5J+n6a
G9ikuzgb+Luc8FPzwwX8DI7XK97yFB9e7NeYLgG42ZJ5O3jXZ4d/djHd7Cj4w9Pn
HyId1SuQ3449q1qvTCl7EMXDx69lwxU5Be8/ChcyunfE093oICHBfNK2GYqkHfIV
3WGIy0QW2DL0A3w2/Q3mgiDw3oAUQ8JmhbseDrpYTORQnmheImfLM5pMN+XHRrX8
BDns3MLXewJr+UhxoUGDEOiihERyHsR18oDrbu+2I+plj14B7Xegj4fggi3CRsfm
mjKx5caH6A/Eqxqou3ihVZhF5AT+jvNwyJErnajASy97MHKggxuGFRDdHGSBSywQ
cxwpiP8jcrR/F4q/tdDbP0Agfp+G2OU2IMhEVocNRbjgYnYiqrV7fTbY6D8KKULw
GVgJISLCQH61a/tejIXykwdfqHQfI1ZawRFVUWsKGx0mTUIrkAzxH2Nf4FuKK/1z
F9Bnpb9mH7LeRxrQwaTdluy3EI7VgHm3GWAx8WN4uS11C2E+sH9tYA6Pbvylts0J
9hjAC+xxS0WZreMqs85ORGMCH9E1zCD0ZT6pNyzw1uS3bXJC7BUEwsX6x2pPvMM/
sjFY8Zqd0xQCBe2TlNqihV/uNVnusVJaueP5OTGbrrzB13LZywP83NzLJveoIls0
dRsrZOhCUEZAQ8rmwlO298g67rWyF9+BSQPw4SUEKGUYP1VsbOJoNHMV8HlJaXTr
w0zSdjdw6MrnYVBvhpecjXB7TfohcR2vCvjYyvWfHg0cNtT/ypeVEZwDc/Alnmn2
hKbWO7+c6Ew1Tdn6MfWB5pgp74cE2YkvkAJZGDohK8EBLSfFQ+VFqdMhe6TL+ANd
aqLp+XAscviOMViv/RgnHiDVcvI25/zh71XZ3mLaWp/jUpddMw8gmlFg7nMQvkYp
1oagdb+SEsJ8xFfUiD03sn2kZO3jA20ui8Sj0RV+6hcecYL880XSrmQOzrUJgf8U
Jljrs9Axt6lBe5Osu5WGt2lBPWla65QWyi6xqolyqw+R4dRs6R/UPZIepSV0CB2d
CGRtR2Ns3Kmjiw0daWY0o63unDHg4NKxgw/jhSe0ieA1Hh1sb3MUQbov/pI4vb+4
qkCK82cybOKXHLjMIBesk4aIGNbwOg2fKgcHVraQX8H4qsyJG6kVOCD/NdDIcBZ1
XaAW8UsGG88QsnD+Hm7p/6/Or16FiOsjt5OMrkufyBkrDywLtYVuLTiCbdcGLjpj
K4o48Fl0AZ8GL0S6z63FOA+1+BA/J4e0ACaOJtJe4xW056TwpOnBaYR97PwhCcKa
7zsEyxohY5VN2l/trWV5iyv4Zk8mfHtFGft0jrAY15izhnfJJ+TVINMTxx9gFJBT
MQLMgqahC+otgSnf5tMM6Bk2Yg27GEDnCIZQozS68UgeA0RpV/hatTqjzprdqh+H
30qXVEnRjvqO8e3IAPAej4P2eRS9yaTK/Dd4Wja56bf4htrOTQImRcibkUqiUJpu
sgTX+d09mQCjGz+kqMm9S7eTP5XsHCTmhrVF/Sm9EIhgmA7MSzbqWXaW6y2Gmpuo
8dpX5Xiw+5Hywr6dKtgczyVmxgwwK0Te2CValevFYPtQzUfq/7HskIpI1JepZNWF
PsqklGesVnkVYSD0iybBbPzzgixeHJX8BH8vQHbX1wpkwu2zO409mrEAEu4LnX34
E28J2+2kmGPcgmOZAxzA6oUXkRX5kGOIvzUHjWs+8xMlO/jZD13c/gNoBfEkO1QW
tVfVFMr3zX6gDdlWf5WujJU5bcNk5U7RB8sE9QYoo2cDLmOCb8NyYB5pGJdN7hKm
RK7ZuSgZEjdX49TYbQFreqgHBksxBsQTMsEWXkild8OnNO/4dqjPPVHx5/TPEpo5
VM7LNPJhYif6CS6jP9f5cJm1swcEa+HHu6/3D9m0rltbzw+nqqO6iVdVWE9Gj2fN
/N0LHoCr/WItAzFs9FnIn89sN+3gzDIQCYPWwFeK3E/RUieQzwsRwZCXzf7EqFRh
lb3Va95p0CQa9GkYvykepi86shQyZr8oNEEE0JihPA+WzOvteUDV0hQ+Uv2hm504
McR8+6FgY61l0YBAt0mCtYDf6qnhX/r9Lu06SxMHoC6UJNM05YQdDfBiuL4wj4MP
htLNbxqXI4XAOsODgv7WLZGlezDPL1PkgHhG0Rqw/eiK8eXFCzwrLZgVSR+wGN1k
DsCTp5TSGMQQ09lyAyX5Hkxbrpvd7abu1YFD1GFJvPMte0FMg8rqSbn7pU54NauZ
7pI7Kg9BE6Pc05z4x1jJRVULpPI9hBKXLq2qJCwlkrv1chSrE2gTIqcM7W/9ULkX
i9FaDML+ma7Ulu7328dfo1+o3YSo70g2jG0ZL0WwiX8A7naCz10sEVKrqJyc48fo
uBQTK/yzSVENHpZ/1dS1o2wEm3v0Gr+w6SZJ1cxCjJvnyFXrX4NS7SKY659clVOj
ICEstMYH3aGXa4mwYNYk/4yGpVFXuyQ7VBypTZtR+eDmIYEbu3ADPHC84Yhk/1Sg
/+xVpWyqwGnYYU6qiQ0wlWcm2noHRklqEe8xDACoeB8zfmkORWS/wnoDfQO2zuOf
aQ04zQ2TqpPDl2hwbjUh03Eob0yJdd1C5mOSjUn6Z4STaxQ9ISeGLdjrl6g/l88r
2xO24DTFpmITywIWDqjLMTsI8QMsBdf/rz34H5OqXFL0WZH9jdVAjWtgqVs9BxE9
vE5jNjvKBAM6YpEzxZluWDO2J8DfrYMWj6uXQyrK8VJqtyJ4eZ5c/xWY2Z1jgI3t
17k/OTN08Kbm+r/2jXXt+oPwrvfOldLi0LfF3FUUPMaKerMv/i+BwA21/EZ2k2bm
hE/ldPFc/Nq3wMjB93zvDU7lzYTvyrG37IbZ+/JxIMQAqXxqGD5DtSeA36uUx+T+
tfYmbWQJaW60nphwHmADpz+PhsfA4NX6VrMYO2VucRdXXVXhH4uH9lsv0XMt/5gl
I+x6xhlBiQvPzqo33QN30ZMacOoK+FRBVT9MiOMnKGdn8ihl1VFVJ7HZAwgHXtp2
Cd4G2lvDdRiDE+U862+6xsYNSpX5bk2Vw4KXGHxo2V59q7xFitwP9q+5bN9Fm6N6
y9p9PPNaagjLLC0Ch0C8d1M/P6hZfFgKMIAR/5wr+XQd7pAcSs0wCvyjdejqtls9
CfgpLC/AyUH0U2Z189GYMmS+4ku+vD6MZZXF8T4n9sUdrBrAD5S4QoR1WdakbcLh
K1SyRU+7HWfAzW7ZnSCokdiFor4GHAbUnhXiA1otZOZlL9mmE3zLzUIbgWJdPHGC
ArKJ2sxu/GJzeuKzvl9ucDx0ftWAK8Ma1Py6onkj+NQU1Bw0Y5/JelggTN4xREeD
XGMchJ+v4y8/kyhZ6aA+FAaI8xp5K7MzDWWoPu7qHd9o3mUoVR71TQ/m1m1kc8lS
C3rI2H0jTLITmzyQnwJi3UZip3EI4umXR3jb8ngV4cnU4YkAmxtwM1CE1OmjFWeu
AgmbfSEXnsEMzlRjb3shLyE+dS8rqE7JNOwhtTADo2T63Yj5qiZUURKecUSIQqr/
q5py0ZenRZuY2MNKG4b40kZMbda5gxyPFfHyupM7xMmtvo1teCNmrjXmYGpRt9ap
7GBPmtTlqWOPOVTg7GEpHBnOFwi6QBp7JK1WSewSkTLuZI5w98Ad1gEEsABC4ZF0
TFfJ1Q2/X5JuPkg4Y0iy8UtLjDQz/1IGEmkcisawFADCsch7dPSSh5kdGE2OnIT5
eiXC7D4beumv7QLYP8/09sBe5RwqXcmLrhfHsuzR0QsLG/Ue0JT9fkgx3WGhJUU5
cFE5cT/qBImWTYgO46wCZZLXvxJBDyd249cobkZlBKxmLQpEntkGUP321Pi+Ln++
17fCKdQ9y9AAkAa1C9M+/BTvEljwjWbDz2RqZnboIRSXK5PPXglWg56Y2gV8fzKb
xNnHw9muUHG6PF5RBzBeYpReSE30Ubaz8kZlxPIlsm7dBoG8ZFEq/qczwTs+iW0n
7eWFvtoXBVfzx5d0N3GPbHxb09g4Qstj1Ct3dhyqWJXCBbFwANiVDsTedJdy3hbf
S6jb7DLsEzrOMaJtHDw0Kg4SsL5HJdAvmCmqYR4Y8npxmgqsGA66KDRxmwj1AkhS
7Gk5Q/ha4egwDYKW/6QhiWQ7kp+L5U76GTuTn4VCu1ZRmeMHMuoYyiJ2SjCAqBRm
rqxre4Dcq2GoLWyz4qAr5/V3O5hGl2xhQBEC3WHLhZMWpQM/zuQCAhUksBtGNAqr
B0gEKJiEUlbc+ahJlgPWDJ2Ak4OGiKVGYX+Xvg1STHnXj7jBPMvLfcPTQg+j0f+s
hzu4xYZwg0CIfM6UJNQwcXhegDWUn/5hayaFqOjrRFu6kbcKkW0G3sf746UdryZd
PBdzgsZTfdgKfjBaTb5PK/xG4XAN/mdlYE2tGl/ZNWvJV6N3L8nPHoGTUS/m/8iH
X73+Sn2yt4NLhS/fwhdfJf7O6JJPa18hXEs9lbBdnae012Xbn1LvEgYSjH/NwEAR
A8nZhdce4rdHfmB4aSrQNcUuUYOaiXWLIeHPSUpkyf16laUIQYHR1G2yuxnb/QT7
vah4C3mye+J9RlEF+VBm2bH0TPOpvQrXBtP1ueOcdsJA3YQY+cE9CetHfAhWEv1s
Dmoewm8Fd4wkRbc28uZiLszLPA4ayFjEpRqpDGenBnu4DQ+hni9mpOO/v7zEzd8f
DNyl4svlzvi98HKTCTWxbS12tSZ3EznUQ10CdskndU26aMZx4A8+Q0qVqcFL1XDT
Yhqc/WtyuuRW9rkn2N6h3U11/GxSi8VXU4JJQxzC65pboceUI6wicCp1oiXgI4HE
ncYiA7qkcz2u4sG6qAS1JkbGNiBmcaeqiwjHBZq3AwE9Gn30ZzCZ2wCuue4AdtlT
czh/+YTOOre3AvOQcyK0OTjBwxHTlW5auSQESTnUKg5hhsSAnxxu9Gh0PixqwWm1
LcS++zhdNLIe15D4MEA70bdAhofCl3RAMdAIAsmhUHARHUIu4SKpAxKEQjuztSOv
/Z98i+e7aBijQOv2Qsnok9bcdcG71oomJAFscRRJxfTX+auUpYa6VTrIZ+vtrd4H
TnAK1VesJrcdQP4XsDHflYZU8ti6wudFO4pQivlRQAjywq4i2aGfwyTCSiEeLAC0
+sKi0wvZE2oXLWLRhQsmwFWTZfb5EgyyDeUvqeQsRL6aC61xBwD82Soe33bhOUJj
d4yjwzokW6SQfJDBh/143YYzO0D5w9hejjyx86iHis8ms20mkVT4WHq5oyW8427K
ap+iGzyKGdIvnvIje3CujVRVt2OQOAPbONP1txqLs8eFPKkeSk437aOw+MEv5eXH
VTUBwGybDBj1qLtej2fC7jBXsxEaWqydle/v8myuTm1Z8lQh25GR48S88LjdrHvR
UfRc2ebfkZtm41FQCf6E0rM7wxArhPJ04BmioatC5kuPw2/5W78gVwyIQ+JMbZ1w
STgvNgcAM3bqnECqiUPNBTV0LgYaZXtJU0nrpZ2UwZzDSNmOM3L8H3a+RgqMiV9E
D1rK1SK8EW+ziM0uI5ORzdkmYMTZ7HzsaT93jqEBpFbsmC+F7OAtBH9hhb2w3CBM
3vhfnvjreQ+/rYHwuzv5I8hXRX0dHr08wBN/PLmiO8yuzkWpuYXKktb3RVoK99se
cUsh0t7mFXk4joZtfVrWzM5vTbjV4S/CJsfueb6kVp6FVm3Zx0GrJ0eiTX1Dc8Xe
n6lFN8SVwf7baUTdBR6zmP7cxY7pYrXTl7h7LEOnEktRlh/cwxic/HP3JZvisyPb
igWEJHD00MHZV2MA6+gkiaM92M/RApYZF0XH9e8XP44MwBTZfvlS793OfBZTvBEj
12TC4BDLQuMNJzk6HnxegX5hBTnXguDd4eJ5j7i5wd0MEVnOGGkLQEmsEVLuVCiX
/Joo6//UtZHpZhveSAC4lMiF4uTSS0m1seOHHcT3ZpcXI51t5fyOe60hkPOcVS5t
ipKWi28b+R+4SXb6NgRRTYzChohN0mrUdGEW5EWM14GXAD5daeizABBUILVhEXBl
qT07VLuAdLBJMApppRaYVm8RwWVX+4aR8KbYsx3MH7lL9asrtWJKFxJkmMLp8tqG
0AMEuu4o9uOsHu0TegV9CHrrFzNV5ZfG10bK/8dFtEjJTOKczk0xUQExhEY2U2QQ
kTDwmN26K40ASJSyMjiUes9qagxJDxkW2JE82MQYG5z19ECeWMlUkLcdvtJsP575
MHqXbaMouR6xeiKailrEuNJR+5rYuFhlRP6ZOx4lz0sRTRwGWmpajI/WaiYUoiPv
CJkZt5h8qvmod1ZIwEx3+9Pgn5PS6dqghBltquJxxh5k78dgnZ8HUyT3LMG1Qg4a
fKd15IWE3/et3PYAVl+EQvPjnkH3FzpHydZKQerNu1bSKL33wEfaTu3Npn71pL4T
qGNNZGDScs0a0cEFlh8W6j+b7av5mbHStPjb3Ag3tViqO2Q5qDjvokjK1DrUdbOG
WgPWoP5+m1kQC0YZclp9mrkfpgRLu1CsJbV6ixMbWEdZLUE7X22qtz+1+qO0vQQn
nFqergNmgsMAfyqM94ovgr8mZ/uQVpDOIAvgMHx7pvmGtsXBXz3mkg6NlCSE5qds
OuZ5X4sat/ig6QLg43L2d9TAOvfTt/+dtAXRKAQXzQEjMKAmEyk9YivozjePV6DT
nS8QtJv6X7uvhBCRATD+zOwxXJhRXum5x0YTiNU4LWfn3kQh0ZjFuHHqDO/nEaG3
E0FMPxT57vWipfXVWvkrZ1iZzelX8+O6fgWcuAW3UZFGzSQ77j8bc12JnHsyKWS4
NsVzxDGm0LxqBRgQOPSoE55w7j/1jn1NoamFXOiY/li0V0Usub5uCPRJncpV36h/
LbxJahZDq3pfgPyzrHjOw4tKZ6c4hpCtEzzFzPgEmEYsBykUA9pjIuNUUh6Cg5oS
uvhtxPGLugEg8X3oz0FoMskneYKQ1h+dmGXStquuWoJzKLeb6jq44MC/qkazZdxZ
FArB8tML9Qvhenn9DNJYBA0ITlguAVLyuT56Y5zSuB+GZOXiRZNaeVqdgsHHoUox
8ez6cS6GlsaTl37VwKbBmFd/JINl1L/APHyvJdClpZtF5vJ//AxxtwuycGQVtuvf
9uU/TXBOw+86zLQjMvkAaOUyUZ0vtCJeAKqbHyLA/N+UY3RIkEWKN4n/vffjETD/
msRPbkG05K9+n2Z5pxBXu6VfmYLeqCj1wWwIUukfedOri1x5/ruMcYa4cPo5KfUo
6b3JXjmhoOBJBrj2Pnf9FKZLlxdI996cmn6Zt093JhT9jhWO3xJ5ZGzYQdQJw3ld
2lD1U4q/kgAGTV/mQrSR6AKJF+GjTei7pE+IEXUUp2KgZnRqpAzF2mswfczmC60y
2cmrWddafLOdN1LLmCQf7tHoJbgOPhSrdOOIAzW7J/JEZbEEZsgIyfFRk6eMHHO0
+3ADax2iZQq/OKPwy2GdOeDKxfuss6SfOaI26wdpf0EpltkQSu0Q8HjLxORL96Pi
/A/PP/V0M1sA5Tv/dAZkk3WWyOBDwgKAS2f4H83wYjs+vDzzAHQN3Jp/nSQYU7LW
nToBSO6IS5IftWBihwOqkXi7Zk7zXLkwvA/rAEfWWGoZBO3sslRnFlK3JN5uHQ9C
q806Z9aWiTDGotrfrXrrOiFfYx9/rzSvOsFA7gPOsc8/mtLUDJTufwnXse72W/sx
hEBa/0ggBYaxAkdE3dXXPCZ5esadc+j4q91oiJpZAAr7ZKDUx1u6E+uGOuhXFiXn
HAEekikcZfXN0FWPQstw8PAlYyqsmp1ZLOslZVPlUg53eVmvrv/Dr1BwcDAOPiIY
htAKW1BKgYhLPgsg6gQOIKXx9rxRrreKBsiIuGRebIaFUAwUfTPpQ9QZTlq5FLTp
liCyRMdBXXHbBnCzIOBii1FSpCROhe03KevEM7/I6z94CUaOtI+3M9Gwbh2vguhk
kK2Ngh0DmmqLVkbqJSegNglt/pH5Yi+Q5vgd+5pHcRo09pLiRJFa+GWUWRViP2xR
TMj1qMd31ex/9gdqW4I9xDnthZbzjItA5c+p4n6Ns6CPa6QqloZXCxGjyN0vuqoH
SDk/sXR0RwVvHGhl+9vrHahXYOnYnrrimEH3KDyDj8DKve4IqBdYlyODFh2wBcmC
wYgdzT8rYqDt3MFpBhTQifN87hm4B6gwsI5XU5HRlzS139xjL0JFYwj9MmXX8uxh
Lsk+2aQGkSTYGH4pgnWfV/el1YgKNpAVtoJLmkY56lIWRjaFdsc1FlI36lwg/OIe
64nVdzY75bdAuVrmnwrYOWTpoCpEzUusO2ay1f1tA3/uUtwJYEpR3SV26eiwy27y
mQv24J8mvHjCnS3NJt2jfgb9SZ4xPcBV+5/NzRjJIK5wYJ2t8usqxNHSjssEmbOK
fkk8SBK294BBpVhh4hExbbDLWv8FSDeqkM/ZdU7mn/lS21V0CenwHcK7Tb+IUjMH
DhyfSgOKIgShRlMpExqVzKi713rY5C4D0zGeJjOC+P4LosGzZ68z0yUBF34S3bSu
Y8DXnb9i+OnRyQSjaXTF0dEDE3D8RE3fIONTGPefFroj6Lyp5uHOeJgvbu5LuAP4
/yJZInvjlS95yfadPhBGnRqdi8dcZoa/We7+6pYRcNsI8BCeEi5ZbO7VJeOwJVtm
xN1nE4pfATyxfD7TcNE5kY/qqo5BniKz/QpOQRdQpDwQl6W21GsgOIebLAEju181
i/N5m1ah8UG5WDswXBSItctL5LAtxBHruqBUL3NwTgRPpeVMsBV7KDiYN5ghFiKx
MGVbJawB5qyKVnG8pKJiNhF01WBiGlqyb/cRnuPzfZE/UzoRJYUVQ8HL+JX5t4Y5
ddNJn2KVdYvYXwvkPRHS7VQIf8KdTH0flgvS4hIHBlplpg6qPanKy+cXwn7JMmSI
O3gLr6YRUjRm37rLyUMvS/LPctqqgTjxNlHpPpDp6z2CSo74n5pfZuTF96P/WMfP
ovYlukFYmV/RY7iUr1WzVPZrl7nTwa5IFDcBIsllhundBoUCWvycXYwP6J56TncT
mwZB/5awObELLGDGG5/r2JHcdZKcTSh0cT0yLYKQEcuMbWuBXrzLOZ9NkQPmGWHP
LJ+HI1q390oJyVKb0FHpRLcS6+K7nn5nIIAxY2L2rryvMkcrnEdUCfsTzi5tLUe9
/XVawRgfUjjr5PkSToyk7V8eVWjBK1dp1kiRXzCx/UVzZod/igh/AXNMU8ehl2Hp
tUZWXBB7T7WDHsJTmyud2XZYvkm/b7peRM5hmXq04Qe+KeEMnPOLM3pCrxaHv9Nh
kg81Xe/dDTeNK4hSnrcS+mf2oujQG0Ni7MiKycOr/kiu4G0Kx42A9pDJbVjYT10f
IBmp/aYAf3Lw2MnrfLLXGt74hZQXvKFn3OqGl2Z6SIL+K7Qa3k12hTUAkcbtSeqw
TNPD5w/ReOnX+EvarZKeFhw5ciNlTRGgyyNUKPi8LvzlBQ1biAWoSD1+RT4MMd4I
fbQbWFH93S5IuosVpFM3NoUvKCZdfKc/GSc+/0h6mzTbQTDXKKFKQLU5Rz6IZB9U
gGjIJnzkPxe870inv1qdsLTy/5OlvZ5qvjNAobKwfj3PLlPC8WJ/Vfn3PD74hmyv
7j0pTCxmF5yzZ/D3bEZhFQGnUrd5eNFIPfCrZ2S1djvy6IBbHRZcoFWmTRVM65Zf
62p5MYF9AlcDGFBrJvP1bneJ97+h+cSvLei1hwECIy6yBJYNG15akmTh6E6Ba778
+vFtF2/9Wni524MGbnBVpisvBGlda8EkaJDAXITbSR9i3qzg0RR/ROMGlegJfrOt
scYUONodWJZPwOXiFmBpFXklXooSnxe4y8DAXO7Q5lRTOZoLNLhJqaSKX68H64NW
TDYbNGO3BE3r54SzF2sZ7G8BzF2L8+fBENjQE/sQmDsYsvx4bDtKDq7BMLX+Pue5
h4trag76Dml7k//staXklp3bSmPLHmXqf7UAV1UVjq0GT2zpuWuEN9EzdkfhKp4R
yF9NjqPyPi27j1gwNcf1igq/d0TX04wk5Dpl4PeGAKWZaTv8HSmbTbbat+7BSClp
dQj2GanhxDjJFtUU3/OKgDws0nqJCCLFkpYQk4s7ZZP4Y58QO3WHdGzsRr06R0tX
yXBDSVFO9Ez3MDD/rKsj/0Z5RDSUWhPVNSVCzaQo44+0RkpDjpoBXEU66LW/hoP/
Fg/TcSdKHY4OY5bYC51/9oD3zPGc7DF+zTzYMHcsLacZISY7XMowoSCbFVocq2XY
AS6ottw1iSFvVFQVprBp2y4Gzh95+m0SA1grKjqTHAFWG9VuV+TR0+qihMOFVLJy
GjSJhu1eLhZV3aHRO3Gdv1zcfsukbEoERcEyfNgyWgA5VFZpAc2UdaQR44K4Arlj
+bMF5wPEaLPK3npKdJZOUek+T08ekn3WaLgYx5A+ghwjns4DefXBXKA6nHqHMOJk
/uXtHbvsJYHYMtyz2eeT3fyUFic1pVFSC0Ol5YhEDMTkLnmTgUNYo6r2/iUAXqKE
k2AG/ZP+uWmeOBB9Z7Xa+9GwGEbpidiCsy5+E+jkUkIOeWicXQvoCPsC5Wbshz30
swhVpOcw49oFDFVlFnyo5ENBKXD6Dvt/EG5Lzsyy+ltALHh28UwGERb4dff/PDxL
iuhbEMxPDyBmGbaJROeUguzTimrM+UvwfdS42+O+p1CBLqxdJjQbNFXPYAQeCLIM
K85+jXbbCOClk8SVgbzu940mOCq9tmP6P2WvAM2G3wgbTcdnP9xw2B5PLJcjqRad
uKPYQLK5hEoTOlotIKWS2GC7Lkdtza5Rd3mclUZ7m0RxIAQ8h23oC/9/NeyOaBSA
Ed6CPsMuCFx2V9OD/flNkgnzosZXim5Ii2O45cFJDPkcAn+Lao8LXJBQ7+h8wrRK
PI5Wgf1ICG4IvNsCvHKgUFwBEAGvOsjzWaQFn/g5yU+JGMdRVptc1qrFa3+0clv1
P2bs5NLvmGZGNymUG4kQCbKb2iNwN8Z0hyyV0gk/rqTERELV9/Rx0LnWKMNKzHlY
0CKVrzDlp64bVPUhx9hq5hMZx8JY6RcRmpjTgf6c7yDySrEvTDuqE69K5qqDsP1C
rInHsviWdImHZAlyLWHx4vhQh23sTmGdqInt6Cno9b2055PeapllrUYp8KL7lK/n
SBOp2wywtX/Ke+q9XfP1lUXrfiTfMxBJsPj9v4YOekbGvRHAR9Q39hrhpZ6NadI9
FqUSE9tJ8kDG6hb8/mAr+s/TtxftApMSYVkruc+PQE/K74KpYn3uonpuf2LGFtoK
j0WYvN8jswg3QZNKpTG0vN8GtDCI4vZ9zem7UrkkNfblFGQv4b7+f06yZFPQOty/
CxJrtAffsgs0kpNSyGCp5MHXJIKCiU4SsiiVqZguBHnU/LBQEzukAKo0GIRXoBsa
+13R3NCI+/31v2DXquL88GF5NMz6dDFVUpxK4yuyREqzYVPiqsuBBVughQ7NjGB3
usAX8sVfUyt++o1a+v8BmEfPgBQGlK+NrEgmU83fXEskRehb2EwHSSJBBT6WqdYy
QMUMHsubV5CJKzt4vid5JZj76LAAAPeQEZZ/KqpLRW9lXlULu03VvmxPRJDJwdjJ
AP/8GoKTUiYnEPvRSrMHJguyL1S+w8VAc4OirdXIxtE50d+8hiY8gn0tlbwoQvyt
BpFHwHWIEkQSRyAUPNLoFz4ha//eyw7x6X9H40tgjvyd/7vzqrpMXFGYTXDuZmnX
JWQCX0njKY5uWHHC3JVNoHvuJHpP86ISPuYA69zNcbWYt+ChiOwiNaHtMC6PSZum
/i1q5sM8OZTj8fYAkZuTKOgZRopN/mZuzulpW0S8X+4FkYTMBLEBQdEFBTXBRmD7
ZLSAIaynFHZ/J8gh6hsFTY6+OqvnVhehRZq7r3AMHTj32GUMkd4+UzBUb322R6ZG
EKpS0vbdUdbMfoTt5HwTrDNg9mtGAnbdtb5s/DAErB/QuWYJDLSvW6eOvXIAVQlU
Zt6w3j+Zkp6yv0fqo/KAqscUyE4uNTkdepDWbItobe9ncuVo4KTODfdCqnZODZ+s
7+rqLaKEU8rq3PpMEdbvBr8vuhMt1NJ11hFDKukbeZo07QR88/TV4dcRwxyXH0qV
cZhMHQN6RmygKsrmIoMz2Uz5GIGLj6QokLW80RWYFixxNy9Ik5YWi4qfdn5WmPSv
Qxsq0lS+eMeRG6Kp1+NiwS3XX2U3lAWfSlNXxyF7RjJWSqvc6qHHuXieiudVB7HJ
OaeqFCwkB/rLQW3Ey0xGy+j+FCJ9hub5YaeS2fAWfnoH5tZYZhRnzi/i3T9JMjje
94jQebzcZ2YQZ2IIdXccMeTxDNA1aj4eu/CUdyS8Ak9LIReeadHChVzLdJRTDDuq
oHRtylxu+IwADzJ/aJBfVgzvoUMejvzil82fPIGvXyTzs11urDPZjT5NSm6YWbtN
bzEeRwq4UXUbk305LCgvSR+3+1tjU2fHEsJ4i07Gvj6taTaeH8fYCGYW4kErTCgx
qH043vFF+LCueC5muNe0UxGDxLVptP6SJE/KU+gRm9HsG3RKEfzhd1naFzK3Bt2y
FbXymRQaK2Tb9/nve0SfR/0FRDegyPmEcgcr11HucBk85FBncZzEEGCGMfvPM4bR
nVQNBDdPaO0EhrZ7EvZqXJG7pzCV9RhcZWp5afZa202wjLgUPSjf12ZD+5VqPafN
Mt2WyC5m6jAR1hCjt0VsgMWa1h5msyAdcTw9OvcKGPKJFiyQUdjrBMYfqGsiXE6O
z7wrfl5AKt32D6d7nwyhxT6UAcWbFbzyOOlwBsOP9zyNy42Ezd5meJzDz6Bwmvu/
n/TwEsOz+44wpXIrK+fquN53GOJaVacc/dd9CbfRKTACW7yrrYcdXUIOXXqIVmIG
gpRRQ8OgvTypNSOiv9aoX43SCwwdlKpVKfMELSnf9HNY4A5hcvo/HAlFHZoLX49q
o4LE+KBOlpCIJuY/UZLyhII4dNcGspOl1f+WkpT9FuieSw9uP0oMMkymNgIGY4fw
FvVmJTyJAVWrh7NlQo6XSsPc9sVN/geCNo/ViFKZo29qgNA7mnMaBqafOkvYWulD
5DE7fp71yyTgFo17NvYNFNPvz7QxcBfU4SaFId1PbsVyDcvbql9LBa2oh8jm9EG1
+ijpv0g0BbWWppzkZivXB79nz1aIsR0ZA+B3kxD6wxgnxUsEvi4fVW4oyIiGSgCk
nYNKVCCpGT4N6atTwr/wtnf0eYXUiNvTt9NzGRjOfu9DOVAFwjxrc6SZ6g/MTh+3
BXEXHD2W25Pz1TeoEteggawlUNz5yZtY5w4Wk40Tiklgfr9dcWNHx9V/2UZVVnGX
5eiIxDtmBt3zKp948LqTTpBUe29rZdkfSTWh/1/k5lShoq+IViZgGKof7z+xA+Pi
78tNsTRkBVZ8z5e8aZgFnE86ETGQ1cn+xoeE6WiH6CDKlM62H+3dqiSds91Boqh/
oUeZGtdBh+mF7uF0HzMhwb7iulprCCB++DEcFuG5ermwplSh4ZEA4STuuH7J7XhY
e4jo3Wr6TIlHzGAbV8v88actf49Ov5OusYwQo0neI8S1AXiOYF4BZl87q2nIhJlU
J1gtrqCEBw2gs5/fst14jAjlmkTsojVqhth1SKFEL/EJoqNRaOxvVgYswfAXyiUX
xChyHqNa90PPazV3+USBMqvw79LEUNcj8q7jvK8BVTk7mpN7RmMGXodjg7who6cr
MRSLj3LGwkn7VxmwbOlcs3AbnAtCkg/lEOLlVnqgKh7J9aTThEw4HUeV+lZZCda1
TWW1SuWd+i6P2n4DyM4q1EchxwjfMXLQUuHO1ARACk7I1W7r+Ny1BHnnT1LUmLU7
Untn9SNcet6a4Mf9xq7aKntb6hIjYaeCoXP+NNx2W2TojvqBqwkp45MAGIn8GFiK
7JcFnQZRNLWsPv+VuiXYdVtDfKgBidforW+v7aiZf6WuEVBPiHNtNMfHsznlOYoT
P1lxVR/3ViKcMV4lzD0nMQO3AyH37VbgUq69h0i1IoSo0jqONYlcknejU9sqxUau
+iP08NM/LxOhlZFfPknxCFOCR4ocy8JIfUW/zMk0djGp1HoJaQOJpSlrtpHbwp5/
kooMETtnVJtqLa25/hJ3lEGDkFmTBjEmOpyv0S+CllfB9gf9+eRoRuX6LkmjgxK7
9PIZ8a8WClGN2nWbKSCA/v53oIhLfj/IP82BOQE6gmTpjXz0p8c0PUNGZkyZ44Gn
fSoaxFmLDDrI1QueZ+mtaHReXQj27U8mTronAqqWqAGieUYHYoJa3ujPGpSJuhQJ
xY/AvAm01hv81GRUJTwG4KIhnXcQNhhN+evX1Qj3nsqhOpdpEDOR94qDb1eg3Zne
ZBTRMmCV0vSjXRijYgR1WgdWiRhruyWM7QEMumktFpsuf9LnCNyfVY1yOsyfF+np
8nDSJB+Y3UUdeDXL5TQ56JfBkMD+NaMaS/Ih1w8Ry8ZlpDRmKRjK5+aWuAkoJnLJ
cvLrvVgknWu/oIj2YgT9uDcDUws/jF30NgYoMpu4/7Ag5TBZzRG0VjYmTmacxWl3
AavjymxS2YqFlZ7euyR6JtC72w7E0UFsQDSVxKy4OsF5sEFS3lCyL4LtYjw7Ac5a
u7STIKiUxcn09a4oRv5flmnOukfbNKGsDG5wioznmRkrdrzOgR7790RbJ605Q850
ckyviiVlfqG6Pho/8gami4eOy6Wtnla6WN259OFPg0piXWNyUs3BObPG/x3HQ3Tg
ZU/6zJqJZD80iwh5IJLqQN8hTigDlhQ5SvNx6O/EfbbR4Wj9is6pem8VqM3SHc9C
8/InYLNqPViXosJsEdYSKnnszUbTi/aLxX8CChI1Eef49JYNiAOqtFSozj3ehu0i
0DUy3SMYwrDVAU5CJcc8rgDNf5jsToi1uBPurbJfmLky4Wf6p5ZOxyzZkNEpBzGW
HRLxKuOQYYj/B8JQ/+NRfRZpH98dTWSZr3RhbXbbnxix7ZMxpMDCwlSTcXq6kiF6
3+mz59q34m5UbQsfgwlmrN9vmbRG2O2w5XOseWS/6fAbBW3Zl2uyzN4lG4Z/1hgJ
5UDl50ZL7JfElUGXpAsQwYBejSc0HpH7Klc28izM3Ubh0VJuBLuGTir4xk40g7P8
9wktYCMytqWZucSzfDd8Uvm8i4Q98HI1pP7ppQVZb4bXvGyLciXpUy8q70M/MGk0
LCL+4wGAgpUX3oz5Go9PpaOlMtTNYXwB0Gdzn5nC8hFG9IlE5jeLYQDoVyCT+nwF
jGF2GOXw86EEGF4lkf0QZDqvk+EROuDRxFgUKGO6N7YtJT3dgYPtBxsTup+ua60m
c+CrrEbmaAHV0D27pyTKx5gmx44l1b7bYHrG2pSSIsD5z23jKL7+AS3py97M+cHm
ogTWEb+tACwd9ayeWsKovA7xR7g/nTTUNd7fAaHd9hssvk9SsUPSYjH+CLkOePwB
jq7mLuuPw1S5V18SxDPje6BkeDw8ARHCeRwcSz/vPedeeOrr/2IAQJJd90DYXWXN
s7aqMQp5oaA31RLcG9Ysilns/7D0Gd/Qe3OqXwm7k0vvsac/1iKN0ddZQDFr3KNn
/bxi3NdrWwrP3S9hR4EZeLl+WSPcGcPpepGAUN2ECKf68bVVzPWgOStk08pXKXCC
cnVRM/5g3b0n2NF7oTpd49JMpeJ4WEgvwsLEk4G8x6VfVja1mADcMkFe9O7N9A08
1RSn2ZodLD6IXsL2lD8rT0S0JlJskdSlxEGz42s818/9wfpN2n5qYzJ7258C2zRI
WIgt6Ol/6r5dpqFGrqq5k3olZr1MbL1kSsaIjy+UPMmmXV8pGF2+pdW8nT+5HIPm
ULvmWih+y0o100pEuof6u/BaZw1Nb7rqTbIsJfojE9gff+urukuy6VnJngc46IHr
lUQGtuFkdrXBh6MXBUK7EdU7ZQJDy2XtN1QZyqGcOEA0AjRU/jYuuiPLzcScpbtG
YweQKsvOKAP9UKXaoKymU7GJzRJzJEV7E3tvUbuE7Rl+gUubKbkwlSzN2YSpWL62
a+QN8BuZe138ZMKTq3z/70GDtd6tq0SQEgC4Q/e0FqWUmG5FZ9SYbQiTKtxmI3SP
C2/V/xenD9ED2kgqaujrho8ffTeRrRxlj4oSsqkBsARmAz+trMj2IrOq8Y24Rjtm
jz0BLrB4GJZXG+yHUFxLZd0DqT8urBLq0NqP8nCmMKjcHL1w+cu1BOVIr3+3+wgr
2vWcw38J0diJBpesxork+K9pWCEtrdB6nWjArl1R6eISSL7BckyH5jOx0mCf7uKr
SDxixAviAMvoM7a1fnxPSpLCUh4oI1Lh1gLBO5/liP2wC1XLgvNCkKXePrAYFKdI
meAHJcLgHgf6fsawed6RIAzQQ2JrjRLJke9aCAtFD6+tcKiuCx4U00BZsFFiCw0L
4KffdFSrNHfMuzoXQl7d3nFqeco43B1CejeF5VW2MwuGpipRoqOnHz/PCGzF4kGP
UQLPlVQnvcAboVVuX8nMFDbpVi4ULLCm7nSohCh+kB1S/kDN2S1jj98ZgsonW3rk
k9Yn/JAG9VsEDDi4TcbXf+w4sPFRgUXs2w/cuLGrcnQrMd/OpYtZJQ82o7vqFDz4
VvkU9KiIOObvnR0L0GeVfqwmUbEtDT8iGmfGMOShoK5V8cS2Gz8ocHbNPEAeoNnm
vQXJoO4quom+Lg+MpxqzyNy0S4/0GhXGhDW68L0UYosMdyTwEnmb36QymgLOBqYq
A/cxDbazE5yelMFFyhGTYkk2W4BnNlQ7LuHvdCbGiwr80SXmG7t35cpBecT+JIjQ
fVP6okBG0H9gRHFQOLNInGXsRpXYbiEh0xDgKH1WdvWVYhyaq/B9BLzEjfYIUfDA
rxMhlxKBmS5dT3nZvto7oOOZGcyhXtdE4wsFaxyXHRnYUZ2vV+lEJzcVWDX6qTwx
M4ZG5bTEJDIZ7K/H/LDpjzWhgSTA8K4mftOsfpfLjbcc7dFTJviFQSY1bnaq9wai
ctYaZVYM1yN/WSRr2/OgnSzJaU0yKbm6igkztOplsZYTXsJSMcB8Upk0moKCxFQL
9rsJCZgGVMNcbrJ9x4sqChEmag/3kj/mflgELIPixyiHsM+SRaSwqU1ReSaJTzfp
7JSYa6ipJwXiPMFoUhPU15t27ARGoPVI0QRNNTpqvHhug+iGmQXLSfUNmsDtxu0v
TkfM9xqUCGcNoZKv4WjAugZtjwI5W46poBGKR0uvLfk4OxhVqpV+mG4fgQNfEd0Z
YHUDvNX1goRf3qklCyISHkveOCVx0c1A/lfGo05HBaK3BLEs6nL6NrCJfYCrCpHl
xTsF7XhIKP7Q0Rk14HzbZpW6khPI93VVDC1nENKkghcIJSkLIV2aBDXPPu4/In5c
y9O0mFc8qRtkrY6HLyDRovsVrPoLiQzAvhx6nh2/LkvkBNCilsgR4/VPEFj2+cp9
GvrLsCzKEUsf+Uk4fUV2P4F8b4/ASdh3X9i93wq4cJ/dMUFKNI0/xd9b3j5MfmSY
hmA6gSt3ykzG1titQD/zfUxzHzkRId48FRWtDMzOQ3v7Ed7Pt92ONZvG+jCZFyxd
nPtaKefDD7rct9ZhzcX8Yqe/Jb9DqYzRqvNTu0grdka5B+rR7s6fIXFREcCyWFYC
JED1f4u4lJhIwJJeTOyysgrMi5StlcHNxVxZWUc+IrCZnnINQR8UBHMxvR8P2vx6
ETy+4WeCcBl0tQ9LLL7XBbXCLn2lIgIQXaZFWUk0NFWwQ6HuvVdOZBtJ8plz/59p
850onV71yBtYmQ2pmRK5DZU9PGO8jaZlwtjVq7e0o1qmW8vFsuAMXjiemYdFaJbs
fbvJ2YYiEXDfX0S5RKuCa5ri8NhCg23qziidizajWhoLUcuFG3iiGbqJUlwuM8vG
SC4PwmX/XKfd1BDzexhnRT5r6AHvvY9RnUADeSUikk39gpHL8XSPkuDuMtybazlT
nDKc/J5IBTdqMiXhU5Zjafh3q200oR96vdbriDpntYwc0yW01MDuIQTUUjT0rKfx
Wx6xnBUwoxZTeeq8B1VvIV9xOvnn7unti6r+yWMaNCEClCyD7quBkFwUMr/aG1Z4
LtqIEBMV64+zXCXmIXJtt/kiqJBO0xKYU++MjFbhs5V9d4T9YsIQaVPh+6eERMwO
zqXyWXvVb3d7jVGda7ANF0xKo3QaCLRU5rBl7hByip074W2IDGdoLhbnBPq7mMnt
ikYIRXdkSMq1JJJetmerA/z4S1O7CdC7H3J+ryDqh8mN06bmpgC9fxyB3CzawIPs
bzsDWOQyZhlDhDCT49U9vhWydPHdmDOYPu1FdLQFC8p7fG3W1uTcm9NnRo4ItaDG
Z1aXt0aaJt7DmPqB/juQqAtMe9/JRRHIzbFYKq1CL1QdXbPuSiid5wbwnBJ84kOZ
cilzEIqPU/cArfgQN4PZT87u4wZ1abmzHEdJH8yr3qwNTshO+Q19avKybS6M9eDG
yN62bmBTL+XejHLSrIENvmM3oRsMwwaAcWsxBVn/ORS9oQVeuj5yKnXuzvUTxlRn
5bcY44emAvdYO5hesmkbXei7kf7lqNms2IesN4dqi8azjCfzFqrQFEY16OGhssIG
d1lir8r3GI9ntoeqkMWDugs4xZRqSaYNaMvJ6ht7dH0zZDMUJKICiVoTlxlpqQli
cBN22gpXEUA+vrSILVVmH+G9qTlKKVFQni0b8FxmB4lO2sJTuotmKD5QAiIGX2UU
bI39xxGlgTvfGHi6i2MqXSNYSdXYT1k1duU6Ubn859mn+nwDXFifiQSRP8a0jOaq
4mLMHO8DdPXTXTFNvlqzmkUHbiI6h6TlTdjDrfVAXQv1s4ZtOSAO9csGkbdGp0qh
u6LL0CLboyzhQ1fnW1CMXk3WygtfWruPOk+OCD45Xx0XDAXLZ+Js7wbFqVfQkiU5
M52VYtra/m3J4Llyogw2igNDB42gn4sv50egSLgMwuHO+9xT3eDIwQQJBm2WrjaB
gCZYGcnok+HZqvGw4l6519LHrHIqfJOTHzdVUGQNMJKyl8LhEaQvXb9LT9nRcgbn
Lc/pHl67zOATz/ogo5Z6q+6UsOSEYnlmfJgMrjYQYxdT45aYSFS9jb5HtepiOCZq
xxxupffDCOpyvMEAhea7dBmfNWG6syydYDtBIYbAB6lSqbtkk/spNs/H34mXljZ+
DGhFztxz+vObvr6/9ZQyLkAcXxFM0CYPFHPqjAK6cvO/ZwdTfbH2bt2ejAw8s5Bo
Oy7dKL3lk5wO8Jzrthw9CBSnBju2FMb8UfRev+2O2nIqAQDyiOaCn0R05BxOxq+R
OhJwQIeyh3ZPDtoZ+WR9uY7hqR4JUi5Z4dHApa4JWwSqevcfCBToqVYYxqPprspb
2tqtUyd3pqVaJPqEjA+1NxEbfCHz5VbWRgC0ONFMVr9mskdYdq83LkvGCcrbI/PK
Bxo166vStQHAjtajheOHToVJWj7hMs3GSIr5T3I3++wwZ5YPtkO04Y1U4RQqRDhu
N+BrugoGIchteUxYIvLmCNhFL1nBjEwKV7VzM+963uIsnOPg5poJDq0oyZgxoml7
rrTnHDRfg9OmAm31UQRBQ2HREWup+AZuGUXJ5zh7hr9kvjs8cpbDOWZp93VgZVz1
qUZISlxywT59TXMWkTzqWWG03QggiD8MJhjX2ziK4ZByAbVzZIgbijgccd1kwy7R
99qEQPy1aH40f+6+pyz3SQn93xUxzSp+xS+7vYHMp63IdRnVGISkWmLw8Yyzfqgy
oqAV7zdFbzZ2Ff6yfaWFLi6+uSE141ETcCGeu5QfKMq3cWVJ42ik0aAehm7Qgm+1
331F753eVJKHTDuUvYS2Vd6+ZOxIRLxepdHEftyMyiAhWfPjui9wgb3S5gqOt/BW
12k+nklV2WemUiAU5Owg5TcbAS82Q/EtKfAuXwv3xmaogv6rE5G4AmnEtYvfGq43
5l1Z7qliGaLD5/Nn8A8ckV/9pgy53LUl9Cmn+v0FegVRqX5BtQwMhASN52D22YIG
+6NDAe2TFQ1znf/2EjqNqnxJ62d5nHvGNXS1foToK7lzRMKcEPXijPu1QtGHQGoG
jcb5JRChz5cnSlLkTvrqd7ffZjzdokRo0WT8/Z6Zv96EXeC9gsdxFX2JDuQyTsDs
b8sz4gQXjOZPDmsvfBxIzE66ccFCHfVo4RzoD8yzBX8BooEPw0fEKHsndNX8gP9A
/iihdQWlYzaM3Nhr07RfrXZhxs/reia7BXMEzqZuZLH1zPW7fL3d9CuqASMYQWX8
O5kZmog5RBmS7VwJ1WCJhhiKWw1NsTu6WRDJYDbYvxNROJCjJ4x3B6qpN6XmW/ep
QnhGWvKamFaDRrmuvc+A+AIxyZ1cDdWQTC4twqoG42JUW39Uf/hFp2kSHiTYtZOc
cCUd+/5S8FJ1vxzk+uVJygzPOklRKSbqzB0emGP5B2/RhFrTUrgg/T21Yv64ff1I
O7sqyCK3JfYU2LXp8GHKStoANZyc73cQYC/r8IoCRkGMTcbz7/gY3zmTX9U06hRU
u27H4BGfFFqu03QAOlxgV8F5zRhZgCYeRA6mkXvhjQFkQ81Q9oLvsD1Zw6a/aAPc
YnltmFJadOeAwQgFJFoDXmelLpxf8STdArtPCRnwaOFU6Rdq+uV46D6RfBUpbcDu
YtXYGpF95D/hqSTHqdCaEQ90uSMaaFwACFuiyg+qzzfmSZrqGXU2zHRbvWE/4hsG
dEjiHTP++q5LzipHYodrOkw/ohJ7Awwl9Op4NHpghwFsmotidFoJICBmSUXeniR4
pBl76+YJBT8JJbIq9aQi0d/bP04jtJA8vHhJ4Kf70VcAhk2h0JPr4nfdNvv5Uh7P
m98S324xeQgfARfsCPYP2laG3U5yHEW45/Pax3SCVBiHbETSFpuSUCIri43hcCW+
ZQioaAd0qKsCq7Tz6kzupoPL38MJu0JSvECSLiOFUsMYkmylx5A14p87cJsMNZ0N
lqu6vsREzjM0KA051OHA6kQM6Z8mOMTHJWihhMREL1cTXXLwxnVG71pPaqwQdtVX
2Hyi7XpYSkHWK7cT+ur/aofzZIY2bkxDnEdShIDuSrrgakR2wET/HNVsKomID2T8
JhkpEQekLBhyMXXsIGrLIUtk57FHQ7i+IfStp0KCnC0QSdq7tyJ6SMtX29zpYIzD
SmF6eiQX6TBVL/DOOB/Z1+bJa7T4HSVbbANd7jI51ZKBkHBhLuXpn413k2rJECoH
BrY55VbsI6H7wpRz1KIJbpyUB0Mt4yVEAHAA2j5dQqkxEIfAR+aVVm1SeBOMgXOw
dBvggGhyHwdTw61vJR+DizgkzAbeCx4s22r42KIkwCPGfMsiwZ6pkvYvRKNvPZif
N1BNU+cwe3KxhlyL650yHsX1j/m/4HrqWGAXWdF1vNunhpseXyYdV/0/yX6WpAVo
zRUJNWmOSAmz86wPykzjW1BHet59CQ+ZaY63QctcLvJpfrVqrlWfeIjEke7d0h9X
418rALzD2T4/tLkyJbi4UkrWa/dFeeqputMaerT/j6+tAP/C2UlyQCMIVImDyQii
I5/0vCRkqq874rBWtSMHMumD/USRyTczpB1QmzCOmrpUA361rQDe9w1N4VIo8uXq
r6kPIwxvx1OZzlvd8X9cnS2/1KBfzph8Fnq1gnbNKwfIB+tLcOyr5HwVlZRQY9si
Em2Bb75xANpwLnvlgU+qZz+yThA5Fp27moa8R6eF6aYTk6cdH1jhPBMYNyZuE8m1
zFUWbsY+/tsfx7dnTzvYaQCeeYPb6eymvTuJPXaqjHAnofi15YFlCjJ8U6QxxL56
x+/D/PZGv/staCqRZRtHgS++A2yg4AFKW6IfRYjJGuh9Euf3FxGyVdVEivp1EDwB
osF+I+KZEugnqyWYrILKG76ZeKw/xiJYoGutMVYTGoWuCyNiBgA1bF9mQplrBzLW
0W2he/6HUHNi8bSzAEuxl3itmpcXI5JnCWGYVE/4rLZj5zcIoazFz38yK1LiFzVk
mJ3ToZj3P6D3MZIWLFWq5HgjgmjvUdiiBPK2iLv2S5CQYECynCpg35gyN9nmV4Ml
VBYB4PBAgC28nwUSCvhkHJ+Glrl8UauozUMBpx1QP+OlEWyO03eet1Bf3w/R07Qf
DaWrTzM5AVSGApE6F9dISO7L2SCRM2wjoQCOVKpsKdgPAMeY8zvhBSnL0hFF8bHs
s52YLx35FeUv1ewz4xIQKa3guDJsMl+FiszmvY8BbEN7Bq4mFCWpaCAt247A4wvL
1g5/CvfWgyi9L6/12fnxVt3K2lKMBSvbuN0WFxDvSrz0HCak0q1OFZoBG8J9vcmL
iuDNtedW6rbcaorqhNXOT5AIG/4VhwKV/bjodKhaxMETo11qhmagn0iRjsii/PMN
DNJtD4S7MO/24et7qhNwKMsZj9L1hsr5L8aj+3cM8TLqbyyuepejNsk76OJy/We/
08e1+lEpSscGu5eApW0zeCNf+tXHRfrasfgdnYhqRdLHNQBjD6NRSN4n22WqpchY
RQdnmLmbTy0foLZ0rCrrqqVkvQEHA1sdYMfL4QIngtGHX/3vJnV8MXJ3XVJjkaai
2Ul+X0WaLzn1jJ7iyMYZEO2aQSIyAVsoCpMCFUXj1ouHVp9RD5cHo3Jhs09jwQiO
OACw2p0WsfjEVaQ4FN2FPDnJi+Aexynx7lqKAmquoE+elMzXjUfRiI7ju/Cygj03
XTEtsZhgSj/OjPhVyFoE/bq5SqNCn8qjNQWav7Vj68X7D0MiJeQzSavMpKYXkdps
345ok6mYf5YB3Knw/xbWhnjCq+Tqiibia4FIGu9mc7zQFpinkOAfkCAuvOxPXNsb
w7IloDhSWdOErf7B/mcMumyWd6NaRt7nFdHV82DZ+Jr0SRFj6fWBrGs5gm3IC6Zo
Fb/5uzgHFrRWe6VFP4LDIbfTav/g0aaOGzf0iKD6oxLr4BuGSrJvusga6gKBIs2t
Ky65eeFg9Q/lMJtMeg9gQa4p/9MjXr/FS44mmIhw/GppuxOU1XfFeI3znwq0yCRC
bZJkQOwcs3qtJTlAosrGz8f5fEoavtq2kmJ17fSXunkDEz/l9xNn8hDjvGFByx+v
cG/B2jSkuPmR75rO/MiS5dW8chMGMBDNqxBIotQ1sS7lzkxPvhg5O+wSGeINe936
PtbmuW9VEfZPQYYhGoHcAPacU0QDmtqIZtWHlWElfZdRG7cyqP91ZLv+DYBWSMcl
J6UC6Ej8QaS/BM/DL4kGyZ2BeeIBe5JU/VtV2SKKM3jMxfJdklR6zkmFQFDmoUEO
ClDXo7iDbYJrL2jj0VDUY9tSnnDir41D5qS0d6Z2BAAIzRilFYtiuAg94bJ8LTOb
I7ypzCtriNvCPx3F4pPHTD6yuSZJqA60YVvXSP6b9vOqPdMumNkqPVwDFbH/agto
6crtO2p75wQDFCK+21F+5phbHQsgJ45GPHMt2NfrB/ZjxZhfaw84vpH7BOsyEgIU
acCQgFNi8l5Fpq6+Gwp6ihdN86hi1tr1mG3lfQqHvDuQs/zO+DOzEqD8GKjQMq4a
tSeVBWMxumwPslV36uEuYGTQc+wM+Qyel+6uw1QsH5EJGt4b1Xz6zvUx+95MBp1c
c2OZ29TPGNGkf6f2CHE3R5edIXJZbVoILWQGZaKyPwnxNtZWI4cecwmQzmNFi5wa
GyiMpNr3DiO1h24BTYYFSpV4zpf732GW1b5kssP/jWBJAM15nIQWv6BTqjUNxbYc
lLfQts1lBcEJHARL7Y849r9CeCgHngDpfVmKZmxRA1lJBGlzgawaR5GGvJHhF0U9
ZQMaEcL23mkZj0XsIUP+8RyoTTdPYHuInR2El/OaZI4iCBQ+Pikrqtl/Fdm+uPxs
XpHoJ7BS1J9ZSdhp3yUf/FL3HjJTOksoV4wdWm60g7MzgEF4yQ4gbpU12fpiz/nS
GJjw4/T5oxhMoq993rxLZ96RLrszXcQnGOzapUhpKZA3ZmUnUR/c+oo7S8epTHcm
yh6OPyOI82zxaaFGwKMmfOulCgJofGup4a++Sa/UtgUgJmwTOb5i9dlLFz324IJs
gBCE9b7A2PvkAKKPCZ9ibyy80XehSC91dtt0+bXpOcXsx9Hdaiuoso5Bn30gWefi
NUrSCRBX5ptvn6zDDdhVLrKBiLK1QBHiV7NA2BUe4nhdLTpYPXA9a41JestIEbkH
P5320UO2WODzX5Es2f/TLOtKfh9zc1hwKSPevUAfIPScn0bvDORNFXdEL9JLZDqE
WvfPHX1ACj4X3WhLqClYGTgmlg+9FvtbKFxrnn0KgP6jxqMLuTG9t8EuiF5KxMpj
p2cgEtbwD/RG3FeahOS8cRs47/yjXZ0q1DXOwhhsSHnYXphYB7cD0BUZTGg+O4u6
uq7r8cF84xVY+xWSekT0o7Khu5nR777xXsbRhaY9kBdFuFlDhERujTlr6AURc/XC
r9RtFxigT/m6CghQ/x9bFnDgBJiwMy8FAipHnhNO0np+deqdCT0ecmVFOFMwiWIB
E+s6p/4xuO/D4++Z2GEYDlTsDOa5maHPxRpm0Nh3x3Y7Idn87wtrFqAGIkCqvtYt
ZZQyv8JQCLsGLo5xPt8etcsHk2FMutTtd1LGHVZ6pkTovldaO4enIjbQY6C/0y2Z
wslSAx+Kg/HVO5Qa3sbNj82PVXbkFroSDY4eskwazhGW5Edwa3DmP8Tk87Y6ciox
qV5JI3ltVXhY0xNVMvKI+qrQbVIKMxsZffGJYqzFDpSX+FEnDa+h05/l9XMlWxXd
HNANKnE4+061JT+DqNX9EZhlPirv9KuAU37e0tkp5rMvy3MhAhhlZgz2HSZQzjea
v8AJZtOO9v3nIdZI3yCcV7a9zwGpnKCHmC7A/+livlNa0Azy7yqZ2LtrbOIevtGN
3mhKkqeIewiG+o19u2G8FzyPIOASYkRL5RSkOaaVMIHY8kL2WrPXp/zhyZ/cSMIO
5K5hdUBSrS5g4wmwqkVwOdJjK4rs53VT+drRuXZSGaHN/xId31Omn8Sm5OM6bzpp
rXh6LXqgFwBS6R0Ndyij2C9ND/ekp47WR7cisR4h+0+1g7a7sK7G/HRibyQh/MO/
/IxccuIqdExXQJYz8XQcyJ+riupEWNrstvqhrocv5W9C0Uvhep30ldumy0NMO98d
vFS38n3fh9sEd6Ma8+Qn2ePrG1//OY8gphalRo4bYD4/oJncNGHelGYFhFMNxkxc
gFW8614PpBQPjQ30+ME7aGyZJZnecsQJcIgPn5hO+fQ5KuZtZaNu88+TOzmnRGRv
zn/d9Nt90gfDpM322fds1wDZxep9hIIlnEXIw/Ak8Ze8s8UNNQfoYHdieyTyuXbG
0SqK/QFvOEjJGiak3Mpc8GOUl0e7dcHgQcapnTZIcsquiuyVAAEU7eljhbtHrQl0
IVKfc3KLtryG5rPseR2hRiyQzBIZKtG1Y9Oh3xazMpdI7TPaJYOHIAC38cfVz36m
Z4wgfIuosSBbCJ0S0xF34rEngUcVkcgnMn1EN3BjU7pflprFZgpp9yLyKD04SWa8
0rRmE263j5iM/hrt9ONl7pzez/1NPNg1F0kEwMFs436tl4rMdh9Yq+btzsMhJ2uL
VXPPqYO/zL2e7+0UKwb1D6aAYNRP5te8S83jTBb5c2ACMhDkencGcf8ZnyLc0LhV
w64+lBOvdhASx9b/W0cFuXW2rCUHv8PIzqYX0Z1LTUUYCkEua6GpNtMHsPgdEJeC
i/+ZoteTDM9Rg3049nmWaChHraFdsgt3NO9UaGS3oE9UNsmnWk4tS/FYMXmxNQLr
Vtl17ct7BOpW986RtUoPo9hFxt7b+D90jUSMrR3u0iBxf2sALXLU/2CHCuOGBloD
fI4H1x4riycwXTJoVAqBaT+YtL8J7jK4Wy/qRu4OLhC9B2KHkc6NOJwUL3C12qNM
MsAEoi6SqjxA33q0+Mi9lotL6iUqdFyCrnXZb9+WP7Yyrap5mMPJdcAiTsF7zZMd
DnVUtjp00rmi6ZStUTILXH3TKVHnOeIWCnWpemrDQsApXquonsxIv9G2t9f/Y34V
l9r59AgETYxGqhYJJEM4yFJQoC2Mr+QUgcMoSx19UHjeRu7dzIK9qu+OixQVM8xp
gslKC7Ob4du8W6EcnCevpDqL5cOlYzkV23QuCcp2uAcjQJcbVCQTFMK0PhZz1H84
lHIxEC3roaSvMm5QyEVh1i4eMHBOXxXH6rPZp/5uqnX4Zx5H2CXaHTgwZz8CU4bO
dj+79nC/TtolMNf3WHGHUmu0umlFx7O/+I2SM5xDt4TRd1WKorXuMkoLtHAD3l/M
g+8UP29abyHoUsXwUCmWITlVn6lhqrW5h03yzd0cvWXNPrF2FTfSX2aN4PpjTB5R
hZezyAVKOY9aAmuc3TDJHlNYv2SXPd/wmOC7kfyWiSkT7EYg+rzYixp8YU2TkRYY
+gnN7CgRgxUY6yoUCSsNQHli12Znn2txzqv/RYz5RM0tHURwMBjdzz3IUiGQCQHu
3yvqyw5W+j+mkE8tsN6cjgdkRfSUmRcAT6Qeug0OGv1iIOspWDRGlqu7COqcDw43
ucqwIriXLpftR1mGNrBmdUc4Tpq/myPB+kAR0zRC228yMIz7aQtBvbWH+L2+fgCb
4gvFUmiaO59bCOMWeN3HzGnY5yHajm5JTuURW3Ns+kiilVXgDXKi/0aX9l5gW2AU
+t5PJl1zuNvcDFNiZq8DnySEBHuAve3KS5idA71jBkESNH+sZnxbevoVgqa9NTBR
m/E9DxBaiPOn2g8mVLfT7RH1TvWOnsNRPHpnbdizhhEXLHaobQCw5slFjKMVzURg
rpOnz4/r1BFPJRJOiHzUTFoFEOzN5WbakVGwPWPkYAEotnPe/A8yqbvQ+/FyR9+u
M9ZZBN1sRCuwXIsV55wU5On383OGIsHSnUA2nzJ0WM8VVpbvXcMvzk2JLGdeoowq
gHrJQcWkTDcX6JRezfy3+Klaou904FQzYp7xdsp6zFXv74z9JKJfu0WP38h0HlZ/
BK9jRQXknes0P0wIn8MWNHUnDqjwXvncz/DzK7w8BXJSWrDxPDwVUHvqraI4h3RD
Jar4wdTaj9q60klx2KHHREPPI1cFQaehq7MXgYBQL4qCiq7R6Td10Uth8mRqVCu3
ioZURTPkTRpl0WQamx5TKqQkmw+JUQZq0FSOYDDbiZrL/rbmjd/IANQ2i/g/GcEI
xrNHSKIPaaOJG3hVUlNKnBM69oEooglTYGnko52+OXndEKYyZzkfIOiDnBHPc4z1
+92iKZxi2h+50BV0OdPp/ijwPKdcKn0MaRIJ5MlaCgliyJF24rutjacJ4x6d9L8H
Txpf5m2xkuLn6ZdGHB04sqQ2si1s8M77B9jAeOo0OcG6GEtrl2C6/a/2oiehFRIB
9aGcVIOJmBuOSQmx11uUVmjbqml6vLF2nNBWolOG14s5+JTgW6FljrpOx+FkEj8/
EFU09scw02fHg713X2Yj1YxJyF08rEM1GoAvbIHtMwgQ71B8HuVjyXRiA3nAAlRQ
eaZ0uqBZOPd+HNKeZIWVkVTVgNeeOzdWR5cOarrN1mudGTGI0Qv8HVLsx2Hxw6yM
3lUN6BFzVWBnx5muyJnA0/gga2AzthUeW6t6eNqHvXArkqkh5LzeUJXdTkZVuCi/
0ikClAsq/yvFjJ8h+/KaGoR+JXY5EhtPA9cGVSdPguvK/66MPcNi0SrihbCWs+p4
FtO9bVq4TKRLdZmI22kcuLgZ110xTkSg9GNzbOZFy3HtXpbb3S7tS6u78oMbq/cu
TyOVcVbfwHHYr3dQMCE7azsbqoKg+QZA10rRsZkFT/BDQHXKp/TObrTF49jLNLiu
MGGAxquIk35inmfAzEOvs13/EMozq8Pdff5K0qyxECVWL3gD9QDGLwbgCFJSzqN8
mh8SmDQdjL4mzPzXV6yh28xeezMAezYDenpzQLA/pykQBOVfNk0ndt3efv9Fl80R
wn1pgmZ4AgXuZswSkKCtCChvyARZwOtleKB5t1mEOZK3oZ0aljHrUa77xq4QrAKN
se02dgLfTiEnIhgAQSV+27j4HKHwClgb8/gTiIgDQ+7z+cvnQrb+KhQMazSmHsa2
NPRLNaOO4QBB7bsGCFnyQBuBiaSVPwZhh+OBVI2DXFEuY5U0aEosbnh04/8Yu16H
r6C5O5ljcBdqeW7g/va+V7NA5NScGTBCwYrIEQxE2FNWQxM88xMIgrvW7hggi2DO
vtRiSdo/kvbsumti6jc5dYKJZ4OyLh5BmqW4TvgdvhkQZFLryq217ht6hKPQI2x7
HXffwMqWplZRUD/5ml7O0sZ1kzjeXd/nouChoexYbv6aAIiTvZ5nPhsmb/2kAVq4
6HBs11yLfTLcG3WfbZn7qlB6bYD1POvjuZuNZLDL2HuLJ6E4IZgaFS0Y88Tr+OIU
HwPP4UKbuESXuqfAO0115sNHTVhe413i29RYttI8xIImAuePkEyk7Rm1MErHTQJK
aRZs6yzFbibq7cIyZYjfLVipx8BkaQ5GwM41q56sMsK//RzjC9MbzoDVFiogrfKS
T48h3wRHit2SceeUAiF6SsIp0xj/RM0bf3gl+7JArKJAjNnUgX2ez9vT0ZPvNcsg
cRoWrNWX0nb4BikfwflbiHmbra8XBkatlmwdbYG63DAto52ijFENHJUpqPOTaN6N
QCPlRBJWaww1UAM38HkW7avgNF+3jUXkq6rq/1KJRiNJvlXE+K3eATciRMF9NyNO
x4vEkJwHBZVMaJaDTozS9Mq443OuRzorJ6BBsoGj5MTB/oBtJXtph2pao1Cs4NR1
ykjbvD3lOt974MCqKjL7l5cOCoa3QsJ9usE3Z8G4dVbx19LBO1V1mP7/HipWJ40J
NQkViip8rSFSqAsX7Fb+tDiCwFBN+5uHWuSHuOut9ZFVSvvunYVYX7aiZZbSx5yM
PocMPa81EA5JWX0MMudHc14A0P9cTvtBW7Kk1S5OTh7g0sMxVEwUytXXdn3MuZm6
LvBgFNNMpIjK/hdSmFciYWE632grz/JrARAqN3y/HYr/m0eU2Sdp4E0xEBm8y+LO
e/e1O2ib7CqhG6hNCao0OrXxI8w+68yM7DKUi0mffFcUNeSla2WS7apAKiLemR7t
ILQVeWFSgnf0YwjUJMNKPf6pcQseicxqAWxbK93ikN9TK6HgumxRs8VHIEdhUALw
oXNkCF3Fawo/Todi6XTj7TA2hUVZntMI2OLWMYYRJ8NMwCb4FQHiHqkHD2OIH0NR
MhDXcud6ckbP3r1gh6tFtvbS2UFcwk+dR2i+6kH7zVXMPSSvix3wSL45s7wDwdkj
8tdM0w+7zUAv49d/hRGtjtGMIuDjI3z7nYN6FsdPSf+DeUGR/8BpLrxzT07lxGrv
kfAxYrotn/qeeiL4HDzO94K8LpQx6cGddEfaX5kYXWEMaMUxW+uKOfEQXx0EjZwz
MqGe5SDZ8TQoi9C46Nof6NddMwJpLdnow3kM0hEy48gGEcwHT10xTUm6uqOKx5+4
LVspJne31HGC4HR0ZpM6voi43Nz2lsvBKy1iQb10wCF+Jh5u7Shz+0bCRIZ341Gg
fJlng0ZsT7NwVN+i/JjVkmf9wVqyfTetL8wVL/UKc7SbMk3L5eV3uR3ez113tsEI
7fnmP8K1YbY6Qeq71e7FUQRSs1FlwRy4OVDLVR4Y6qEpueJ9fJEALnQy4ry9wYFU
umMuuy0PVkGxiBwaP07LvlrbKAgBobpnI7hlt4P9qMV1zHdYYmuZ3ulnXXiKrnzh
9+6eLs9c7516GBGoxoUYtN6+IYh2qm4DIBe3lnQaRZyjNpfZv9+jfoEF6+ZzLZ5i
M+EroInbUTBd2xAGhonzLuBVTWrluPDrrtpUmrXpj7EZEGKmheVt2XYNG5pzg1gG
CcIy3HSNPmvzvF0lRC8gXIVU4A1osPKLsdBfL3UMM6rDTUXMsgPNFHvuG0tNUzqe
TrP0+h4FpwZNI7aRmZxvWSAnSMHaNHzWJtN/4tO48eYLdT6OIXuxJKrKPd8K9R2b
v58/TtIhdQGrjE5NiZ2tgh9PSlHE9CoSaU9VeV9LCOM9PRF1buUqGglLzheHlMMg
lMP5DIpLUtnuTyrItpGMiUYG+86eh2lMw24LYiSzH7xRbzMb/qEzYRWE9plQ3QZN
elmmrNWfSsjrioMhrWQ/1CvmfKAcv2AmJaQcIgaThzc3n8Ylm9LljjnhfQotnCsE
z35mNnaBg4yrPEVTBQ44NwwMDIXpEaXD4J74hDPyrYQV0U5jXM5KFfqXwgjbUAuF
jfq5jvCekxhbkgw5UboXDixFiSukihP4leBkLYwrqomkQ/+UEw5np52OJwhi8wmc
kGmGmjd208KGj59ox27KUhyuP/TsKhdJY1grem9Rtg844Fbavo8pN0r7TqugPVow
M4BnpqUeDM1+4rAFc7In/6fuJ9noFSoStYobqCxlynbxH3s+Dde5V7TjauDR1xxP
4LjsUWEgog81p3gWWljK44U6hgloWEp1px1MaK9b2kDpSD3w4Etb8I7Fo5ImMt9A
ZBU7F0p2arQw5fS23WNzFC3q7OGmRxrQaH7WiPuu1JM4LQk74vsNg0qk1Jfa7PLa
gis1aOuDWCZbSlnH5EA9ZNyIsKbHDjhaZFl4GjLdMKWazp4omVlHjvqV2cfZ6b9K
ZD7hVr8LntsMzejXwZsmP1kKFjZqRtDrlR+zUUeKfRID6pJT2LWYS309CET9x6JI
zq4Pr+M0rWChFMETjETdBYwADOoqeSFHKMtN0Skkta+xIMq5xpk7zlS4+z5dZHk8
T3qzz90wK+SZw+i5Kxuq4/pFoLcE6pF4OK58Sqve8wFp08pTPnpfd639QZMqMCvb
3LnzYdqTuTxWumI7QQ1iwrUYUNpMnXVJQ0w6BDly8yg6IR8PdnmA/IexmP2uHsg/
kcu3RVGMco47UHDQ9DnKgxtZIsDhpFBpDiveEO4iHTOQv57xfvO66earpVuv3FJn
2weXd6UXRljo5WpqFdjJq6oUPTG+r8RwP2zhRJGO3FU8AHkr+mgccv1asDyAr/Lk
X92KJdITDgivN8gxaNvUFJbkXg/T8nDmMqcfaod1+42ajxVh/gr/M6Be7k4VWrD0
dHlWemE+DWzyQQUFMOLFY86J+jJcyJXa5RN1RmAPHXO6rMIcao4kd+WmBUkE83ec
Ol3XYu5yap3qf6vqMp48Ol5KlG9fpE/UOEx2zqlpxSJzBYI2rOoYYcvQWFFzUe9m
NWAYhT8mIUhQnFo6oyocFWw4OPBfVzn6bzJVJuulFR7LaXpJFiDEn620ps4h+jXX
YDBuCJhx+FDbikCu+RlHsOdz63t5akwhn8of15gfoYKsBlVMSQJY8pBSoBM58MDP
9AGVOl8URAOlfPGqNWApuXsWmA+3Lap7XLcYjN3RVQ5dP1bP8njuuVGldlnMgSX2
aws05kMVzsu7LJjfOXiNLx99L3WaC9DR1gXbekv8vruH28r/cg+IQxIzSlpSeRUh
IwON+ayO2etQQhSIBfSaj3zAkAGi/B3PIbgu0r88aE8IGVBOpxraQa0qv+DkQBiC
wfPWCiml7lt5eR8JcjoPrOpH/aXBNXB63OaJBhc0bFiCBS9iEnvT2bYrCANgtjSA
1o5UFu+YhaL05yeOJfWGl5U0vEoBko1CVXGOkkj/5h61ZIw5NJsV7DnyqF2PuSHC
6V4oJLrTGy3rj6gfplhCumbBClGI0bSUeezZb13OQ0LHuw9Y632QIB15XxAGONhC
AFPagcR4c7bNzCtO04ZJKq7a6RVxOdX+bJsSEAJsrATkRK8hP1LRsP2Rv/SUpF3I
6p8E/aDl4r5tDjh5FkKoVH4glscBaNI4kEVDFCR6Ki2azTQRiLrSz/D6cuaNgNQD
rSk/Nqpip/AxIR5QkVF6vHM6PLI/oKDQoo9QYob4naeX1jYuqCkIsEovBKwgDo9/
UDL5l3eFGKnEWDk1wNIsQqd+W03xwmfLrlppc7PpIFEoaHZ20ZrRrz8XlGJNlg+p
Dinbf199iNjRNjsPvA9pHaiR4vm/+wBVKOp2BCQCeJ/8E3Iv2wRuChNujhCqlraF
DZoWZ4NPpY/2CKuQroJIzXQtbLm31d8Ww9h7pb8G0Nnf2g4xApCs5sEyTqOrWA+t
czldDGIaCNV+dhlFPUHkIE4QRwdLzEOZd3KeEXnPElnvnyGdRvYXABcnGfLdCgur
vRhtPEHF8QHMmTn4AwNLh7Ss3UYfshZH7uO3zAKCyMrXvomtYU1jNg1Z3SU9R0Nk
uT6hXxBTa91J+6/YA/Ky+URDKlyGrEbltcnZMhH1D1mdKwFkZoC5tPaGwFcYf2yc
2is/LuJiIgldsjQIm16ZqoC3hSrX8KOo5rLCl75v2Sm91FNJZMq7bh2FnRo58z3Q
/JeplPDmqbdqj3tEqHARVK14Ria8S8GGH21S2NTnaoIOPsBu2Rv9ifqQfSpZFW+a
SgVAuh/f/uNEv3YTEHdTtEKbGGKyMjIWpon9b5///c78wXi11p1GTCUTIhPEgoj1
48yhDIDVTYINX50B1e/lRxwARLLp3jDbKPITNpB0yKVdCWAEL8+B3cX7AYFLXV2z
Z/1sBltMo6Qw+dDeTOpzYy7NX3K7FHuEklOFeyMkytXelmVZQtW8EkPTP3R3GfWJ
TFfvgaUMpAsnxl2muJLkey9Pjmc1unouaMOL+WDds7kjGNH21puokkjaKTyPVqC4
QJaJUcDN9y3GiighIaOiMoVEQMo/XBJrQeC9oR+KrZfrQWRKUZpMqQAKleveI/JZ
myS0a+Jf+w2CDg5c2uNx6uxEX0dZ8eBhhAlRbMBxLQZxPqDKUz9sfXB6GUKFkjti
/YW7YhexaXDQy9RLkA/jEQ2sS6SajaWwZG9GyvlZsWYCQz7JL1GM4sVGbEafkFDc
UwsYDGY+VofcUOYAV2kNVvD38JAqvlZqLkuJfgZ7SfPZV5xLvBjcVY+cvmxBdhaD
Ctt2J2FVsaYAzwhxNykYh6HRIMJwFb7lEK/dqXbmG35vCyyc9SCiOKR/RahMLDlj
AQtz8+giJxnKqE3B1qpVqi5sm7X5BWz6f7614Dn9inmFIsmpslPNLinpiVrzNlBr
vMN/UMEOKfTcOUC+Em/0TjRgcHlsc4mELBs7ICijTWFID4E5qvgRI9GNJl5rUw9P
vyY9txbyUmOkf26bF7ssT5XHdX6XxGQjLXGa5SyKFJBt6BPy/33k5q1jKgx2yexT
6igL+Luke8WsZIVH9ePG3jmvMW/s1WqLZjJXFzQJNrKXEQGVsBTbHenTtiAF8xL/
IfujYzoL5UvnvJedKFvUTfM5N2inZzsy54bQxaFARP3X3FTw3u6ITeWcFT1RLcvE
n3H6qYqgXaWBIb3Xu49sL4jbzocV8pXtE41f/8Yn5UndweTSXt4UbK47JnjNDA7/
ztY1XzrwRECekOvJ++KZvG113Prz/j20cMZv7H5BUyMwMp602lvA5mok1zrfyoc7
jsNdT/Z/mkwGQliQZgVkF68+V9zdiIUjwUV8uxscktNaNiE9c97z/v+7Qe7fA/jV
fY1quN1XY3PTBLQM7v9qXQJeXwkXcs4iQKjtQ4l5ClCuSfWl4fpzoIcn/TfSJx1V
PL6hMCq7/kV0ci0SDDPn3aJFiV3uwXH8WSHmeHCC++VI9eGwf+7L/8HEwhIJ2KHs
DO4bmH1xERG0jytzw2O1iIc57BVG1vwWFPlvZF8Im/2Eo372JaneoOkj5odOW6IR
pm4n7Xma4gZ/EOfUjLjzpOFlQvBY63aaejfjKJor8rIvUwKwY8w1Zl4+4qSs9A+R
Wyt5R6iO5RIGuuCFpYXBhSs7uPkzf8Er0SFoT9fnFzr8qB4Li/OvNdw/6L27gOEd
yvrKxlZnv/k9SXAnUN19Hh9rvnv/EWHJygFBEvHNxQT9jaHx66dURPvDHTbDYL+0
Idf5kWuZl9jPCZQf0DdC7KRDNXDsmAQ/KaVfnRa/gzSYEgSNpc/CFFHg4mV1tf0m
g75RVbHTxOc/0jaX+OkznhYXgTqo2s93dwsIKCrl2DLQnraf7GE+X7bQAT3pgja4
3tnHjVhAFJ660ZdpQyxtb3F4VKz86v9PhmLGOhOvmJp/x0lGJ8EoBLFQVpozTwNX
avHX8ERJSTkDK+miXx7XTjy7xiYTTpcc1wKZVMqZKSULDwl2SfzF04A63KsunOpi
80INwi+lkye3KI3POjQcC5lf/0JvC9bLD0bE7Zf3gvA2MMQ5QsN33BgEc9BzOGQ7
fm3Sl+pdhYxEkpB0wrVjGEevdmvEdbzssXeEauWFX8eB738bZKQqXeNAuADyGSh6
P9/CYYI1TjHuAhUbFQxJJdxy+b4U2uSTWanikQjp0zEVsyEToBp6NgV2kiHYL04O
rUKf4xFxYHVYTElqd+hGvvjVFr2FD27l8q9P0jfRDj1DgdIAh3HIPSVL0u0AEqoG
TS3y320rUiHBM0ZMUUfNMpPXwJ2fsX1qjNSg/aMHQ+WZXyFyYv/qROh2lzpjX6aX
o1PmMYSkxbNfpBtGMwerwzVwXBAy3oM5jQrt+zlthpcoqro3lmWXZrUe5v3bMP/m
fsCOWfN6nnQH0Z8/byVZTcPQARCky1l6r9TxPKnqRr2u7BMUc34xm1uM7fwcl7Mc
DWH32Z31b7ewKr0xCCgUNzg8oZoL+aM6wU/e3KzOJNGNsTrMZTxarjQe/xl7Tk6D
GviIaxj27yP5zTvdd7c3drbQ+vQfBvCPbQDIKWFLGOQZFh30UkeTGfllOYKJL4BI
ri+sZrIr1AoGUOl82SZA2SU7rBpGQVoLSUsn8KrBiIQgrD9ticT8DxUelCCEOA0H
WoKMZ1chRnbRIwqIUYMamSmFH9RkT9D2tn0FwpsERgOV3REIOOhsTJdRZvCP62jw
rNIzFAMC6xcUEmiC3RnehrtVDYspMbQ3/L0NttncLwCtpKdIAoxpsSSxXmbPKLmN
F5Oq66I9D8aGSN+a7vFrmwD50oBo/kLW/glR+blnuP/Pv7yoA7gdSs7z5u/1tkLN
xAra9k+DF9Wo0SNhRUYM1haenGrSUp1C/J6CL/8YoCeOLZpDGsIjx0/sqUa4HtR1
hqxQ2Twq/Bpw48P+ouSuDvUBLKyy/+JbG6mDcAu399WEjUT3pMLYsYVqQTjAgm3r
5HvcuwBJN5j04SnjhLXIsAjosKyvk9WUb5grOG6yH7Y7JYF4u+nG+s3/wjruhmvk
t/DlaKwUJYbmKWFWXB4eprH0FYb7joC7AoDwHHoVy8hs3bYLZZGi1MAC8J8gXmhe
Z1a3n6BcH9ju+J0Jh0xCQDBRUbdvPA9eGcbmYwrO870x3CbrbDZjnGPcDoeEUtWr
vQzWJ+ekXCYCI9SGQz23LmoIW/126vnJInRvF7kwj3Hdpz80U2Uwug7Elmcb8Tg5
vkTfgGawSrxlt5QPCxou4HAUiKZCx4MzgVvaGqtIxFv5lJVhU/8kv7Op7H+cvTZW
8veNEKR5LPPFoV5R9wzXnxH3XglxvpyQsP/FdA1qijLlebx1XlWAZnyhNnBE4ZYv
Q7ah1H0hAJNq8Xiaj4ooSa6X1QEQuoFEWEIza1z4Yt088s7CMr1Mt41frBJThxNh
hcVEkC+6zsWBKLZLuB0Ljga3ih2edzn6UP2d3NNZ9BO7lh5VGMIr9yy4oAuHAFJN
7xhPBbDVs69IODyfn8zKrDXJToRc5p5WfEZNcpXMEfK0VRO0b4f0e2kELtxdSIZ6
zjM4AczMZ7MLyPr0ayERk1LrvoM1pEcq3z1jyeRtbNQRHndarXcnaNQcAvkD2tVH
JFYzgCfszqOiiFIpcemD+bz8I9Ga4y7oEkzoG2tUZi4VXwpH8ImrPAjItgP7Hia3
iFYbinIAVnqkplvpDeQEvwMskwDV0UVFDDC11/sI1OluDuvka8ACHpcNKCDCBFNA
0bejfXaINZZiuyt3wBL90X3GcO+ZzFZHLbdDH5RLcMas6OLBsMP9hvDHZgk01Qny
VAJR0McDtvjqJE1AzTRPhm4FB4iUV1yiU4Gn6r1njqMqxA9xb3tl2r6YCstuRuQo
cPTuDgEbNIg6vpAgEW4Wj7WxZUFo4fk2RkrO2sJOOsnfOKXx//v5v6zzX6UnyH+e
O0Qcl0vcSKEAyJwzAkjGw2l0ndJ8ZKplnD5713jt3xMErUH3BucnJK7mzUiMIpcu
JdHPCw5s6SAUOH+qeHcHiJ8/5LiGVK1pkhv93g01mfmifZ+VblRR+Bgr348gm1rD
2S8n1QwoBXCghuSB8eVz6fAdjp0EKxVnJ+rJO6M2j8vq5vl2u8TOcqbZCGO0EqwN
L2jJ1yuG6+zB4n4y73IyXU9d2sRsZVTOm0ZcPIvpU4slqo+YH7txgjgChDMmTQbI
HBnS16OoBHUCQ69vSfrNGsATsN38+35Tatzz0BWApG789QoExU/hBCvyGkxz+36n
X/k0jxJvHvU/4xa59r9Q7M1MNmKzBsjQwfU/ed7TBOAxV5M4mj6zYma5z/qtoBod
eyFBRriOjdgBMz2MGv3thEEf0GY66E2UMDGBpPpdTMtd+dNNiBgZP+ysXJ+a2691
sBSXS5a5z8+bc7RRKSmqnx9op0kq1A+YgH+mYauLIaIKYIC8fvHnuAuj3NM1cquG
zw5AuPCBxxYpOdh6DP0n6KEK+qIe2P995r75UdhzAtwfkPj4QoiOlqEODKJnE0Sm
h+XgQYsIaz5fsOKIEI1zgPJf18fAEggSwacujAkEWAA3TwkadL6Udq+lXGiiEeK8
hFnlb4vCeDWnnu08HgbFEZHl5UWoSYVJPHb4ynxz3Zac5M6t0+3hKK15rtcqTvId
bt8yyz2JoHpAG2q0JUYIEGtQmUmx1PFJaGNw/wXYL663NQNRcD05CvHvAQJD70Su
SplPgwstrAsB8j//lAFIGXP2miOj/dcGBjCpbIgGRQUKUCsddRK6uYVtbmfgFuTB
FNhtIzjlGoLuBc2MkIvL5qNdRpkVwvW8upL2Z88dwN8PIIRTGrPyJT9ofbnWzIz/
O4I1aP58ByH+Z36shfKVCDCBIZZ5S0NgMeNpvKCe8QPIXie753iHJ3Iqt5DAs38l
S0ficbw5HKivWN4y8anPa4C3EWX7MMZWTsOf8ncAfut8YeavBb9WTyCybREirTCE
WBmPgaaY+SqmhAgFwZhfbT85eLotf/z+8BjKrQce7bMyggcx1y4brZLB9FSNJ/Q+
e923129+zOmNAC5a0W78tYa2rO8vc8tbJxXH4j/REnyLdnf2hlV60BbbP5NYQFnf
vdFr5YZGb91xMoY9QimLPwumpZKt32kL66q7Dcc2MhBLNK7KrUlsC07S/dEJHukg
0bxL2kUTk5JAJrzeuUtWjcEByP1LUNPofUkoKd0CtUlHC00nfylKzGfEjg2KsL8B
tfp+2WVv9f+ZGeMuFbw7/7WuTKu0W3Tismql7nV28xTj/NWVDGjtf2VH8u4J3s93
M5zXQyCchZcTUSwqs4P8qnJ7t1doVCmG5HzfHFDMhTdy3qR+Ryw5BuycYwTF5//o
uTknxEOr4nYQVXc6A0Ej5VLPAOPeFGxVyxtAaFNqQY777yoC5AgvmdNmkYBVMgqB
pcH6YIirRmB5cVZdTj7lgZTRZ94AmE/mKDATwN3UEygtQk/nNxWSwKx+N/YHL8a8
MND0rAL1+1PUdgUYDxxuBVzLVw2kQ4g2XiLryqNDrxc01z2xIk5aSL/Qm9H3makN
KQLyqwFM3rRBvRMtPCnYpeE5dAS36chINCHRmaxnDYHqmaYOoAbepE+21YzG25th
ZmnhvhO45MgLjvdjXc5yJgmilAW3jvsqm35S+ZsEMjF0oS06by/E0w/4cg00TFcB
dN1fF4Cz0SFsHA8gNoWxMFy8t3QnqC0EN7FPA/B+wR2cOZS+Na98xRY/iYnH2BtK
exc6/q5aoFQ2kMxu0+M0if/4lh0qrGvxTELDK3SPtuJzWxgVC/Soo2nZK6/qtcXv
4m1Ip89P+AwN1Q1n601KwRjaxHciHRaakvwHjq5P4AE2PFHsMvJxj8q9LhfxvHgy
3EydeagPmrqz5zNZnG2KZiSI4d+Y1t/4aEMX6Lwu1LPp64lu/+Nvb/envVyHGbdx
ZNf2SdC1h/YeOWf3bJQrCLQZUCECEMH1FNpahD9sGJ2tldw/AZs92O22gJUNeIVr
fS/EmQwf9/iscC6WTM5YyXQb2GKy6F5kpj3wSp40po585QbPugkkm7MD+qfzNryZ
FQ9aNMuKa39gbW4p2fxWgX0nRE3w+vhs6NnUBifwMkUUo1qkPuR3T1NApAVP+Hrn
mzXXAga/o+NswflsC18X8V8eExw8qhOQOnqZ5LybPszYGuZ3vjfQURGQ/ciGzyNf
RPPaPJu9GBMMLpz+ZqNUaaoA0N2TOC5rAoorZyPUwKe7A0P3w5KAoQmc3Erglh+1
jI90t6xwInINJvjII/1yZtJLSAT9/QXMxEPdsOjQQezfbwlMz0WCcV6z1LNvRdLZ
uoBVvKeT10Z+KPnKYOuVSJVDveiwiU1zyFthymXTyU+STYXgVjm8yBSqKH1ApvRY
sQ9ijBE+9nmaDl46EKlZo4KfxHqTJcbKaa3GT4XlqXETiy1f6L+gCGnmpjzzwR3Z
dTX3lB68IfidNwmAdpFO9g9HkXFpEABJm8YY8t12X3rjHyFuqoZ8EN5dqbjmfY1s
TNysz8ZSHDlgNFt4KH3aTIOBY1eCDSifztItKm/ZokfLMeg2ZdN/peYRcf2H/G+Q
b9yCrsj/GzswOKYkWaJAPg8Yt0KylGCY1Zj7Er/toHupEtZXHzp4ojQBUWy5/iik
07JNyxU6seNe4Iey6ydeWcC1RgWZ/rmIOoY83F7MzRJfa0Oy4+H/y8ZhBpFhQ3cH
c75h+lXygH66+1g3ptaqSsSjbaDbXaCjp3XZ4DAiUOWHRYcRvu5VVpqFH8gDLvRL
tb8Qb37EmuH6iK3xNepoq17vvryYNXHvXLWTgwAj04dAdLacIB40oATfam5zjtcM
YI2rqZgJtl6KGwsN3ddNdiDgfgU0AVBTyyiSr97ygWjp9zmOefOkeBCbbR+vORPi
QMzGVtrNqoAQVdY/mqph4YWmQ1tWeILm7FTu5hMbcKEo+hJ+pZv21m4wadwBAxJc
iSVVt2BYeza5NfvoU3pRfCKhZsO8xXk37w1Zyt9W9ivTPlspRYbzll29yJq9AX0x
jIv+66h89stIrHhj39axQI4MiswldK9rSc/ipbbnZ5aLJG0xA3H4dFKBDCPf4tot
puQu341wzNRATDDE1KMy9GoEdhDfyyoVD45G+wFdwmQlgGgKENzsy5MoSja3FcIe
kQmVnOpItpTBs0D0VDuYU+jfL0Jz5kXzDscE/ZVjy6mbs3NlVPJrV2McZOh5qtks
QeaZUhmpE/CuVt1Z8cOMn31OWdd2lT+sj8qphZjw0F2WKVF3KqrtZfF2TKdnTqms
zcnQm4DMW95Su6+V4gV6YJkkilhxjvAKod9TN/IyFMHlHZOcY7ScGfnK6TJsCi7z
CZABhpDFqbRW2W87zlBf5mrTkQcBTSQETFwE2FFp80egadjZlhAsTf6WAKrGkeB+
s4OmPJaUsBmuCdvObx1ZyM/q6NnMpFJdJD5TjNRr8w7tU/F3hnhuVNDlurYm+QfR
+m3bMkwfchXvXR/mKpussaIEeLT7IsOGUv2L+HAdZ52v/S8meHzjGXZPcMbqHfuC
w7n3iaOaso4necz7YF2ahdQMZZySFP/3NbAhqxuJZQibECC2s5iqWSZLkaEBnJhj
MfhrWDaPdf3Dwejh5brbS8rjt31MTk8lsjEoMJ/iFxDZpbtorKlM8QR6CErvmZ7q
YGCEE0b62lgAl+YX7BUwE0Lk7/qVauRis9/Ek+oy/94VoX5InrLoTt26f7HwU2LX
j2C48FZJo0oBRdiXH+glqTNZ4tIkJdyYjxusKxLq0uIhp0BOqK+W5ulY++n6WhwL
SDns8wVDvr2bi2ZmY562ZWEhgg1Vnz3z5dglNzUWl5BoTNrhMF6SuuLM/S17HZjE
4dQ0Uk2CfI5Y5jrzBwOfdD0DLCrkov5CGTigIdoS8CHlXm16mgRuA2UJnopdPb6H
a7QhvqNZHb8EahzPp9PRVY5NPmf7GRjuJmOTg5CbqscRpPZ/yWBkG3D3DTdLwjrA
MRBSCP/I+HrgbDiYs4NeGl7Xjks9y6DpgpOl2GDgZy5jJbc99soSo8Q0AfenCsrJ
aOqAfa51SFBhlgNQEbnNEgMeP/L+WeoBf8UaLW9i7ZbHW7Y0NIJjPvpVvSx4W/xt
I1S4Q54c3yHvKqouTv8y6Mynx315u355l0+nkt502euGIo+tQkRwFD3sj0IPB5zR
/OOALmvtcwRxB1FxX2R/AqAZ26UTeTZzcNRpZNhVc3ethdAOJ4dIZhD6aCRBsk3g
wstiiVCQgZA2AQfBNg5qV6XfYtwZAd6CWnGJxaaYkjKVMjqtAcLXzfFsK4dxJQ7f
7D/s3djx4ej7tZLS1W5HLHNz1nNhV6bgjC/RlsBwOWnwmepQh1HyC3uKvzWEOC4P
P0o/7addGb5t+EVoPah3rgKzqeWrrKKHeFtSQDj8eBTgXPy2BYt0cNgwmzSOxh3b
RzqPr6Lll8U9q7DbsyIcF5VU3eAs/AjhBCU2rZe1m8KP0jJzwXLlJ1HrlES1aTzy
BNS5wkFzFoeukOqIjvdk3UnuZYMozpz9S6fNSKAP0PYQWi0gQfWK87tVNo5BjPc/
HR4p6w2SXtA5UqsrKdaqDThFrbjCvK3rjCstH+hE1+uqN5NaMH+7hBY7DRByOAPJ
DA9JLTtkJVrsz3zyZaMXSkJjzGc0Ush0Dt45DP7+S2xKgWRcTWS6lPQKMVpQ5gmP
s46ndDg7nJ1/v4JN8PzQ0ZMErFocmWqcQoKPUVSnvu8e9Kq+07TNqNu0OAUk2oZx
nluTaYHWjjtAMMe2CDZVl8XenIlbcU++n6sPD+01OYKMWPU/MZPUYbTnututlUHv
ovBBACS6xkX6UxvW615xftKMDHR7J7Kgi2hxNzA5YtVUbGafHuNaScnyjdIr/LgN
MR6HplfMmnXg1B6zrT+rAGq1ZtP6BdCi022bzwjLQ2epw79l37lHbjirKWjRgl98
GlG8UesNj/mlgB3uAyEZMGC/xeyd0vG0Rke3zW9VAITvFSkcJQaFSefOdzgfu0FL
1tDSuGgshgwPXsV8vXDvnIMD0Ck7CP8obVISjAZKc+FXR4lssKPGpoOaVlpvX26a
NRBVom7ap3DBwxP/mMKt9LjvG09f5i/sgNOE0TTcHVO1Z6Yn5sbjGXua3KAqELfI
cEUR6XrWL4XS8CVOOaRFF2laIZfIhpbeurZuDC86vspn7xPxt4rMGODBTpnzSdGy
0vS4OMxWKn2pzmF1ZzbdpyBMRZ3Krb5IxUaM/xEtqhlDdrSuom5XlLz7F1n09K1P
zMfwyn4WTOJfaacQJWUzsDoMwci4FQulWejSMiFVk7LeVPpyJBvNRnpAeAFTwg9p
lcYq1Ku5+2fHF//7kWMxunBMY98wC8mGKeuAE3sB/lQr6H5ZLR3MMxkecWI4f7b8
OKhVWqXeSGZlS3rRv7eZ9wEsaxq9AiJZdbQCBfm9zxv0zynfcwPpRso4VBuoEYhA
SMCONPw3CEV3A1cNQFtGPUyxGc7/bbRsTTnKgd4c4fpfIPne2dcvOIaJ3N0jNqVv
bpMXzKQRsyV5M6/BESgfzgUyW935+7kFhkb5Z6eJRXbMlqSmQoxFIrpZz4shNFtQ
35+WBCmMGJO7TeGuhMqF042fEi9DdPSf0MlGWTZVpG6LdF3/QhPsq8p4WiHRZnKe
cMA/fw+ejddIOZuAcKaFbgAC4vtrJDWmWaxm200WkOIkh9xxRtcUvHB1a4HY1CDn
+/G9Tpk3QFHg/GjCI92xigRUgVZpOAfqqjmzRnWfxEQyAjuaZRREZIPrTx7An8vU
RvWrZr1HU616eC3XG57XTyKyABb+FXrGuy9sZF4awB1AmCsIw2+WAcODuZjbvElg
aq9W4oo5yUmvtZjfe/7INuzSrutoYtMeKz9fm+mcHJyMkv5x9U5ze0qNcRXjJzE4
mik1F2G5re0E/0zN4GTuxWFTiCsbBn61sDjrV5bGbe7z1N4Xmwbv74ilphkisVO9
nLnwBZr+TQo/KS2Q73cb57pPbyu2/xWhP8Am1m413vvY/c9yxYn+sxgDjaxLiO+W
noGg6XBsfTeQmbDxBJAfIK7+rgVJLEhuvLiFlqSLVLvKFEepTiFzbQnGElKABI8q
3IeE9DqWYJ4Gfk8jVQ1dMsUScNwtFt2qkF08L0DaFg3CLPfhUiPw65IC+dp5T41N
XR88ozliFFEy8zjVWFFDtElS5yKtaHdiUe867/RqcJKFDm8KYEm77foMeAu/R6BP
vYDW+XamPc/nbV4MviJyuVbbCo+H/C2dsyud+ek58Tor2O/Z9VWunLyx/twGr8B6
Yb4JS37P5SfxGefyz6NXTQyBqe5lvgFJ2ddzR/rhZ/xQ8m26XM7Om9vLvYplB0rQ
qxYQMNH172t5EF9yLEJ+np7IvJzayn1GsxqUMcOlf1rDNzdp5p62g76Bh/yRfAmH
k4rqiF8M7nRD1eXUL4AK6t5pqnKS+ger4UKYkqB5vNkQf8HC5DjMBlS4HrMHJoTR
1XRT7+35XGe2ISEClLRazsFSoRfRnwoQPFv5PbYLsAi0oX25ZgCAw78uUSyh0Z9c
k2ZO0n/xd06bedEF4nUtco48NW0iJbeqgYzm+EiSr7QOMCj14cSmQfNGSEpb3J6f
wyhV8dxo0LrY1BSUzsKL7USzGqbuC5cfem7OOiezm00ca2nDYPNyxYIZgrz77Mcd
vsVfTbw70+FYMUSwIsRyiLv7J1WmChyFCM560IdlinR9p+2rznssQGh+wpEcDU6e
TNkFMjHmRdXuKxCdo1jJhF6v6XT/MqzjgtKO3jvrnFqQoNRZiCGpJpkSyRy/uXdC
8d/dGkGbVnMgqc/smYhMgQ2I2whyQ3171UxV5OBM7wAd+JX8JqWKfmlqtmbpaLPn
fJ08AxGMpgY417x7lANrsQwdudjsJG/3d6k91L4P719JnDVY1ZKE2Qw66mXbaCX2
XDHDVz+28AwhbhHyGhuawPtqxkC8W6Hx40mD5n68TM+K00hoHxD5Q1sOKtB9R9GY
jpCCekiREyHozq/fd4AUdC2SmV+ITaCXct5ccxB00CnVcQ6vbrJSTYRkqxXCV3wW
kpTDAlSKV9eGOx3j+zDP7bnc5+HhzDBhTNLUZR+qC2vdnNMgAKs4cyieGn+PlkzH
KUKP2UP/a+94l8jMUsDV50fTVlJS9KcCSSFMkmKjI27xb3BIiA9lfAfP097Li+4O
5o90jTH/YwyScHtlXE8kwHrimLhWLZaj6yPWgH9z5wiYSKICvrpfSE5VnwjJUFeh
VKYZS8k0xWdcYQzDtSqsyTmASanynwrm765ZCp1na5Dxa3PJIlzciLGZHjVanxVb
hTi1Q1CJL6b/KFLu38J609Rn54WWIwRIJUcGKz3V52NzNFUv0/4IZO7rr8teI4S+
uhx7ZtwTIWAJGD0Ac5hOLrttY5Xzz3AG63OHlOsPk5ocN2JHRyC5ehmVxRshQfGp
JEkrKBgf54XDR9J4EC4/UCGNiv+4Z+dlySte+ISCjsqU63n0JBoIxYdLIVTo79Kn
jYUnxOUW+MHChSY5LDFwDnM18cQ3AYzplhPbtsgGq3QxFLx9CYTqOpkmddtJF8Sr
XyxH2VdwNhqWfs2ex1pGil0osp1Dz33y4TdTDkv03IO4p8M2zD5jqJMd8CFi36/k
UzubnG1XbxuyHi31YdnPLTxm590Z4AAYIBHVGeyYanBZiqhRJgWS1Wnxbj8VPx/d
mpE9dQLlpH5K/SwsfuDYQYnE9IbEYswOrXG+1RAZhA73J+BSw/Uy40yUesTx0d91
EMe3sj6irZDONShb20EQWm8zoC0aDneDOZV/tov20UXz34Mw9SxXSJz014m4MfWN
JnIqIRAYlAi6xrqodrBk0pTaWcIt2TbcwdsWb/ipC6LfQjDCPUEo5APzuYSE1mA+
EHRd7sa+Z9BgqVS8681Rhd7hleZQ1g87lKsEdSwS/BkFugpLfvuVdvcsmoLX/kqD
EA/p0tFsPzh1LqNRoUnGg/ln4eqE8Ae2VZpSwLi0ObSzaFvBta+pO17QTp8CV5E0
4wEfmmB/fT2/BiE1UChbtawqWbfV4sN5Gs8qSYcbR1/5OxkTuk6LSxr3o44TE3og
UuD5lqoxsf14jspa4uLC3wCX9dtb7anx31sdThLfBLq7ZbECU4SDN1SO9dfH6kTS
fOh08/FP+GzKtPxUFa2hTmJ1coOq0Qy09SDwekvUr2rTwa/QZrZIf70SQ6+HJjux
nwzw7qjhXqE2KLyQaAqWOd7r1thXSrygzzNUseeM6OVlQdzBZheD2ob5u1wqxrm9
Y7N+RELu8Rtlugr1jcXFS8YsTu3xoX1AmvAEj8VL9OF7RsE4UH27SyR7PS61kQmm
rTUY2QaIoQOiTXJKjxZURSZ2y7tmWA9snJZueHwE2M8V27tx6DK07762Xl1MH9Gp
Z7AeQN9jcMAWSGxtovb0Ru0BQVEpLhJMGzla1ARasTFWlZmVBm52fVbFjQHXhi9+
OuJXONBtynE2L/vmVm8Pntjq6DTnrbAeCWIabrHIfIEWvRcS1PSVn5HLNIAB73Q6
cWGTrnsYrxWKBCW0DIps7wGCokkqKhN+cQ1HGXmA+5EC4CZ1mlfd68Gxzu9jLBB7
YgMY9VO40hoKM9mfJPwjw8tSu/x8A2E/sxUM3jB8jPerVXBSxbU9LXFid3nmTnfj
+uhkR00HV1AVc/RGSIYYkQTU3YFPFGpxQkzYxUPPIp9Zp4/9L3YuLazFkqWHbBxy
1uRdtRgC+/tMYfh1v3OdAhHb5gqRDTyjxSl3H+YqnDCOREX6bPcaxH70s/m4uhQ/
uA1kw/nDRCeARMjVVsIUpoySb/5Vcc0VOZHSfEEF9FM+LjqonyfoaDIIxwaTG5G1
S48TLgZ2kS+9oPOx94PFs2BE0j8OIzxV+V7YMXN08l6gJV0y1AATJ6kPMDagMqtO
zAk4atlE/283PGSKns8nVlFti535xqi1rX5XTehLay/3IWbmxHRD/ETlzVQAhZ50
ZEHilAJzOj1d2pHY0VjKJTCrTtGR1nCLPp+7/QWhE1HK3kaA7M0TAOc4dp+kdlrc
ePK4TbXc4y9U5bazO5iBLAh7+60W1QHTnPTrnsqRttbqksG8wBe8Z7NpKlSXsJ08
QD8Xdypz4LV60+jsz5ClIOhwl6Sh+i71UOkHMwSqHMI4UO0qk7wW67xSs2P/VP/H
rCYHMYm1dFjHsKp45muGVa5C2h8s/EZgSJ49jNo1DbFWzU+zd9VhOod3nQnwQTTK
Xjm7odrNMKkQPE2JZhhFZ9OyZqQuQNfp8aE9hOtfCOWd01O3TDTkMIWxXkFoNiZf
idm4pnJ9PUiRJsQNh1Z6mBiQlvthlGMyVCCnR390xE35TCIrM9ZVa76V6nYeLZGh
/8NpgBoZbOdcE3801bsXZuQAevdSVB7J1ZfXarYQ1ht0+tT5DgspdMciGStWwsIL
yF3nq9Vtm0Z9ZCkehXbcFmR6nJKhf7UNMnH0Fz6tuU8+E9zUhabwvd4teTGoSCDT
7Np0ySx76EmnuAZTIA7OCoA/GByDEnxzEckMqdkkVSk1PSucc7/TdSMfrIO/QeHR
uaYFO/9QpNpoT1DnzUhBvQ1irR5VMPLLAoGcMDRKnEq3aKj3/3LXJaCUoFld+7ar
7rbyuqCmHXm0haZI0Iz1MQvl8GGTHBajhcVAKXBqxwN6ZgXHFMIIQPjwb8JMlAI5
3RfByetUfB3NWATGqqwy1ZeUGIcAQBTCWTJJTMjldQRUhyroKuvwhPAMd1Nn3Z8f
o981gxdOUVJL4AiG9nj5B36+DKrtOvfsS3eF+W9dCC/a0VIPFd6mrHrtoHfHNXZT
hfgcMy4yMoKvQ5c3t5aWxwEWMQgUmpyQRAqIdxZLCscQGzmosjo0cPVVRHJzCe7I
apefNQ5XapcHBD9HERlhLqS+vJIidOJxShBb+RZAIl6x9beU7j+ztmXkArdt65XH
02hAgpxGppC+ZsYiXB9P5O8EiKGqgdklen2NTdoB658Vo7Y9+Srh4sCm8aSgn9yF
dZFHXIIQ2E+szGjbbaay7HXXE+8LMFltlqqP23EW/YatfpX2JuRNIGSmG9H3W50L
YTVbv4R3N+L4EDPzn+J/u65Ra1oEqvJfp7cB+ER7L8hyQr5JfSJojjXdF0EZDwRH
Vpxa0QD3VXJgkMKOBVNHL6UBCgnkUD4uPUC8/hzpJh8kqAoU68EIAIXAP9KPKucG
R2eVnjF1Hkt17hApiPveHqjRcvxFSmW20D/x8iP/JX2FrUH/3c42DTAW3yguyjKj
8CzVb104aS7qgKxnXo6t7ZiGJymfwlZi+pqJr3+kxpLjotZIt+cZryOSRWQ8rv+X
AO0ak+lxZm1LKfbejKOmQjwal7WoUdoj86tvMZB94yC9WT5k3PQ6pC+dutZOvbOU
dMr8xYtJ93rL9G/OuQrq4rVnC6i27TbHC+biiZRm+RPnjHoRrMf3ZWXr3HnFBU3M
1wqm48CMH2NbhUVl3Qw9Juit/kvM4ASz2gSb4YhWNjeDe7Jo0YXi8ybwjV5zMqqv
0hzXEgnFC4KhQR9W9aA8ksYDH+vyxGNxacvC+9U3agx3igDhvRIbfif+edNipn+0
bZmmxOKOrEhlz7e0IiCqzjzZlMfsTHDwSEnpcY+c/4OvFPLkIc/gTeJDCGJng6zf
ThSNJwzGYxhFPy07ikMi/sl59CtCXSYQsihlpTIph4HVpIP7nLImFZx4y3JliVzD
fyj2JSiBOdNGxYoBCjxARP63lcUdxlJlfAhwVopJBQAj7kEpjGjVTQENO3DOvaL6
BTajuERFGPXh2NsO/rOVSFzS538btF/J0crdG6FgmFAabf50FgMXCasWTZXTLPKd
Imo51AhQWIloYlMwVY1JfNs8nZJfRFRcefc+25c5+AQDkJkMLw+47ctpW4BRKee2
g6TY2yWOwNFTRFOhWt3hQBu+sRzdGUiRGsYC7wO7gOcpvMLfQLIV/WIWSRulVFLy
3FDLlzpW9NTPeBeioAz7nBYDoG3ilk3VuTPVOMKxj5K8enmgyDjtlKf6LzL2VErB
kYdrYTew+XAk1k5o/46AmV9UvQGwvuVGZOYCdOVhknsmVgz+SK1oOh52LAqOZm1K
WEISgOM81t3RwebocGoJAfBHkV21vUEkG1wSmQusOrGD7c5LBPWIBpMeOYf+6ZQx
AXErb1Zc2ji5kVu3pwcr9PitrM8hDTPj+jOVdlXQCPN9/XKTHQAtAIC+y0RUR8/Z
5iw3daGpYAX02jk+XKSCHKQAg44OkqaEhUpzvoYXd9DoIJsLOIvclZ8hufX68GCf
2WY6KU6rJlndpERBfND5xr9IE7qJ4upqdWKZaei59R9nISmMvi+iWvIuBm980emI
0j4PvSP+GtG52y2nxuc83w7sD/q9XclOmcw8YS+7YHpNmPzQHNppEVvTJGTXwtlo
dYZGGz2D7kXdB+LPwhcU8oasiWBAh+dn7slgrFBHHEVu+YnCtALmxmgsjtX/E3G9
jXxo8voLFkYMAoE5NZaIvAtv/ZP2QTg7bn5jfNxSuWnV9cNrgaKtkE2NRao2jdFH
Wj0VZDnW+vMs0544gxbrTUyjATc9St4Ro5pZJXrNdqZfYxPnuxiFMQl12706Topz
xJUdAqtk670TVzbKogSzt3KJ7oFux2bmBPb5RpkC3m3AII5wgLwrdpQMy4FPF/fj
dn+9NVoen7Qu2UsHzJYtwiH+POILysdearTAlMFnPk1qEqHSt08fwZZ9pxYEipIb
1f8GxVUj7Ap0azvUCfRX6R1XzxQbpPt5sT8Ca93qrmwA/zhMSzAYKfbA3nSZmyz9
FHWPlka+my/3+Y1Qinn7DZaAhGkgXhK+V66Cpb7D7GrJHnk3yrsh9TRsjYFpihb8
5MZOxczX/k8G7Ak81+av6ibIB7WRjnnnaAGKklNqyluyfiLyP3ab/F2z290F+4KL
i7K3p5UICzLytFZelGqd/usDI6/Oom1o5ij2DY3ChHaUpi3aj6RdRX0S+CJZjbwf
/E08Wc/VXjJ1twWAJnv9Hqsy2gLzaPPkuZw4MJalUwEEVhpCfkpYO633tsts/j6M
vcoWpEjbtHMymb+bKL7aiYNcb/buQxsK6aAaWwNQsrQ0igpCaVtkAZYdQM7qph1V
QgJNtY9kLHi09KwXYB7SXVOco6p8MgLNJGrboW9cTcai661L9BsFaHTuIc/VQvb6
skiqiQqgqT7JOucS4pqspzsuj9uDO3PgIJA5qbKZwjqkXyT/KRzHP3g+jI5oXtUA
YcW/qc5O63yGaxbu7Ob8UxSL2R8cIrqrhLeAYWdtTigGruvB9Pk2g5jOFEbhuddd
uH81ybP+JzUMWqHGF/7xjHM92ZBaNAKHDBjyjP46/hhF5MVQI8t9aepDsBBSwmU+
J3RmKzxDOLoSssXRyyhvdb+WLDPx23DSoPkYBDRLNTGHl4A2rQ0WY+swBjlzUMfh
tItpxEu9jEc1708HAXbiju8I12rLYFZ5z44bPP/AGusYsw+koOw7uqF3PWKT1bIx
3FyUfzkiCJihmEAO5lrwcLsjtfQvKA3607a255FGq3+dPyFcuyNw8UJE5h/9fdNJ
jw1RsrkRbHR2i0Gl7sRFIRvliMugrpg0cbDVoAQw56QLvz9xX7RpDda7FUEpb7VP
FSGyYzCmcpPWQ0qjvZGzAT9FD1JyCmiLoMUbuawrRgea/uQiqQ2bYGIozNTFmTyF
0BNFjcfghXa7CgE0geNE7rc8R7d/jneUobtN/96O7xKBVUinP2Lc+webDu1PXzdl
Ljzw56DWjpFh6sl3k6pUCnqhmB79gNG1kRH2aDf7LGO2JeBZRZqVMT07SqUfz/3e
94lL0z0fStsF+M1KqzQakGJ5A88hS+lzb/gl8Bn2HYnt3URcAz11qVkZY7I169Sf
A58DwittumnMFdQJSTEoS3I7DRR2jmd/bHM19bSnLiDA6SHPjwva7eCEgvBe3opA
4wBVk2NNvj31v5jwYq+spo3UqkiMnCku13RIBvKy1q4anKnJFoiFu7mIoOeEj6Ng
diV2RD1MJly7D+Bvvk6phx8lZu91DoHk3VIEkyfcGK7A8ogtsBPi89nvaO6eTCLV
p4GgChYUUOnF7VxRTenVMuPc1TehK/TPhgCDFTiyDWgnlqQjR4FEeDPMYE22OYtR
SiQxvosEfZddCLrHHDP35joEo44aUN+Qu+3yYtZ2RxqJ6MbcWJVkTj9z3xZzZtQ1
nAxW1Sd0LcOX9pNwbbhvlFX92TiB3S9iSnuz0umbMq5OvQivqQgsdnCVGzDe+w5B
IK5DeYlKgVd78ggod1/FElBHlotI9gzcUABowCFF/uCCsCoc2VL1IT2jv8/ME3g6
yKCsSOY9Xg7BZVec9iU/3A2SCZe1xhjv9tJneRUnv9Rg4BkhX+7zpGUIc1oI1eNl
cOKqononE+DhZ/A8f/JqmFA7Aj4HDKcN95kxR+kdnkWxlk7rcuijb6GX2L1bvo3l
7QktA6L4UCflBeszX0KLCbjJvBGdCNqLDwgZpp5BJB5nsWurOM5wW8EyBNIj4DYH
mo+pZDGdC+VH1yUQL8iLkTZFh20BtSKOoYYMlQ7Fg2Q4HppzNRCz38rg5kBzNFNi
IGe+nhmcQdENi4EjKzP3MuRpgWE3gaygP3LhGIsoBjS0Fev2FFsCkGiQYm2X43++
YIXGInw62ga9+xBsNZxIN9yqjJ/aIabywImdRBZ2gTbHWB/HVBhzAMbTeFf0j/aG
1x6bF3wTm5tRBXJvVNU5hMtsiIEfIWCX0giANdW2geVcN3Mb7iOoVHgPIbyJHH4/
PAkpjrZ0Ev8ZEslO1ptC4SJTnXzSGT1IzNfyc5ZHZrcksPLqxspButRm44iIw3ij
hYTdUwdi4mGm/2L+LaR8YAGmty3kMt63w+8qMOIAN7X8BqvsK15nE6xUKhhlqec7
ig82QTYOTNgrnEwt+Xo7HuWP41pvnjOBu43RRFCe8wQG2LdFuOBnLbk2Y/L/HEgh
yHpIwn8ajCq5ELt3HXY7ZLB9XQ6BHCqt17rLB+UiOfYuN57y+WG6CRA21nTGX9HH
Iyl7SRNS8+jKEP9RYf3zrWhIVMR4g9pnuyCeYLw0y82ODtZB5+L/GJichUtsWq78
56ouoq+21EYVuEzy8VdkgObpu3Jijn3qhaoi6xQIc1XLLTpBxjBIs7vYITOqkLjX
InjnIUwVkdhoQpYPNGH4/PEDanTvJX+rZJ3SYFaP3RnetU3x0XTBU2aQHb/VZyx4
+4MRmKMG7WX6r4ttFbTjnGCYWtQpWVcvh+0zU9Pp/YaKe3umVn4kQBdrArAzuNth
bxAkutO5lF9AVOdXWu2uVFmyWmoRYz/qT1knuJzb1Ed6lQ3x2fUEQxeLRbDGUyA4
p4nIPEH4mMaPGSM85tQavnh/1ny5YXsAiYixm+keR1o3E4gUcmPsfXD1A+iXJOFZ
SQhTROUTJKsjG7HLfk8IJcN2ITTh5OLfm1mwKVHr1cQ5hpMSBJD40bs+ZVkiFvw5
2EeL2ZtvmbAXJgqxCKvvb7PqhGH86YRC3ohXgHWh+TNIHloGjSNaTMweXx+Qq/sm
Gh0PEVjrCxh/alWkP3TAN7gC/224X7UVVZKe4bObYET7GmFy+sFrcO6lIsGS6+aD
Hw8mpPi78fRISmNjocilN/rBDwBk/PHRWtjzCSBDi3q4X11mZcYKqbP4p3Ba7bi3
ZETrqsAMYgdNNW+XUOKB0Z9jXja0IkoFfm0nOVAHp9w90ihQxGYsU2WzlJJxbRr1
N14Cc9HvE+ooR6uaSSNdoP20A300Gjzlmd1WMj507Ko/IP6ZxjawuFOtMhz+xrhd
m9kEpJOYeYVY1q2pUuQzKYYmPflGTP+oaXtalteJo7L4v+WfyWoU2zydrWpXQxGL
wn2uJTZf+hPMb68FQq6mDm2JRkjzRqanSIAkUMvkJZGP5cW0Rk2QeBNV9w850Yq6
HqGPpVg9aHW0cicfT8V9Za6hZ1cOF7GFAE15Ab8T+svH/BpxAaUzkmit7tn3TrBK
n5MBqNFOeWVw2C3gXxfzYLCjCh9uP0AiWkzgoMHT9umQgiTOUmzcpUoCAT0VuemF
PrI1SlfZrb3MYJrHHm0WFAx+MAnkV2zwaRu9gqQ4FPEjCF0DKgHvW/RXcB79+ACn
uZkkxbzAhdrYwyptwJ94UccOCZZgk7dyaKkOpbV2WxBUH9cdaRXSg7Pcqar0Q00U
R4w+6l4TN7OghCsk92hEDf0TApq15yYTv/iLu8CXsAYAkU9EK8A6k4wwjQfF+1TC
qHJxkPSdmtVvFJKH5sRouBz3NuTZ1g/JvwZ7Zia2VXjhvNHPFcvghz1BajnE2dY7
KJ80JqhQdS8220MV9Jl0iMgK4TeG3i4KTurm+48y8yPDflF3RFy25rYE7pJh9ieK
tRuR10s6hvXEFnaFzfDchCUiHrttLkjweqCoCSePTCMvfFMwjjprnHhKE72yTto6
3uXpD3TYVXSL12yheDF/kM6jHub9Rj+wczpvZu+bIbd9FcuRZDYFjDOSRrfXdBoR
fr6FQCFHe4J2Ll9dF2U4Bie7cWlGRAbZNT3DhAXarLsh5fIFu2OGlkjVrQ50/3jU
REVhRno9edD2Z3GS/mxl31dlaPwUs9kxwL7px2VCWWAb8a+AUszB64M4l4GnbB7H
v/2+D6qYN+vecQCAQUNkcK7Nd9eNPdN6GLZfNpsdOclSuS1XRloUznBTjWFoiYDc
H4eCWNbrOFTQHvn5Xg4H4q1jDtkm9+PINaJA5HNPuEO8XQ3Wox+nSfWe9H+9AGDa
cIV7UZosqKjMOFoaGiPJp9cpx4adIRGxn7wPi9CRckMEtauwrb/hL+EqYkhEDnu6
dFIv3/irYvvPpHq3d3nTGiEJECSlgSveDRcWGfwppyq3k0M6WiJf/bQNpwoWovag
L27iwYV2uic+hDx/zD+5AcxKoJW/HqI1OkVPsBo7Km4ZBlInWNowD7lE6MwMkPBN
bzIYSnMCIhPg8oRG2wOJ/wvDg1EkqqJYf4twrasFqMclRcjWmfn+Ct4SBam1cWuy
RsV2oU7EU741K6kk8utsgbwNbCPdq2MEh0w0gjpABOFo7RKGI9BUypR4w0c7Kp2f
J7eEqZqVdkP/fEBotJWhPp54HsZIKqSmvyAB2ICsxtTfUPKpqi/5XhAkkP45LugO
gs6jZ6nMhX1+uvRxR03sM5yQlkvOpkjtkf2n/oYMxMfn6+jdIG/Q1E4KZKnOav2Q
oIIR3ePkYIDjyCF7JdY3mAESUSzRNZ6fj2N+sIecIzvFMUWcxIPLC19EkdGo3EbJ
w00cmCogsC9RnKNaGjyDQb5OAQq7DgDGs5RvEMlhPUP9aeiR/HBM0grBF7M0s8A0
Jiq9IgO4duLR0MN2WmNdaQPqNwakcO9ZxX6RV1k4Pz3H+zmg4Q2lkQ8tI3nFTjUx
E42+TtnaPjEfKHSABQv0xFajK1c758GtROTPGenxNNuNWe4cLptH0Fguy0Q8N4JD
R0DekwXi1F4HjUWWMUdxijX4bXEnwqnjVR0xh2SttILsEJ6ysGN1NLkv/rzG4KHg
LX/S4kL6Zgv0XN+65lJYNuklo6RY0n9uVhhGJuPYabidEz1B9kyiofhRSd78oKZi
+RQaxtA+Amr2T4OeHmxztF64NImMfremUUH6P04hCN9oxRmwHcAKSTLzTEXflYWb
SxBz8Db5G2IiVJ2H+4SkIhgjz7kpB+9o2iLU7+6iAle9ZJAPT1pCL0kgZbu1hoQz
+fPHTEGunnCF6rAai+p51f2ZDumdOnkJqM2IjDouUJv6K0FC6Tvm3/sPnUiyqhDT
jG7ArJRb0FW4zZqJsqv8lxPRujZpM4EV4qFdfbeb+2Y0mp+/AOzupxAscVRrPE1e
Grj4FuTBgQwtvZeeea70cylkG0nrh3cLZRshpXg7wKVZwWAK8MuMkOD+edJRhXIM
ZKS3ucPM1LkaWJkk65MCHPe+F/uqDqQUwXDtXk+7tWP1wqlVa5Vp1SG1hPUsptVz
Ew8ZeLE7YoCs+ICBE1BaXdQXTzFIWYXzduzkeyAyyBsF7RxohfEl96TXdujOT7dC
rRlu4PQC0Um/4rtgXSSfbkhhIZmSHxG96UBfsfnT0jHG0DAbeu7uIRVTZZQjsCTF
BCfPyCye+t3Vy9uLMxbM8guvXn0VgYPkMFDGXtEG7hnWHaqiyVY+DH6PtxM0XT+8
7ZOAff5dgAztfMzkfSSkIY/07fhrWsapZVl+Bfb9lJ6IkmXDWiZHhozZkmFuTgQu
jVBbVpsJNmVHjY18n/2ms8ww3Xb4Wif+ijWMoUsRPqIc7aR8OHOc2iyAfBXXXxKV
nRJtSGjcJV3zoh8e4PTqU37C25k4vciCBAXq7hMkQ5QuPSU5B48UtR3jXAmswMYL
GvMgDwi7WkUz3RuFo/R/HcV3cKDpVyHeAhIrURB3PsjMePtlCKRNyycEy/IyGtrL
seD+opwRrqwbNW9d9ggjnK2NdJzgcbjq+wqQC6K/5gGjIoHl1k1jotSsG2rPxj/l
3SBJ5aX/Nf4Y7Nirtvt84ChG1qIqed4wFyiPZdnMnWQBFfSWGx2pAgbcHMf7qtGT
wBTVBOxi5epp50A2hLBIWsacdjRQya9aI2Iom1XtQ9bsaPE0m/s0MHkOOUenYuF9
ZWHS+BugV5s10OSscN106C4SzcyxSHt9PtNYzSsIobgUTqbjci7IQ/Od8pBkUKBL
trFeqTase/kJym0LbymWWS56wemOCgpRZHomxKdXTQ42GYJlV8rbOZkHvCI35i9m
sPm+F6OyYCBb+B9/JGvDL1OgAiVlOzvy0wf8mOsi1lFNWvB26HhKAaAfGVukb1BX
iFuWt45TORGL22YPEI+56JGFUVg836Ls9JMDM09OMBgjd5xVOM5mLIKALkDKH+Gx
2IVKzrB0GbALdNY+SwBnv4CA7zFusVkSKWCxTel9uc4xmPubpU2CTZ6lb3cAOL/2
jFdqoYMu/0Ph+7aKCTad0AT1iTXB26OaaJ0UaLLmf7WnoVTl+665Gqf7VkWTcE8V
tjr29jPaz6AAMiMs2uW/AScBhGi5BjWbSr8+jTtJS/8Xi7bm1FrCSAIycYVepv3f
APIrMvrkAbcz/Mufvk7Ke3Zfrzq3Wwok8ZsbaLmQxdQ0GOPIr6BuYrjuQ15ty4S/
URJhsmJ9DAYEF+fvYu8mmZptt/jKVfTldBG8KuhTwtdU1C9V2tniBEuJcHsdU99m
l4Qu7f1mTMdJhw5LWS3VdoV3kskdiyvgR7qMcuT5UPVvnaZwFjNxSOS+uGBHPSBL
3zBlb1DYK/xnEPhMBn5QcAggbJJYW8lv9+OFt9/5Lcrq052fP+vNMYxkqrlxcmSt
XLuX+RDVcVbZ+aFtduDruAg/CU/Ft0XKtxm4ZZxEW3WUA9l7dGXbWme1AbZtfgOh
3OzcdzlFj5S5BiMW6qFSEpNhFvWHbeGcFSW6Ra3DgJ8cTzyY2f9tMqrxuImdb66i
zkt+UEH23ggvxBpsIRtcA7MjKDi5nXz4a9AF4XFRHJ/Nscv2gW4oka/eBuFzRNe1
AvMh0ghSMUubS8fvOGb98Kt80T3Uxhg7R3iXKQsJfk2qj4KvhkGRCKAuVkw7PnAG
TpImZGN+ed2AxC8jlSqqCjtfU00Zcpeoq5r3DTT20SwqAfvGI222BSa/wsLwvRy5
nvPcxbEU+Po4Cbm74j116Rlxo/UmbPab7Reiu4sFP+UnQdwHu1+y9ncxRVRwq2ON
xFRXFX/QBnBxZM/ed9rNfOcTezS7cJqNCGxe/7/xqD0FVIRYqk+/Yvg3TD9DO5vC
7wRSBWYZj6u2XsRIMW5XHRpnbDEMONKYb4oVPap4Ceh/Gs2qFopyAzpHfBkQbi1z
LmKl8jI2/eItDqpxOvIN1LYeUcUI/X9cThThYHsawjeam+YWz9JyoCrVmzHVnF3A
GgdEAMMFwd68zaeOL/vTdeOkLHsZS5pRVGVoJIhj3+TWBYMIqn2xMFdHuUh+SRJ5
nj0nLdItMEBC+iE12CQXx/qpAoAWjSZBppbk4FQcNox8WMtG9wqDAQfnW1CervgG
WvsN/wrVQV+OL64zD79mb/S4gdB3b26YKE2+ZkL+Dcbqg6/atuilkc6SLq+vCGcy
ZooayjCyyK3iALZ4/rCFbB1RQrXSoVfxAmciap8SBPmbvevwJsmnsG/jN7lHUUbA
eI16joFvtKXW+Ao7ViG46/q6wG/sx9PScb3Oa+ZefYyryEHF4EzLRLP7LyVmaPEe
j0l45OKYgEq80sCx8jLc5+zSqzNHqJ+sytRwUdfeeY61xQC9HqguaMhdgbUeg+nX
nAn71LxN21+RwQnX3BEkbbsEqp31lpK8HJspJvYRRMDlpY/c1nU4pnyNWQaco+WT
hgJFdeJLUoylQkp06Lm5n7+8mZ+DnRSB4y5LJFGXisFyzv5oukFB3kLAPRXCCGp6
MMCRxN4jJu+wiA/3FIIdoN2byU7Ktuz3ZTMD0bwBunOWqiCzxbR4ornrNTQcJesq
QJe6KyC8uSM0G1aJDXfBifu14no5VprwMWfwn7acEjLw4pdIjacnHbGf79U82Jyb
FTJBFUC0VcyQqwvUTrklXxl1YBtJmYb5M+bq3p+WKpNy0GLDUgqiQY0FJcdzo8s6
dCc8Br5wWs8ST1rNd0W1A4OWCBxBHMOIaKJgweeH/m6IrfAiMneZLhoXW9jESBEu
I89asyBt6G4yCi9V0ZwtoA1C7YqiDZhUiZuFwd/fHffEqJKGhOnRSJix79SsOOS/
ThFHpCdge2yV/J4y6T9UvHWPAEFXFF755R6nfuWA38f4HMDl2c4P5e4xyLxYZckl
IqaVMdnK2Ll4gJJWo4OppmObiKM74SSvaz9bPEPlMe0Ms0nHBnrvOHt91dyqoxmG
HG2s/qmcdSMwLFsFlVPnxQINj16JSS+qqiA1bSuCJNveaZ2G6EZaoLZMHJrqITPz
dUDSkM+Mp8jnJOOXQcXrJnorCpcWWJc7hgD1qw+09CC1IcFC0d/DfHbBGgaD/8q1
XSEGZY60brHin0dXI6CXrCM959wasggCGDL1eqhx4D6EZAShIPcFUpNGoatj+lKT
M8JaolcZLK8m/j5JZS8cb83qogmvDx58VHY7axCnnfYOZYCrm37jYs9lq8HhvI/o
mdk6gnkw5MtU8ErmjSTfCQG+RkTmZhh6sHrjwijwgWHX4vQolbn5bVJvfSYuK/x+
TdGBrgMXXd+SwGtibJGpIvf3bu9bzkt7fb1fki2q+V+6aoyng5S0o+g5v58GOlgl
jQENtQDk1gcUB62Fvje5Su+l/8v0ugEdA5879JKASR/jgYB5p7ecyCkEjRESU7FC
TtaZ39pxcLbNMXx2ecgBxCVdJzw6zx+lOC+8Uw1soNSkDKT3QvO7l4uBEUfl47Ae
2WMAwDJTwrcNnLWdNQm2SHgnYk17ifeGm0yx6JTKmTnydgXDgpsWQsGRPOxKWMS8
C2tbBEYnYn2Toqqvxnq7DZvNxEsRZ/dHadQ+vYmq9lFt8M/uDuLjZN15+BSP+Rvk
Y0BXGikbRsbTsSBzQUPZHxcEOREuRu1Z8ELKkM9piCVYYqjucuWdfRrNuPqvRA4e
n/VkfRCgOD4/35j3cHFzON+mDGjN+DqwSnVKOWjHu8UFyHPUpYKTDgvQarmTJb8x
n9Aah3anGwN5y1p8ghiaeF3N1zyRG6gpUQtQvdjSadJDRKPebYStJoUM27eiOv5U
dMSCvz/85KJ1FT4i85isOxeZ+TeJCfBMIr3Arg7pXMP+8T85DGe7sdi3TwmK81QD
FPV0EehTYDsI5o5plrV/lnkRa+QHaNPGBoOzeZmIc5zWQMGtNsj4QZDmBBwXVxqd
gTF6Q7K+u5hPRB9KoVf0D3huHH8DEErlYwiVf94+96GZc2Qh0RxgkGFrLRn8n+hy
00VpiZ+f8N6jWT7J5ALqtpsTguKiihdjhNNsotg9sHEkr5my5fIwynlg9BGmQn1l
MlLOYZ2rbaUJCKqpKMD5z1NRG+W/BRtsbqcWjdbZd3shzudxWxabKN80Su80ycBo
QwJkjPywwZZz8sXGMceRl8JOWN4Jtymw4e3dDOmQwxeFbEtbUQSfJ0fSFGPmx2tl
qFSx9ahCfYjQMupa8SOi72exAZ6ploIT4CJhcd3rxYX3KE5Nc1RgznfT1aIHT06P
LalpcC++l1qdwcAd6HxdPMaYZpv2WtGlZvLJoalcJ/UciMY8QaYrJ7pCQYxAzL01
X4Sh2eLDwVibNBbKWyXVQ8ZeFZEsCTBcpBKRLeZG46rMvUWdPmaqJ3RYT2tMr+cv
LWHppvubhOgiWVyInlLjZxkMjl377y89t6TRaLCCt4pEW2n1z05/+5VC7+Rc9f1W
+0R6sJTSP/4oeNCMRvR52+LbtCWuqQCKIv/qcDf6CRb+E3HquoNlCkV8PyuOBX0e
VzUKqBAbrktkvOWjzUUWtvsUcO0alTObdjpp7s8TmjY2emisIitIvc3gNva1FOEH
yDZVi0gq6GHTQ2z/jVf10JdEWMsU29kcz0ON1p7Ku7apcU3kENblDvmwIQWbHEWR
gP5frIIIWtz2b+Ac6LR4L3xG57eLPVeEGfgZVQbGqgnNk2Y2ZmuzrcA7TJe0OCyk
5yM0y1hIAIcddMrVaXr/RedahrRgKjDrMN3IPZDRKiPWcgn2FygMiQDGIajraA/T
NeLcOdvmm0twosRVL8quk6YxHHFtOP1d1gYTsu+p314r7hva3rob5DAOX7E9B54s
ualBnmsoNGfG6ri3AwOhEVEmtTinL1411Hh9Rgemfgi1CLeuciDa79RKNQujpU4I
IDsxeyqrHXEWpGYQrqIUTLWOQ0cE2ivgPKzIaZx/tWqCdSB3r75A5KALdxTfeSIv
gk5Vn2Z8ve5lef93rlYxKR+AxyqkHlKDe+99m/Febn3v39hZQL8YkZGTFAnaKqKY
/tiFSViBbks0kG2+u/0fPxx/MlbG/Dz1/7iuDHK01o6OAdCdBkqkLNHGPBDm521a
7BUg/0buaYK6zhCCP2DG6DgJU6zzgOwDnhuYqf9K43NQ0EfAJaMkyWfu6vaLrwVZ
TKsnbWHckHHgAr+HusOZLvqBvaOUdDZ6EIoobFPC5N9hp3z6Z07M4HJnHJgvkCt5
o1cIWNtyu1iqEDqEZ7ixvS/ZFbzXYILxzman0rEEH2TNrZbW9fDra0KY8cEpRRdD
xAnkEsmuelFMmtNy5NTy8wSPX7rZXh1mPFnyj/+9EV/heiaCIzYEchLV3NG6gkFL
z+hFiQ37llFwtChmR0sJxWQoOUaJXLfzCEnKB+7VgSTyJzwWut6pnDQsMdOug17n
ySNL4g+1k+ST+N9bmw1VFGPVXh3U7//5knra+QtSBrR5u6ta+439Cj4Hl5Evd2Gn
XWCna4GKR136jILEH9IDrKF3yxHfzEmSYsNqQV1pkR3iFyu1GIaqRp39cFPebj7t
XYAuyu5C0bAeFNhUbH8zyZxHy04jECzhL21KO0vrdX0DjJfOp9iAjmCdLdC5q63n
+tekN2wP7X5AZ4SII7LJQ3Sq3sBC9zBr3Br7fLT+OfmtPTAZ2e/bmCn6EZk+EmUz
94XGHKAF2PeRwLkeKAN4I+nLFvMAObyyJqIGlmYGApcMZNIhOyL493yZ1MpxcHAQ
Vlo2ayZyT/T+nYWvAlI/I7oiNcPclprxpCYoNfvsAI7vT+uNn5hp2H4CW25jToN2
/CaXwW63g2GGDJWPnPylvxn3ITJMK9myYPC/X1QAJkNmJDgj8x3Xg7d+fTzh8tMy
t+CIhFb8qwbWFu9Te/mL9h9AnwXrVUZ6aOgfyGtuMgzemsszmHx1sHny+RkRcwxt
9K2CFEAKzGtNBVLa3Q5uY0eILR34LVc6hbXmGWKx3lzaIICxoLSQXDiv7dXFdp2V
4S9iGKcmdgnCYvxkfeooukx/t8Rb/h7Qj02FMSxv7eiCaUtXSD7o4dYwxbd0AiCS
MldYLdx4tiA4Ymw3BZm5ZvhkMIl+Qa9r7lQ7fhcyxus3ypir7OsxDNUJ6onm359u
LVD17u3bUwsggBt9bk2KCD31yqDgFDLuzVW/sahaQnhYnNBci17ziXSmnwtNSWSg
uh0/bBAOC5pUns1gSUyTbHc0m10Bdi/8POCFB5HVEiEe3vPIElcUZ/2YPXPsJx2A
cDt4KBGq8gQbpe57/Tp5IqKvI1pu+sXo/+OMxid+MJgsC66WI/6xLbHWsUX011CI
/g42XvJEPCLiHd0CBG8bSMqQzJgrIonMjr6coAfhliMfFjA59VXuvnglcJBL73E1
NhCNVXmTw/vinnWRSAsRLA+mOyd8iKOLSKfX787vPNyWAVq968HxPHGWjQ4bBAiv
aS0OV2zrHwcLHEaEtE6OK5HT7bxz0FgjEFY5zb71AEkKvKtZ1iPiio2owsfd4EHv
hYfjOs+YaZRI28Xoq54dzK6WeKVgtju/8qOLCxcKPZCo16Fjjuh8lJu/ER/kVYJk
VA7n1KbWOUrVi4U+B2uuY+EXrC2t8VZCWmOyVVaGurHIdoWEkFEb4qm8ea6jRvAv
/L7/6ehKATptYE+xFn0tnz4JBQT+7oHXWyoO0PIe1I5NY58x3lOFdI9oG63QUJRI
K1niAOS0OPsJHaz3Nv2Rjqs6lvOWSw1EjTfaULnnUdgC93flltZyiuexzl5POtjO
83GyGJwpgESCuqUXklnQg7Tvt/2Xqs9/C1tLRU0levCQul8jTUVy+04aLiDGXpRL
KTgT01Zlre5/FAvu/XV3ExGOU/LN+bgU8Idgr0TQPXCeSWT2jaiPHJqAjVR7u711
qiWQAcXO6IHSTXJWowSLDgF98Vk2o8dXiV+tY0/9VaWjLrsuJHc9QiA+D+ZULI+i
SzH5G/OlaN/lenvGoye0a9GwDz3IVkxbEDyZ0PYalSSo7IRjBEsBK6QJLq/6SrDy
iC4Oqj2lEik2t+CMWzmp9fMHGh0h1ILsUmHY8Gj+c70Ic4mh0WkUQvBeJ1caz2Gm
GSMsHsC1c/or/Jy3kHEwnm4qwFiPP0hdD4lxKJgtRqHB305+BEyo0SPFGra6lK9l
cXOjAHeW/mqMC6uLsV6wZY1T/WuovnvjdMiDI0wzWIiQOTGm/DyyRnadiAg+tTni
nA9TxkLVXBDr98FLIr9V1d6sBS+C0ZfwFowfrqRmt8Vt99hCUKehF8ewvPa1KJEl
pLxbyg11dcsrvdQHygt5Pi0vci88mcB7+mC5hIJpXemCubUvX1UYvEgEtRlNJG/y
wtet1PT7WE1dSlVnPBdA2qRwCROaMB+bXYVKzqrf0SHEzxuY0COcSWc9xhu1SAz+
KuM5ZIShC2A2Rt8Jmi9lbz0JUXonVsOma2ppTgCgBujMUMI1obWsBraxrbsEbpSt
nTvOZkzt9CfND2LRa8WF9X5HVBXuFgNs20E0/ilE06KGHSGDByx5Rg4gI/4PSJH0
cRO0gBhkt6tkFHTLm3gWkbgTXRJFyyaljlgjA4yQPMZOVxIQU1/BabIUfRmhIpAA
MhclODoAq6Mv4uRzPePWPXemA9bWXyZM+lbQnx2cHoL2LTRV5Oged4GgOtUlLMhU
uOFcgKhSDE5AxpZXo2nLYKT75nGDVffAJvYdNGd3I8FlhuDMX7NV0ATtWPQZ0odu
1nFrLKaBAaCL6JZD0HXQacXrWzXStphGWy3UHBLovVhJF+TUWeP5xdXw0tnXvzHN
912VpSLJY/K+15hxIQxTMxtKEXkzwdAgrnmwsK9kQuYJYUzVVXNIT8+fE/rgaH1o
Nv8fcHO8JTs2s0nwFqcWbMf3KrsGofidOxGYQgrJ9/2BTvpk6YwtpdnM1hZdrRvU
vpNPCsjoAwa6QQvlBclw5BvekqoKAtY+EHqEo/XP5EPylst7F0y70E/Qi45j9/Fl
pF78EFdYjTJSi+yTtl/ugV4WZRtv6qSZ/yZ7SFEILKsI/UOwyidYxp8o+zEjB7Wz
f2JbV5+8AeD7yOf7jRkkamEw82QdJ0qe6OmAzi5MfNLWcP6MYVs/J9Mf32R1xQQD
thr0rFgFGrekPfXSJePR2bl1J2O/fnZYMPGKVjrqHDlFUll5u/wXy1MxMTSdcEq/
JmnbmlBSQNFgdhjXf4X5/zsTPXPBe9y2HAEejAm75uQMg5wgsXb5jMvvtPDpKz99
ZOp5j6lW5biZwLTYOodEYlLBDQyLL24nkqN9IwfMFhhDGYeLEfgANKL9n94cd7Ot
nitCBRf3t3fm3/OnilCwudsz/ZG4n03hfYQH3/65kOrbxZMmlwRbggH9CeAq7GTS
8NypJeosISzJCcbUnNEngr1TuGN9SKNFMoCjl2JlErZCBrzSbtlGpJQE4niobNPV
kUPo1bf8tqdfVvUAM2syBqsJT/iGKfiOptlwzbMPj+9LI4y1rnr3Vhj1xuHzGdiT
nV31zQmy2fsKC8kwlMKeAGmS6KFMZXq7YNUS93d2jcWMfm0Pw4SJkZby9jPXsngD
0V4OyzeWMlQY9c9L0cZ3wSs3e+jQ9Rltf1uoG/fEFsKk6eppUSIzeQKCYklqAjJw
PGHjE2nN6gvnIvDEtX085cngnbTnE8BqKcxL+2pD8iE1+DdNBoxXk0Yf5mdJiFmY
a9EoF+lAFc6y80b3mRZhJAYFMTRofDOspAi6v4kn/tQ9YSnA+8PCIzC9i+3fTmdO
bQw4Gt3ggIrLVHndNtKWuQnD2hhQe56dAiDxTLWXRUGaPbWhDBvsM846pgyOAB1R
N4KBFsiWE2yrOGavPPLfwjdgzhMNf2iNy8PMPZ7InMIu7TYUClaR/86liz/3O5ux
EHPnvzz2EHqKIsYJpjlu6xCSNuNVgpVmYvGMecJ47Bm3K0QiBToBHZoKj4eL4tqV
X3RmaeinbngN/gyYGKOwUzDIJEc6EUF0nvCFi3sFdFBF8OL3XDa6ppJkouF27vTy
+em3yh3PfAvV8JmyVVpVFTwrs6nWxccWplsVhT4wfu33dsiKV4gCNU3fAW3HwbPF
khoZkTcs0jxGc0BhzYizTKH9BhlWyl+nBpByfYiasZFtEiLhA/6xSVi1j9UdT3Cm
fvY42B4CqM1XwZi7lXDyDhGw2noIOO6K0+JQorKbG55vGKI51e5JqVDi3CaPDlLN
QKZXI4zlxaI+xkRO+9f1nPDP1KVpijZ34qKGdxXoBYlH8rki2BA/Ona4vhy7F1qX
1g9dbFR6WhcJK1ZBDhSNDyTrGdvNc2t6T2gvLtFClxHAknwpBq5La1STftA4V21b
W5H4RANySkWEjOJbw/3ivZvpuDcuXISkX6kWgWkiW9mRm8QK8GAYTjhZ5QrxlGoa
omXjNrYGVLCJwxLswmC7CzkS0Ks2mKNhnA7FKWx9YnnqeL0HbX42hBPV0xAHV2XV
GXDTzt4PfhhEunCHZDrTcbB65yT/AtlWW93lYA/PRI8R+WVfS1oD22mP3LjQoFUn
dhsPLG8Fbyhyof1MurPisbunTvHHDw6FBcn9pBlvjeRSDuyhjk9SwT2nfGDLVx6F
2ws80jfeiJgQHBE8wfqBqjWR3/rSUmmZkmLpy200bXVtbZ6Z9Fx0gRFIodzB8Jej
hHftKQM6LoJ+GwI5mHWJxPQdNG4ZVpX5ABW5TuydpLQrNp58dXZAQgGzDEF4BESI
43L7S9sBzZm+QuWOo4lMOJxHIziO+MXShTXRFwqOh5/2xrUOm2Sypr0C6i1qizG8
qbaWsVuhBVGZcXmXTgJfIE5dRZqqWY9ans4InPw5f17MuCtyNVutiVwGR9Zpcemd
q3Ajv2qQQ4OwM6cYGu31IexB1VE+DdAAu20FPPoZ4mmvuIJ175or1J/9d8ZCj59o
bcsScF+eaB84PsITol306DDtYLYov16FXYFdvVHvRv/8bUIkQnZ/7Cejl/uWGSXQ
tQ7t5hdVpZPA/NTNobXWHRr2VmOQ66E9v5mJAkwEOnCGuudr9gQxpNST2n1zgdSq
jGnh5XazbYVuaBIh36Qe1ooGzoIJAVdTwTfgZzSJ0FchO7U4tEkBfHsj1jOivz4/
3Huvz1O3ktFd27oxmp4f+kWslpBlX7Pq3/tj9z7ll9nzz39U9JUatE+9aeZHtOft
GrCpmFti4DdwHEPN7mJd+Jbbsp7Ff3ZFqlot5rOe8eeqjx0AOu/fXMu+4M2+UDjF
55/4GhiELoW+OH2A7A6MHCxlGNXWcWl50ZaUD9nsg3ttDWbeXBdm+vZ+sk6RCuz6
Pxe/C1cEIePXwbJWc0R4Y5cF5FaxrvtyikDIImzsp2PF0tpIzIpHPI2m5/5g1D87
CVwAXb9mv1y+Y8SISW8JxnwUH6SzYtqBllH18qvmxjjTzhZiTCWzUCtLQp1I3Htz
GrWdN5uJQr1FQp/O5Clf/arrlWQxCfq2QZJG7vdNc7ZMZPfjuyFF4Hpf8SnAy/Hh
pKNqJMsoWweuwxXamlWh8PNn0Ql1Ria8ZOkucXn30SyG/HcG0ZEbuXapc0k+usk4
oUWk34l8WHnL7MqocGqospXSk8mP4U5MxDAu7rzs89sjolIibc47+ti8o4PI9HXC
JE4Q2xGh6BpulaA/R42NrkMVpWgZBvKUtooEcvtgepfnJz9cFSc/dDuCL2+B0SUv
cyMDC2J0I3c6q+7eyeGR0aeRFZq6QmmPg76SCmfWreNcyUcx8ExrRQpTUE8+dxZm
1aC/RVqTPYDWlfDn2lwSlfWItr3Jgu8SriBOl/9znbnu5f9TU0tQm8DO7spkC5Sj
uZbG7+Ait+K9UKhCB4PZi1BgLc0cupnXKcuJA0BcboQNp0rAZayKXeXSFLLy5A3y
k/3OFaatcA/zbon0qnnelgcLMljoOT05Q4KjGzjAPkfwEQezIcorHts7ypRDO/2A
TLi16F7/bSwuq2fyDXC/XJT+O+7RGq1SfHgxmKsLPc2MoukuOHM8ybRBl9wrt1c/
NYSLLrQZFCywZPNFAsepLNEIorBcKk1TqCppVE1Cq5yOICbcBvfLOyrDnEvdAjI/
YnwAZV4/zk6LocRi0KG6EROHfmV1KjO56Sx4d/df31JfnsWDVPG0iMPcs1Oax8n1
3oWjyMNc9E24GztVvLNfggscorRRNqSb1/4Hj21nBwKMDg5i1ROcW3nuNXStzyjC
pvVJoKPVfwTYpsAKlWst4MqTzujO4zbKs5yMU3clamNNlaNwAdGUjdXeuGBhII/a
pPfl34K668S/NnFycYgkA6b9dF+951IGtdLOIkGq7u3WrcMmygKFY6CMcVHeUlVh
ec431rL5AYKYo7ahOLSGe6ZA/nlxbwBPDlOr+0DXG2CwDtuwcE/2U4a6Q0P2hwYp
tHRURT7Bmj4O1Bye98C5MF7jkZMAiDJHGxNUuJzUJH3EOwnmZQblJ5uOe3NxDYp7
1or0iCb7Spe14qvhOMt7yZSaZqezBOC9RKMLxeloq6bAHTo5K6gzdbLZ4oCoDEMB
UEjs2MSOuvK9JEay/GvEVitP+hK0mlw6kkO3/QUx3+sEiIDIEGKQU+Oe3A7pYxQ+
jGNA//e0/+9GctKDBcMKsna9duHvAvQwsycQNQ/EwiOKDoYt2tMfyWFte8HRinNJ
V4+nhwqhUb/c1T5lZDQtcAFLJpFn9gapwiDN32DX/btsmuu3kFGqI4suSFgiSA0M
upshlP+g3osSm3Qc7Gi914CXW1rKJu+WrSxCuOv9Um/HTehAphUFl9GT+VaBVXHn
+uY5Ie5DzITOcWeHkZ36o2r5o8rxRcjkEobNrJck1ry1tVUh7kAnC/IeKubOP5y0
+EVgnPN2Q4b1lr3ZtYpJF0ckIZOVsiB1VRnBWkzztQK+yUL2+x4Kl66ADCQ0f0Su
jPg6w0GrIeSz5BH/xNVGlgDLiTCaqTEMh8hdtrc5dHPJn7OXcgsLiWKVHy+uJb5y
NJTSfXKD79LSc5wnSVExeveICDa/oXWKSh93Z1BNVm04JUbMVa1f7XU9l+swn0hA
hxoozSABAkxwi+JZE1iZ9WEBfJe6owVICMNPeAYAxx8+lRfmk+7hGBXNfkwyTMmx
gBV82QIhAdaWDQ1bdaGFEwPhTB/Y0s874Xioum1Si+f7vI/1zNGOXOIaJIo34wZP
r4ko47c1GwfENP3vNDoppcXSXI1h2YW/i+HIWwEncv75YO4XqX9ErAxEMbichx/s
7O/kjoe1NS8hRAfjq69GDdilib/yRlzOB7g4NJvUmcXhjqhSk3blQpFO+5q8sSUa
veZ71Laf698SlkxtbhNH0y8/psYYTnVgSKAgg8Mrt2vKmsF9cBtE1vJ9WMrYbqwc
XXHFFOZ35F/efCgkflUTpilhGd1NmP94IOlOqTn+EEuEwKNIzGl8AnEamZFJ/w9d
wi6tdA8k2VWQrwqoWWOdln0Jv9rFocZGk/sDFmTMOowTvqKGQCrG34+FcAw8yg/R
ypl5eKKzgisD3nrY2vJS41YD0iN5eN3jbecVfU2b5OMWegdswXa9EXsgB6ZEPCl8
4IbaTd0TbQ+dx9WkmgE91PBsBD6nm1bMRbUCGlVZKKvL74eFXa9kcBW1g+MgrMxB
gcm3Mk7EXnpf8L8tL/Ce8a4I2jN5agNq2ZlRbsvVH6Qh/kCj7M40fbPgs/cq86h8
drlwcbfJFNudBEdqKllhTL8Le80CKNYvQ/kIEkoSUPoGhduk9U8gXYxTskfD9mx0
nTN6wiXMnOCEoab9+95X0RvaAWlcceyQvlzXMtcANCXU869nNDlUr4hdI6GG3wO2
HBkLZ90y3afEwL05+x+ducqFvirvAkmX4nYewop1Jdji193SVRYI2Z0NXrJrEKOZ
opwdOUdi32slwo1ElLVkbmWemxN8OhUSl3PR3cBJ0msSlhR4f3cXOkMns/v+TxxA
etE8ol9nrhQnl0ngrlD5k7U5NFTAE02OAAfBRUz97lvpK1XC3nroT4PyU4lMLzbc
lmDYwQGZR1ffomxHQUuUgjiMyxizGXHz1o8oDEV6zFl0iTvt/cXgqozlOOoWTd6v
wT5b6lgoX1/NFeH2Hg9BGsYf2TPObihNh1MQGqLvDlBA5UkIQWzdPK49oOJpf6aM
TRb5CHeaoWZV3U1bcX/bsizmR3QzkaM9OcVHRJ2p4ivUnhr3Csva+Ufy0x2lKPFA
3jK7LpHE1sMS5ievKsNajcoLpjtGoiehpWundd2dQYX9zxf0f5DcQbwE3XrQ7n+c
VUTM5YVrMtV5edR0/CBpwjmfAAPHp6ufTSS2jmehYbulWcgCvcZoike+4NPmd+WH
qidLqvMfTGxZpNUnJ+/v8c1JyXJ5hhARmelaM6QTb4w044oPsGWj5PYJ/ibT2C+4
7WG0Jvff2jp3bhVf1R7AA1XvIfER7rrFqcBO6yR2ECkwOrjtJrWX8w7h5Yov2u7A
/DBuoyXKguTLgNT8UHhC54KBU/wjkIGLUY0a3iSjyyxbeivL8TRRKwW0XrwaRMFN
8HcM+D06TjJgiY+G1/WmU5jmYa13BCbAy7hZ7m+amLAPVsOKT8MdwyylMlYUlEwa
DVo67dwjZeUNK7Bz5C5Ne3fpqha3ZE2fOYszeO0iJL1N4+Nqz6EYo6ocQOksHHQb
eI0UYydQSx5Ja5jEbCijQR2OpTYjfQhuz285/U21HOejOZbIyASQMAfsc1QGbJgq
kGdQC03G/OsbDdohz8fAa8/w3pZ8fz0cUk6XG93ldm+C8+2R9PIT0y6BziCx4Aqj
nGUaIczLme1ZOtaEa1feNwFX4VnhIvif8AJIOiIl4DxxbtO6WqHJHJqL71qEgbFl
l/ipU1InQ1qfJwZ19PoRzKursgm336OjN/EiQ21zP0J9MMKH5Vi6yJuUz3y7fcS3
Ley2/QxHEX6MJFLVGudTIOXWcpVoMe8G988ca4+hYYkMFbZKXYY6TX4ndcyCXqRc
v4TwGXWsr7bpJcb3YYPihJvoDpCDizEltJCtOXMn12SbL6EG2c6z3INUwZ5HkxwV
asIEX+uxrRotap5y0/Y8I+fLW4BQjKLwJaiFWwjblpVCdaL5BKyiyC+YBisbhQDr
73ycVNoQ+o0TKvEDE4cPc4YUucrzQUt22YpH/zBkdQgG6CACk41Mp5Sr+NCVUJeM
qMM8LtQ1xB5yaYhOkPR181Kndhn5NKtORz9B6ECtM9xiNtNWwDg7zi6WY44/4gTK
zrjYTfFzMe+NSbjtQDUbkDJcpNSZhNJQBB63Ul37RIX8ZLUiMOPk0MClsTHStgz3
vlMuNqnHbaA9kOvRb/eYWbOjSxttV3gimxfykIgH8/XNvjcVVJj1/vAxOxMs+XWK
wRS/tMAStOsj7gLymku693FxsaS7jvP2Gfblsm3SYOvKxoeVQs/xt2Zqns82C9QM
vP+CisCEJkdDU0NkFTuU6zJcqIy9Hbjfk07iQRVdR36WqqEDyxMSaPCCUKHdhuxT
QNliFhx1RWLXu8T4/tdcGr3KWbHEgZ32SSMls6aUsjFbkJ6z4IhqmfwQxyMuwT5n
kXPYIL1xpn5yo7oQVwtJ9Nh1PVwJeIEC/PGyd7wFP4UmDIxUPaKsX8uUEjx6cJBv
qaz6ZXdyK6CqjTWzE8CVgPtGAgvRIqMUuuZC0C6NHt59+3AggtTG485ilwfr4WhO
iSczr+14dRJTYDO73FT5hcXrrAG+X5KRNDqKPDLWS8N+4sWFoEAfc5H7PIvoiE5a
tQo8WK18daQTLaOEelvjBHKMdVcs+jQDEDtKQPjoeOMFPdUuG6VKVcO0NjJezEbP
SR/QYuXk2337Bobsbe6G6qhbrYGrIOO9ZajpKRswbG1IPDRgzPTDXwoQWkKk2a2c
zmVaoo3Z3ySQfQwn63jhQdApMSn53XEN7oOxP7IHnwCG7tSqy8DK5clblQrZHOcQ
d8nL1ugDVkkqQImwy4+8R6bNTrwXGVUqCXjeH9jB72JWMqOFXEv7CkPi9sBr0CN4
ARkE5BgvejGGR+DqX0S9ejwuoE71NGECsX56CC7e0ODFI+zTph/yhcSdr12fW5Tx
1apdq8qwIJ5/L9BxIZxs0UPQAySvVrUFsYpe4/JBC/RNhzdgmNQmvoKFbVbaQuBJ
e+7sa1x4woanvH2avNPBhMP0502cv10W4txvNkQrC2yFmLteZlsv4Ef++7uABzOh
dcNbIDa7SMCeHxnXgUPWsFM5WdUdiv9OuDE1F0QlEwNefpdKDoymL1vUA1qAIy5t
xFfQqtuB+hp2C3YQFiE6FaGHQnUzqomLsaA0XFQtFJ/aFLdAu1qfNGSJKF8c8T/O
S72TuNiiDFGOKX8PtfZOYDkVl8fkDU9E/TG6GQDifZ1PvFCu3WvDmCylvbeFKQq6
iLYI6nmTm6FszespjJT7e9V7yqVhDumD/LwlGwUdF0muVpescDvo2r6rohGuAJUy
KKmhTRCB996WIxjxIgRapBZF0JyE1lr+O90Hn3+WnUPiCZ2K0KQIz35EESfnRrM/
bGf2KltmFy9qTEa5dYd0T+DQS3vMvKrApIdMyLXYx0VXh543csgfrU0ryXOYTXU6
Gq/VBib06FiLLSPbvavk5TeT5ZPc65sb0VrPMzRxEhzwnDYDxOdOaJTSkaIF7YrP
MwoNSnIwscGLAsP0sHH7tyh2bn6rfzm7X9n0A6eTB27KxqkfmHKYbs9qfFvVGBOL
AnrYr1yrNCSavub+rNNfWztBXAFaKV9ciG4HmfLDRLx73niTbOqE9zw5+NKOgxJm
0jhHTu9mPJmAj7UIlxhu9Oo+EMLqVh6DBFowbguUhY2h2cXA1jZLIxaP+m8Kzzi5
13BylLpFesNdgAOA55VAcrJqhBXODDd8Llrlk6OSl+NwtmieJN5uj9hwYV+YYItm
/hYgwVEP+NSrzsZhsid487fT1el+HqmW2JNgKGkhtQgEoaB9F2h9MPgDZFlU5YIB
67bHOcQwrogIf6uzSUqgpus3hKcZEDKUrcctp1lhfXgYa9u2G1epbby1S6k/t/rV
is0tjvNO5UJrmeEfGKhuoTd3/gjcBjQ8lt6hwNE/PXIKiKVBd9HIph5O66vyPy2D
t6ErWe+54opWUoa4HcBVyF8aHUuISNu2gtrma4Js47fUpkEUKMLfVqemd1wF4myc
1fjTI1eE00+L7IGex5uwHTWKimsQlkKjiMk/c42sGFvvXRhZm7eL9XMKUi3VjEAh
7kYiju8R2RhnUD63tcC/fo0+PRGR6rLQ86+bWEWT1RX9DxjE8vfOSKMQFrFCZYdj
eauANAnVFutsAnCe1hCqzkng/P5SPIHlqsTb/Dk3q65E/hHCJlgDN0JTgVaKbYwS
oCvoujD6/J8wHmwSOaNFWarExT9u4aSlIqURhu0b9z29GaaCNjAfCj+vfREbKxNS
MDDnom4pxO0QkfvSzLBByH2U7BHguNd0t1pwFxqdUHt14UBpR9uCow+rsH/rkIVB
a3QAu/BNKin83Du8CUiNv2k8jJqGnWv0hFB/rCgYhaLPOkwPNXrkCgtd9LUQqKdf
O1r86+/a8X6Ha1pTCjPxuesT01aQtVn5q4oDcm1tvSWOun1tCxE286LqOypnWUAY
8I1be0Z0jvXmZOGxFWxF9BpAyI6tDyWqF5t+SZkx+HiVuDrIHuMZnWMnbVXAOWGM
1Ro7G25Rqve4kQojqYK6LleS98fcq1JMYJnwSJBX1/W4cYko+EOsn3z459liLla0
r4UBBFPKcaeptiP+mGnc5K80uPUtekyViy+Y1J3xWP8FxwjEIPUzoDiSL1zV5bRq
CotgIRL7sA//6/rkeJcEreaXADxUVw2329m/atspIar+W9BdyL8FrJiLKx2nhurf
G5tE9QYGknD+Ur2kgL59rwoL9bM+cdoqcIhHH3uOpoCKV+GWRfajbvwMzX//gnmx
ibiXi5aYix/m2VTv9SmuWvH1/TEwWXtyHbsnXnraTvFZIy8N7KHJ0WOdwx+KqsOg
d9JgWCdLi9ze3Q05VKep9pdKtYqR6ykz6u/Ir/0cHnnGAcn1DLVMpem2Fj5yPTci
5neR41Eg6+IttDcOFCoEBbMKBG3w3NQDknSyoZYPZO0fwZ7CDZTI/hN+SNeRfyjp
ZGb+Z+7z+37AYWGMYx0Wxd2gZ/tZUtDQPKOdDSvP1HePlMzqCS6rjuh7OTtoEKkf
S4B71KUHry6li5dFVBY23NKfEqeZjZOkICzuoRCKrZUz+MGmF2CtbxPQwaTs8fUy
oiX8WeG9nzRPcKj/COZtZH1r9aDP+Xsr6z/aIPDeZTMM3eZqcH/S8S1EJPomORIi
N9xImnmjq0Yh73hXrIKKBXT90mvDAYWiOqCCm7jt2SUfJiEfhuNImPZAnFmhW85t
I8S+NY1z8tME9Sm9Ti1F2/oUVeHEZbyVUNYbAPVoWNVVPgz9quBOZeF8DsiTTItF
wSAa9eP599wJxNWaGb/nswRI/1AyYCsbJWzwpRoTboDAMreRQY3YegFQzP2Lv2Wm
qvPbV03bT+PxghKFAzvCxxe6n5owkYI7chcubwz5VYdGwpy2P9vRyd3GX+m7L50H
1/6gS4peptUfcpUBTndkvzeNK52JRxrRL4gTSaef6bQuR7EoTq9lNR7G/3Q9RWso
eSzsivocTEbFJIttOPPwE+43CcVbYeGZga6hchBr9ecljrYMc1wcRBk9zra/63ro
ToJQ6U7Zje3n+hT0pDn4qYVcLYDtlGw5oGDJAeHmHEyHZ5Y/2MsjhCWgRm0aosOn
4NGW1haccsI1o9B8btZ6rh7pRPBXDXuD3N3feJbbuVaEPRJJ91wsVah5gZnTxcL8
1AndkPmTyGn4x238iS/Rhm7lh3Egpyw7nR/1AHlqtUP8w1ZH5IvLqcVNsTgnqKj7
qvT+j/W+PW5PI0Q65Nugo8BDxxjL6oqScTfvtMphGSzNanwT4RkUNgPWSAG0eWIF
HUARn7KQvud3lxN+F7Vb2JQU5fMDwAqjRdD6H/rlZ/qbQk+WPxH+YS84jImPVPFE
FRbgQS9fpNPb8s22LtNIGcKkfVIoErL576Kab9zL8EvQkQtPDGLhbz/y8PUX6lw/
UMszKVeJyXVknCOvcuOFCTJ25KuZeiqA18a153B9PqR/wRztN6Fxk20u6Mt+feEQ
imtxKhsu+XaFpncfcG/dx4/A4JL+wHNi80UO+joSY683q/rwYrwDIaxLZ6BLVY0n
FiOz3cdbl7fakmXnvQFj8c347DM0qnQk8NQwL7VsdvZlHLACB3mSHYzuUicK9Edn
+C6b8Rf0akEfImUGZSis9CgMC358UBxHCvqCtHt2C3DhFhl+iMZ+fomrL63GhG2X
MoXM43Ztd1+fNnu6lgh0lL5OYWp+JXR0YjzaxDSH32aV598uR8Q1k41xSbmOoGv/
0ck+5OFt9KOUsvd6q13AQoJK/oE+e4n+1ecpH3cr/+y6wpCK3qEd+WDy7LKGBj3G
4OYWXF4wOE1JcPR9XXOeoDSKw0xee14YMysDx4q1Otnoit84pYGtTU3Ofsgnl9RN
aUX7tzVJZEoH8v20kgMVR5EraPxRKAykBdLaABeP93ALiNU3CZLvAvyMJeqQqCsK
ykeZtLjBh/RkF9sRPS5miF7pY0ynhEdEyDsU18UIprD36TMVn95B6xrM8s1WlG6K
2t5+m7EhxvdPou+LYjzdySnd22LxJcZ7yE08mHjrLymCKpJgEEt0ZB5sAhDzdbBy
/IPfBVV7XdXFSIwOrHrosAPK1hmVnjMvW0+edTpWEJUviBmAaLRhjtADkfBNp0V2
sWvN/87O1Xxy2ivkSotY4a06idzIrbIHqn8FPphN7+5sHfqA/1R0UlLv0tllxLdb
/ytmIXYWs1VU3vqt4T+C0UAsxmeyPDfywve7w9qnsI7qJxFStiX1MDp8M3W14m1b
+DCoDHYTeMJ/B0kEEfHghB7E9e1m3PBvP9mpHYk2Z/0rzwih/oKLDUT7//Rr4pT7
0+y4t7bVs/+b7q0v9Yum0ryWHZ5GWXU3mv/TqEfM9/Yq/v1H4wExp54bnkZ0JHe8
k5tY3kRJ1/Msj01SfjNBWbwdU7fjOlGWcNXlEDzwgubZMWGyobqCz0diOyBgcaxZ
hfLvunkDozKQqqK2BuWJA2pk7aex3Yg55vK/1pLa22m4BQkt84c+MR5MBNriiPxV
iAxCifoh/bYe3YMayZmuy10F1nhsQghv+pdcXIcLoITXpaeOQOcMfIjpy5bxfI8t
S28gA4GPS9eRHdruja/KpqRIjH9zmBzyVSP6DaeFXsjxTyMwfVL/XWtGghxLIKhi
4o1GBliMB+edxEHvl2VnQevlWMgimXDZquWzyv/ClhlNtS5JvMPVKTfIaae9ZyUC
6rmkG6JDszkyWUUICuwWV0x/y25LD4g2C93kCxzwihhOh1cLJ5cZzkovuOUjWAvB
h4N06u0seDxLbyFhi59zArwVbHk7rmbeTXfS8cFoJmBuaIXYACtcXLSbkDWFMMlf
C2wp6zuw+za+ajkRvErEquflcVGV5S2ap0ym1LI1LB+yVE1E+Ed+e3w1cBkOS8X7
PPa9lisp1FAnBdOx7bt+BbqkoPj168f80mvJYyymJCrDltM75JRY0z/CZrhrIl8f
JjsJg5Ry3XrwDIX7TtHHChNvvvYWTd+im3FV6Fz6ZdJgr/T11eGO+lLbL5Y004aZ
WDGVs0fdgQJy67Y2b2jH+VdUOpqcc2yANQ4gz3bxtmcrojzoGtnMkEgEuIMD7E2b
iDIUSXXzZxWdRGAQGs50pcx/lPjmw7ex6jDUk8cXKWtfbqtCZscVFttWaNhnBrY8
q1jdkMB+p8JdVsZOcsF8ZeatvJTIPfWASE5tklAQkdvKlC0kQia0TkLEuOAEQkLG
vPWwAhn1cO+/f8Cyi45WlVGqLvz/HmUVw4rk83LHC5wA0LV7fyklZJqOeJ4b6nOM
Bc/nqIxwjVU7ZzH1Fh+L3trhdW+qobc6/smWq5SH/sI1IV2TEwHLRqPQRoYcLntv
7n9NUe7gECvRoTj2CSII4p2qvXVie+Nwk2GqoeVrqQU36rjRMF5dsp5v11I9GxDB
+wQVQbb92TGgHpMqjX4q0Im5L2V4uONPE2rC+tW7HGjwTMqXx8hH3NpjSC7nwgVs
MyrblJJ/0wYsdE/rIrYw79YhyBO3OLzahaNgv3v+WFq+7OtK3+7eF6jEfcPt8PoG
jfuXzQs0CYXlUakPyhHQgFsbR2il/6GQL19JgxOMQtknG3rGC80n4568JixKi8jG
o0SJzKP21KvjMU1Pq7OB0vY3TtsIN6HPwEmIovB4jllwjawolWhzbpO5WEt4nHrX
6m/QulyxR/7gohlfyiXA81Bg/JPLgUJRYjvAzSK1Lu6eje+DXIdzEXPVRllNE3Ka
WTxEydUYKiq4e9PgZ9ZBbRE/aFK4JhuYqOMOsDBAvq/Lrl9fWEqVenYS317FYeFw
I+dGzET9q3llRP4+XkJbTuczqmqZnr7SOUI5AW35BT+v4m/w6KhF8ZSIUCQeMT6Q
Rvdzxx1pGb4l1xPDIKLLBNtaVYMpzIXX3VJ3TXxU8dv+J12NgjAg0ghFtGri1wVU
7vnp17QY61R9bpNFiwnNyxL0JQbAK+0+nuNpdwIQM5xM0x0mGyyum+EEx5zey8vA
Rsmqcz5LTQAUi7IiHKmCPUbu/shUjY9ysPsznOCGP/t07zzivW3zKVp3kxYM7iTt
k6RI8yudlDXaHwDXD5lOWYADJ5g1XqRoHd1gL59exa1pLbJ8fXA6VgKpdYVzRF/S
mTp8QsPq2qMWMo7+KCFPvWmc/uLYBftxvrYtl0P+E4MCqO9ywH1POmG46zT+PxJU
LlFAnyHVd83Wx5QIJ/yEDcgtD1DYqOV7tmy50GrJaAyw4BlH3xzEnuMnu3rMUaPP
RrIah8vZZynnC/mS+zOzQ9b9MyxPt+8qZavj2BuFdJnzvZdsiEz6rSYl7oXSMGe0
L2lC70RBSICTYf/t0mGkTWUSbvXmK09++Upw6/8KHXq0u70QRHfIBVAf4yzcoKSX
XyLaLiVh3ScWj505LALcT92DG382JNLi2YU0jQVBgw2pq22IlNgxzZ1lTX3OHZ5r
ERvmXXmzCgFmn6vhGwZ+nyTJNK/D8i3qE8taYjVhXx3TmNCGUUqnaRu2X0ncpq1t
QsL/yLPMVVeZU6gY0fvjgngGKKR3WSDqeImaEAhW4Ft2yXT0cQEjkKlGq+OTkIYD
m9NEg3AQq/RfMMJ7G+NxVNa/lXUw603nv9DBAZyK069Nu9iMOP77ljAZ6lrRT9QX
3wnq8aFRXX33np85kaWY1OU68707XmymN4ENubcSEzoE5xIAaikpLwKsbCSlnBQe
lZ/1+sH7NA9m5jWstDnpYayAVOVZuHFER9WwM1uogDn7GCpcQvprJJ4+FgVhpKLW
/261dhIiNXJ0l4L0MPmnsc0MK3fXqT9iNkNjVBESJFB0SK0gj4XxEkr6rdqsXWw7
/FsqOpRLfBs/WPp8gkdysi7V2eW1WYVavJ5k77yQZjjx8Hz9obCgz3c3p6Jakxbb
rK6FXiWx+wN99KhhtrJO/+naO0p9kLnO66tpse0UZfbNXVRzarcXiwWCp419pFXE
zB4/8cp/ineL+wYkPNXx7VCzN1jAmMHA4JIZ//3jy7ib8EiYA2teuBzL0nsCriP5
Uv55x+J+vlijBsbo0g10hDSLDdoUZZeBzQ6Em6gBJvatQTAyGdZw687m2spGnSk6
ApukiSqa69BYTJ1Ty2BY7ZFefS+1XCoN+fCTfHbSAmbZ1Cm0I1DSw1AUFnFjpvav
OdsNJe62QbAuHHhFyK40YyqNUswEtE81GhdTjL2+u0Z9AaOijcXFd2TFS7BcIPWe
7MjmFOBGdu6+Vy2d/xu4i1v68gUJVsnuJExMT8TiAl3lH97FYuMVpluLfp3afer8
/T0CyDQWFg9DYNLSZyp/OZiyCnGjMKrIn5fa7/d0PgxWXrM8okX09e+gc87g63n4
JMZq+40l5oqwdAtEoQtVeI3tkZW5NvV1XWmajRxoJgPRqpZsZobFwA1VXSPI5BGa
gnzntKwoFVy+aWkSyznTM4sU51/19cekBJrA7ECCxdkOtsC/ChQuYOgU9qw/Eljm
Sv01Gwa+1MUukj7Ep8hfqNWo74JYzrKbvkAnEqbVUFwXw6I6OwWSXZ+WY9GvHoyu
LeJQAOWsoylu8u+AUpJAKXMedILmKCNw2qHaOXHwhbseACpdsi2DpL53JF6G4ORW
SbRQU2zptsSUNTT1UlFby6SjkuEItzYHkPM9MaNJnB/iiqAw9j4Lz7bmfTjZjkGa
r/0d+FVTC2eKMJSvibH4notsetAurrkk0khy7qEAUTH2rnweqf3PiLXmhyo4iH3i
CaMm5rhL/NxABDB/ZOzzJBsVFWsL+/PWhzyf7cijcb7SfWyg7WaWZTPqMhpS0/pU
JfbCVk9xRtbDmWEGCB5lzzAasJwisr6UjdlthzQ0hjFiRgkn+F6sXdiPWgh2670t
FIEmDmlvjV1ZZ1DU6TF/K4djnncCbudf2u8I64O310X3hzQ8X5k7ZdMbkNhEUXaF
PI72bUD/JhaLC8toZwyHD3JiSeu37Haah/Bw7XcUaFECwkXZOwmpHt3V/7FV2Aea
g7dZCsK3kvGL2u5JGYs5YX/6+3Fc36gaeAHMO+JypKT+T9an0ktgTYGwRCW/Bl8Y
3+UcUDv0N92xCWV4Bkrbo2R/ZGWurocSzwAhtfSke15uKo2Rny/U0AMxvekGrfuk
+or0n63LBTrZZ1dZdZwo97+YjIeUkDMsngfEEOIAgNO2UiRRBq3mwapgilnDhxoa
TMRe+nncX2g3GgmEM5Ota5+9qcnRDR2j70qdVCS1KSURD8RK2zEvc49e1ngu6EiI
HFXH6qhLn4c9yOk3iYZnMigOurBG4S/V9MnABLXfIrKeMbMfyzk2e6lIkMIm95Yu
vaBCgy5s518tw44ae4Slz2pwUWhPDd6/qqQtxkKro+S1XZmc1oAXX/H/X2S3uldL
ED/zY6IDK+HugTLAqBzbQE9W8g9x9UeivaNtpbW2hMSXn8HLH0mM6E3Zqpwb6wwU
tnKHgHsUsWXv0iy7TkIfkOYA02RcfHCkpfnpIbl64oDn7ns4yY9yHar8viuzQkDo
CtzkCLtTVkFSoKWsbokwH9D6zj0IBJs9ud/7oPv5hOosC5p4rNCE1vjqmcpIronz
14lHcDhxpKcS3Y9EbcQ1EEdSrrtfzP8Z/Q+xoX9nyExr89UZwGk8Aoe/YrYdkd67
y5YmjgRt7eui3l8MseoJz8GHtl/C1HCQ803URxrt7bsosifvdrkA07b1ZRnReRV1
nN/i8j6rt25hIgm1EoheM0F3JbsBfkoo0EbAZMyDVRSezaH6/PNxjcpMlGvnG8rY
UyB6ttd+IpRUl7JZz4Gijy9RrYVxwOMwWazMeeWdoutl4zuwhSK+Y4JTwC+fTJ/V
6k7KDqllJgCKGhGxY3DGE2kJpgq/g48mhPwj4i1il5pJ4JUjTO8MM8qS1lZGIETs
O62YJGHMeGGqinFMY5JhJEvByZI6U6co71I1nF6Olczrmt1v3zAqUiUbQ/iu8nF/
HFlHeJxLEd/rda8ywdYWsyi+ZawkhOFo69HIkgFGYRM5YI43xqfVIg/9cckPUZCn
jTPuT1J1wnM+JUqAByOKPguzPwOeHv7FiwxC44XgW+1Q2NBf2yqZTwGJZIcz4ddB
Cr+i+6OHivYBSqY499sQoyaOr2EtZIs0woxYDPyxRGlr8EKgkpgqyLK1uWtjVBbj
nEZilaeNzEG8PM86y8VDasxgglEwvANV+VHmI8Elg1qmHuSFgbRBlrLp2f9NQTbQ
Jycr7ZRB8ZoRiwEP77pu9z7RTvhCrSsNTWM9fSLTvCqtJosw+fFb6sqiDXdnhXeb
e6yJ7N8XUB0lS2MNGmcioE8aIYmYdZSBAL1lasZSZyrV8NJhqPx4BNAM3X2f0eqd
zqud9Ul10pK1QhPwQZxsGgAndxkVsXcA7akSF4O+ndjeD/7VGWWHHbtX4iGjCe0n
5Qtkee+V/xj+0CuIBE47X5jyqAynEBM1ciygUyIGl9pG/GslzdsxlzndT4PzOjnA
HIiG1M25hT9F4FiIctnq1+sQgO5AT3uuCXfkh3vKv7VJzwQmYiedw2OaLXv8+OPm
hpxVw+JX5QhwwWSXZlpm3DhZzv7kYQi/Zqroml1h+j7i2VZuq5VZIEeuezz2/2PS
uvUxefeUai+WDx7dsYHD6FXmF82ixtF3OJSXqE9SeyxzphLLbAcZeWMN0lCxA6KB
fvJhzv1AsYTQUPDRTQTdobQQdcTxNLNKxkHUyQQDaAPM2eiLqQwJGgskZFpy+Jzu
EF9gVsFMSIkFM4ZF79gB881E95XBbdfih+mjNC6/U4JrjZhnQqYa8b6LB1LzZsZS
5KRYnKwZEb4UeiYZOA1H0l+97NtzqRk8ff5ikXNyxGIB04xCquWoJiphhFnLzv2r
/6dNO8AvhZvMc3coxiWJHltjYvuzx9fbb6ZvwOQGjAZoyBiPRm8FIffNx2g2xvMI
A4RNH6ySX5Vj9nmmKFrOzxrv1SGlHzYhsiUopy2TPku6U1d/rzdFNs6yjP70++eV
ZB1GaIlOK2e3lzN+uZE/syGjqGHpaCSwHAqAWEW0qopWrn2ygwT2jb2DEM6y9kY/
D2V1YknH7/26sm403TTcDJDw+wEfaN3BBnlZAy9g927MFc61RBd29p/HphlaNZ6n
RvCWOl/a+kuXV/WD86gpQmSNTc8FyVp16r/EP0lrDS1q3MWW8Hsn+Km6M+7F111+
byDxoZVduB3597kOQIfsu8aAaX4LjXDVKCWRcwBN60IkKl2GOk+3muM/1AkIzlsS
KtFOhfVKtL8MtVfrCtp/0xpD9anbupZvlaAz7ELaGkV9HEiPT8kB84tC6MapVMSa
Y9HhsWGoKAxndSapYsz/x/shKv6oOIIj2AlRiUKXOAuCp2/LitSDlHq3C+et0Cw5
wKFc1bIHEjEc5dWq5tpCxpPDQZjOQ9PNple8FUoFGTwNheaS5R7mcVRV/xezztCU
xbjSS3qOUwndtenbBxPYUWfpX8qfJqF5a6SGan35vMDrP57fwCq2wPvwcVLG3Mnk
7YSFZ3Oh7cyjLNHRM/7PvWHt1/DYS4UyvjUVIEqlo+xDu0HMF8OUSCCMe2nP9HK5
FRdKKoBfnSaWfLIM3i+3oFayzZe53vYnalr9+4UVUxEY1gON4ulF9Yd3t1P3gIwQ
mzNu4DWo3dqYFY8DLu6eIXjoW8gBwbi6h7nBBFs+5UCrlQWCYb+KoYWicuZGKuYC
/NDTtqt5NCtuOxrOwRkhRFO5u3+SPtDoSvXBUkCu6HFJqU484hgICpWbYE+SlacC
9+U3yK48UsGT5Xpe263a4aTHfiT3IeH+AD1+Uj4mmj9uJ7VjYQVFEqpxHM8jB9T6
drHPNPfh50L3JOE6sQxlDgL7C+M14ibj740SQgrM44p4BFcM8OuUZdVqDkgbxLil
M5w3S6HyinluO112cKatxTm+3fJkO5ozI0ZXhHn/iMMhkYc3btaS0WrmsOmfCr30
IBZ8qEnCTr1yX8ITiD4+gdImRe0KZNjUxbgzQ7rXiii0DR9LW2vtqfq1T6A53nzY
LoboEb1Oc3/pDLhXA+87qb/yJTiBXUI9j/7KCe83BSf/nBh8xIMxvmHRxbiUZIl9
3O+MYfkqkiyNri4zngJTqqaAgaVUrB1fMEOOSaIFPT8YQBLnJh2YgmnH01UA78Bl
uTf8RU4b+4FxbqssLP6aNgOAE7kvTNyhX1DfhJ0B/gT2cVc3J+wLNaONdoA+p4mf
3OmfLU9mRz77+L7RLdWomlnjhIMvxOA6h1s7mh46YpMiq8nGkeQxLic+ZDnVgOCP
ryRJdXHkwbPZ+/U/rzDTVLhXAsrKyRWZMR4PsHW035LekedKEFvOX0WlKfO43CgN
ggP8l8nMl+ZF9dQKYVLhcj9PZJFTrxjvwY0yeWMqBYDDFaAkY1BDdR8vGSloee4q
5mydhk/Y9iFMDBWP+5A1P4aso2M0yc/pd3WrBpb4/pnLCOE4ip803RJvQpRu38Uy
ZpCOgr6TPfWrT+s9hVtobSMMOk4lEjiwcTp7CAIhEhE6PuWijuLDshUUbf4058Ua
nWYLyGIlSWNZ1TU8rGkVagHWsZ3dKAUmCyp93o3JtFcu6dfLRW9dJyKQYBPctSjW
VZn/isgto1zESqR2eyd9mjzqYXKbxxiAd4kEI8j7LK0WBufswtBrRlEs4rqwJ1yK
Pg07W6XYTM5JnXokdKKxrvqfRHqomG2+ANJoZx1ojHYZzKZDsJ88DbA6B6M9DRSg
2PK0zsQPWjDyyHmG4GhEcv43/0E1duI0n+wYSWj9KjtaCwm73C06t3N9M7HDfkgV
yEAFt71qp/76n6lpw6S3Sn/G5x9BQAiLbkGnMYfhYHWio/Fd+HBhYzjgWjCT2Pbu
7AWD73EtUS1ojasHfQoA4WXfTmIpQ0WLJWqwWSl3cJEsJjtnz5WsRlhf16gy0Q68
jkmNBl+f7lNtSH2Gm96RYVa0gbHPqYaTbRPhYiNs5ZNhFu1NG5VDXNjEUmJf27te
fe3VInnLuyYj8RYw+ETiA0IIWa87/sCNA5Q0A2hTOVUqXbGFj0d8BDHAuEN3byko
i/pd5azbnbPPgQto6C0rPl07VsGw/rGLOz/hjamAKXu8cbOgOy0xQl9dkcwafNBB
kPvwrMqxzFbI8dRB5FOikTDDw5Wz9WJaTRWK28liW7XUUr+su7EUaKyd0SozNF4f
mu4/IPIIUtQ/7A+ZqpZkuc4oapm4A9WE7eWXq1xVGk8FWeikrtDAPADleTzSC36E
0ZTKm05/5npf0/MclFPjkFGBe31PN+SNqquK61rL19BJyVPyDYl1nqGDrL0vmLO2
fKYjCosXF+RvIKNPbzk/FaKjesFyn1iljrx3/rjXc+tqJhmaiRviWut9T/NR1HJn
c4WIHwsRYA1hn9cgWLwLCHVuuvrOLveMRK1VTKnHhXntSMPwSPeYKz9Ux4coVmn+
/4zOsJBHHvArCBFaS+xi3LnSOplsKJVeCzJeq2M7r9NCiK3AF+FNdiNe0JrLDbUd
YJ9F28pSn6juXidiB12KT3/YrmxfvhnWP79wCNv0eMYJQe1fK28ETlK5vSB+jWW5
MIqfIUz+TCP4JaHzPbi0cnArk79KZvgt7aA+mS106/sC6euv4zUB+guwDMVQk+GY
Ikzz2OhH6+17DCBtZypXEE8KSeuF3NwuLTQ+Jox7bDnA92Hjcj2e/cDUY1Ehp2rS
9vkHNpMaHoxhPTNPPDCgW0fsvN67+5Q4TTkpje8mSPippNlZ/UEByPT8xpZMce0p
jYSo1P0MpYkclTtHl1gD6pFSVszZ9tWpYD+PvuPPyZ9G/awJXZYMYi79C6rV19kg
bb2utj5zRWfxZfhq7JZjZcq+ls+8TWF6UFDFoqdosIaKlNboWDCds67tcEcaWWJB
twJaDLSDrVgp7zzUNJ7zcR3aon1DBGslGx137OO8lTgtZqTrEcoWcOQeWDwA0NVs
mG5fjBwM2ZiGJ9y2+T4rBpNK4advODR9oyskCsJdJs01GvL8D5TCSe1rUT/vJmxn
UFPCg+6Z/lLNtDEHhlHDQJZTk48PZOrskrRv7LD5jQ8l4RHnaZG1NBiOkxSIDWr5
6U8OYMjQl6nXis1A2qu30pn/vQfL47FTTxoblAcxf32dKJB0ARE4lZbBMpb78pYy
BBW7XQIWCPkslR4ie0ELDJ9Q0QWt7N5nrUXWagSP74FH2VCjSdn1zbqVgfF4VRta
RaG08XmKx/GcWdoG74SsAwDlZDjeYY8uFeDZ/ZPwr1goeGmZQGxiBuEGo3A4Qi2G
PvkqL0TSBbf81uAS7aZeVldrCurE8O64noJvivax40/LOpJOoRv4nh87NTRb6eGC
b6p8jXNVC8oKpUvUOY3HGKnodpkoUEdzfsTxPedd7NQK+jD0PFbdmWN00I9lArm0
PMkdsMNTiorVbfBpe0GjJ2ieHKuJGJOLU/Bxu6b+qs7ipT7wt+RPBd/cYh5MN5VP
liyIdPNY25poJ0fXlDYtUb0PU2MadBirEewX51cSkhoiEI6v7oUwZxLhFrn5jZM0
fsf3WjBbnGE8ofdp7tjW6FA9BtEOre9KImjfWbixP25vvCeIuiyxZHYR+4dPBsKt
LkJQK0E9JOitdYxxh+NIFEKLt4NBySx6ezpzBpV/7eIcknesQG3R1O9idsHgrSc9
RYfGKbRVxiSUyAX9qO0Xf4gXCqmcEMPBplhW7g2QolLDj18Y7VFAkkaIQZSUndL3
N1R4yiFwFpHaGKNrVBi+4M/52WZH3IW/S/VmyOw5hhlgQJgMWn1a+/5zgSDyZLYH
vDRJs1CerF4kZ6jn2P9HhL/FMt/JFuYoytwXtA3MAgy8ikhYiZTU4gT7TsLQjrIv
AArxSBZcp00UsDY+Wl0a7+ALVnM1cbYA5XoJv5435a9Y2iDZyjrG27sbsekcNFLc
pRySoM1sE0Tzy8Ue1nGfc+Z5d9qQKlkUUB6Yel5bxP12/fut4Ao7riXs1JeUyITH
FoVSE+iyvd90nqY/reDa6dwYURpQcMgtEMrtLdY8k8hl83O2IlBHT2fWnhDYB2hQ
B+yJm2Sl57qpUJ0REpXkdDV40DjusMRJCqBUtXr+CV1jgP2eeLnodjm6DbMAULFD
tO0VCjR0i5sLNk4LEu3uLgrXMU8xfFqQH4BONmO2Y6wq5E6TMeA6K7bT617iHxh6
m6WkmqmH7lhoy+yWbmdudJiIIoNNHedxlFBz0EjanLtN7ApZD+KmwWYGarrW8pEt
uTe4TsjMDPbgoi4Plo8ds7aoQcDt4c7EdVIx/EmfF+U+sojFvlCbzAlE/NLWf3P/
cnWCBqYOkpH81CY0dDBvpAauMdPXdwdEvs7j1ASTrerOItDpZLY2HxUOIKpcuvsr
9JMzhJceif+9mM4iR2y0yXlxIjAaTcrC5Q5GTRzFMokQYw7Pek7wM/5GbICvBS7D
wykfDtmBDygKg3HXFYwdXe89YRoOEFP91Am55bsTTO4XajwnE6cj4GZraHRYzpzt
Gfew2kEqLmnJ3CfiJKajywJJMhUZ0JWQJrdqOYlF/mTLeStI7k0qOWkeEH7W6DrF
ZCfM4oNVAw/FdDG59TiXm1ekUQCzpjPShDi9cOW8oaX1g8laFuaNCGEZ0nuFWLlu
+tN9afUGCW7vl9ZtmgZThLB3RqOXZDCQeIyFK5X6uD+E5DMVCwdj9fhbk0alcrU3
NVDmacjtoJARYhwLq6zYw6GejXUwYomlYa9hG549UTe6NINTA05CSe6hpHioTLup
ez6KfwKfVPMMVDhQCZgDxJLJZ59Pr0/d/h2LOauSt5ppvnF6Qy53/2EVeDCegxkC
9/xwUmKC27BMoHHxRrtiqv6IhD6Sb6vYWBs1jAkdhxUAF6e4hz0mqwoRA8Bt5t5P
wSQ2yzENRwOAGZcJMJu+aKaWFNLAkEnndU+kt+93PZGZuE5CWmaql4VAlIcJ8Jxf
yHK6Ci2yL0z6Z5J6ZFZsc332t0JoHYtd6f7jAwC4vI9Nyw6DRiRZqwNTZko9h9KO
iYuubGOWUphEEmYNiELeqiVp1vCip6LCstG4Te3ozvHWcobH5/Cv7uIwY5k2c4+Z
6flRJFUSJA5iQcAdaZ400nJg3In3eaS06qA9ZKGepVaXBofhqlYK5F+yOHz00FLH
+YxnnnrXbQdMx8ojH5DeBES9DBr71teOPjoCqc5rACjSgxpeWvrWIYh+6mP5gkpA
O7VvgzDgZVW2VpnN4BaSBn5fCyj7miQChqoasXVsg2s6dK7Kd25rmYIoDC+keH7I
0NWN7DfBvJac8kLOUCHQ8ep6R0pAPc6J1XGnoFyYeznmG3fX/z1vHZOcHkkLiDQf
vD3AFUKAD773Ajs0lo44bEbsSiyiPTOgyvTCRovlYDeJQ7H4CoEomGAH3kjm48by
4XbaGIY1lN9/LUcSmPGXfD+BDO9O0We2IYN7pUQxnS+zoc+glcbdtp7yNXLvXAYT
7grZrATbZ0oTduocfBl+X+a5/BnQ18KUA0K9K6Z+0rSXvyMkjJTDh5lDsAWJ+TqH
mgZs89ZCSBPtMvVyEPH548ETQjS5q6rXoakAZAeUCbpyTYTALhERtfBkax5xQUjd
FOErZrE+WEXpWgef8ZtzxC/C3oG2OStyl4ro60UcOc7vCwpg7XBs7213ir1WGN59
qcug/LPPeLtIlqQq2XTsnGnRSoX2CN6qjwp+22EqGzRSIV2HhMUDZmFb8/JfU1gX
sQB4sBE0qLAoGfxPMLbRQO3+v5mTRbuJYz+FK16luChiLHjqHkyjOfaOVS8zwQPo
AkafQ0VD3boULgtiX9k19gh2tOe+stwwjq1Wn6dcODgYP1VhYDzWkotENZEfiiXT
qY9r52GV10VYRoEmQLf0MkGH7Y+5AK0M2VpCY/dJrTNXLQMXChv7HgMiLQRdiQg5
wxzd1Kvb5wrPHLOlvvDUZPUv4IvS8gUgNRi050CCIUuKDneiYmdmz6U/crVKwSUq
EG8GWitfSUIjS5/qD0lAjLhC9Eap6oGydB6sls5bQi67r76lnx89gHElWmomqyqs
guSpCXg/t94qvr7q2aPYITcukIijzdtcZUx9p7pEUq4gw6/rV2lg/fSrBKm6kWyA
eThaN6KWAs4zoEn+JnYZU7ka1YNLzN49TXC6AskjtVoVs1EU69GDiR3yt/jZJJC+
`protect END_PROTECTED
