`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
TzFXkQiVUTmwk+uNsVcbxJ6X2sL3mpAvQs/qJaNHcxJ0F00OHPa1WobI98Ikwoky
P+hus0tg4Mso4RgI9NAbYPL/IFC1Mwugne4YEPM784mdPu3YwQ1orw/NhNcJ6CCm
yHM+CPWwbQLh44AqDop30qX1AH/E6OilrWDhfZuNxIdDLg+XH8yONJu2K3VukubK
eW1fgZYcGUg0FvSz5tNTaHz8oAS2wT7/seDxda5Rw85dGNm9APWgCKynuSVQu6jd
VeYh36Jv99ctYDlmLfdsd6HbDaQO3dwfScH0/XaPdi3C+3h3INo+H56XZdN9ohjS
JXuvN1faAH/EEuO8hAW0t/MeAOfF6aPqIP2WKBX3NqIIh7JpSPuXLbyJeVmhY9EJ
seM9VxlL2CkyF6etP0BH6+JPLvAzPmIs3SynXIhRyKDuAvK1F3t1i/fVal6D4rt/
jPLRddPzyADQMBiPt4BCr0GBERoFAcAeKFuY3l4SzO39TmZG0FN9S1Icahm2mch9
RQ//VU7jzLODczRgnhVjoqD+bwu2Yg9uCZ5X+ra1cL68n78YttKN4TYNOPh7IjCc
eE+ui6uBHO4udKZIsZi0WW0pOw/1z6niTWvSi/J2MAgZNN09KMZ00X/USgb9HcnF
4USqrP+mkj4uX22EW5zPT4+QQwwUTeCTOVZWEPMpbzxvNH+y+hjJBuOAvOuBkidO
CGQ0coHI2yDJe+9GfKpyMRjR0BUy2MwNp7byq30/lp19PagIi8gbpsIFtgmEuDnZ
alxLovGuqTLziyfMkAmDnyXbhF+rMUdhFM0HqbuLsoo3AtRL6t6QvvXppO6+FMwq
yvRYuj3UK+j4VmQy+vDTs7W8ciBmzMCyVkHkvchU2op6SSFfR3XvTcY4wCpEcmqv
8KN6jyw4Ct3HZO5jcrn9ZNEVo6dBX/+9E2Ek0Pxac1d/me7OAqLQAqPcxyRWFLiI
FWqvI8vTzC1XRbFECSgYZVyonxsRCLKsqcnhRWqzRbXT4WOGutoq/AvcM1BgUaGd
B3VJknZt6QrGCrxyj/ezzhNTwkjcQMfi0hrK0KnPohc+uzbGX3ZkXjn7SHLd9Ua1
lZ+zPO4MzKXZ4CgJ8hGic7PqGYb3VHWgsBcxl2u+x2xx/ZzGkMuR0RGIbrR4npg3
JdL915DaKmjfocv55qPSUmJO2LkG3RzS7MFP3S7QJ2hTjAw54o4e/H8gmqhgErXf
El551v1PZpEGaqWz9kMmICCeobZcl9bPLENI4uZ+84frzNyOadlRCzyHcfDDh5R0
KibR+6GNuMXiL+vpbcQruqOLZESn9wZi8A6nSIsB5oTgOzpKXu5srl7B2R1fBo+W
Pyr6qRL/lMXJwy+WF1yF6Duwua7iJ3hHLbEDA5eqVwy9b9w3ZiCuBHpNjq8ooWDq
5KSIQfjQfJdbqeGU0k17gGb0msbl5nKExiaQ6fiz2WKgAcbUwzESZWqLsf3dgF0o
vvesObMuD0fZvv0ot5TGEh6wFGl9wIy3F3hZOaw2GlIKITaNqW4VU3KazINaaju2
NLVvT5pBZXF1OhQiycXhVmWDbznF8/Jg6q3DabmRlQ7iKUD009pKyp65QStVQzWk
Gft4Stu0KKLuqrLyOq6wVzpnKp/SBS5WDNWP/D+u+I6TYJ0i5vl8V7ybsBejC4Wq
P7FEHdrYX2nSM+NgodrchoDLBOGDVAf53toJhSwNNJqt+9VRZUD9O1jNwsArNJQZ
VU1M6rt1WyhpnonTqjLsrvfBp3lKu+3uvsODHaNPW7gX58gZLZbSjETMveLAA9gs
3j60jxAYFXVNKbwgwrKRVVa8LhoeAAUSYZD+fy7+xHHf2Rkd7bRGEG7r5gEtL7co
6++mmZQtMzw+HHPCvYP09izVGa3pwMIkezX1Np+J4s321Xo495doEVIqrJZGOp1h
g+hJ6IKg7wcIzjckyeF4+jb/OcQJGBsSRoBVDmTSPojqy9WPQtdPwULJWOVmiTN2
6j3hS14YvU+UVvNiTyxp2Y/W/+BzE4GBHd4T3bMbpIQq+IKKUjOjie7kDohqNcRE
J8d+Ve9tmop0nNS2ZryS7UTCfBlnfi4BB5XEn98ZJ11MGNPfEdMu4Ie4YXg4KXLI
AqUqQEXm/hLrxXZKzJo7QD4BlckFZ4CFIH924NrsBU1E9CEXYi13U9Ss/ZKDYUlY
gPg6K2SakZwyWumFVpAtunTgKJIYLbQISZLwUuCEhpzb1PtcOIWWCMFSSeLzqCYV
1LpVj+QBLHJ9+EHPJJCMwaIqM0SNCHjmt8SnaKHTwpAyT881bAKtbQ7dxDM4JMuD
jMCn42rq34nY3V6c03qMCdoQmAWUq9XabRPylpm2a7gwUwXLzFtX5rxTfEWuD2tq
87dUI0oFcX2xfD1VUpKYBNoOFrLNST/zaGMtAsbRleNlRnk0CENnvLcT7/Z8KeIA
07OIg90ZavGgH2Vd487L5brf2S3aVPOlU7yCsHer+fgnjL4kDTq+Hz2/4Q1yE+jo
ruJhXz+lKCxDDdjB4wes0/km7TyacI0PmVGIB29ZaJkT0SGGzpwRAWx1LnccEhvI
Iveil1oC46a1ev/9LXeYcJRIR7C+xAat+3j65khk+n4DrHn1GHqwAoa43uP0ldpG
NVfC8exYCDiKrWVp4vO8s/7P9XRMsUV13dLo0YQ2bv9kFW/Q0TWPHtpb2BSAO5Nq
K0y7Pzpy03ldBi48P9EWOw3DHi2r3uOu1UZVJ5toGBuvvXyA3A0ipXPJrbyxwN3E
VN6+GysAI1kyK7yHxQI4g3qDxP7BeaiIyQF+DJvOSIqfsYcRdWuRIu+zTnch6lOx
tzRno1KPfuT53clFVzoyQ2Di7lI+P3c73nM6qvUtGTNLnRN0REkqCNjyov+t7SIX
+X/Y6bwubUjqHeFillraXboetyRE5F0v/Y7Sp33C+bJnhKY5Ao9aUxmoZyHirhbO
hudVjyJygCDYOMwG9I9Q6NNLDYCjzsbdO7QVmb67bxBS6LBFFLW04t6OyesJ6K7u
Vgu4NXAg+TiTL65BjrxMvc4rNBEMrOLjluvGZJgfi3MAD8WX0m3aZZolVA1rfodP
ixRPo0ng4cOnjZ7cp8CrAzpjhOMuUu5s6bn1Xpf3EPHx/QmzFMl5A5sCvBnjm/yH
xJPP633b6+YxsjD4y2psm9uHDE0iugBXmXnONoaw9vjAI61Kz3SS9dgLSwz+/9Wk
89v7oowxIONpbTDxz5OVSwIq2RWXbfnvaxRoDj2ZPn2D+xl5/WuqdcHdvzoljoae
vQaFkW4kQR7mu0aZ+3pF/f03FKlHNdZrxv2LKqFw6TEIJLgznAKkKGKRNroKxDp0
Y4w90/GTZqoK2a7Ng6vlEu78nnh4an1pwzw2GOWhb8lI+tXoMrk9YsFC2OGmFg+o
Rj/TMYerHqCb8bSbMXMqLIiUSRBPqG79o9lwUJciEta5Nax0YHmNx+7tRtVYUwL4
cOFLEjPGW85mNWYR0DJIp7HbgFStgYeSuTvhN6VsjSALySTm2oH9Y1WOh4R9StLS
Z/no9WSnmA32kPmK9c97PSI1xw5SgWPBYdXl4VA+FtP9JPM+hlJAMWrpyZyV5o9n
tf6XfldZUknQv6om0EJ1V6DaCJOg6bICELV+EsngAFToTwxd0tDASp2KIEZtWV8x
6+nN4VtqGAxK294kVDVhkgvBYHR/y5sIeJCbewgqqLLy3SaXeAOcEBzN5+FDHeUQ
k4w9zmeGiuPgNLSzAVlOaVHdzuP/ehN9s9eOr7FOgqgulX04Ta5lNQouyKLnuLWM
3rWtoyZ5wt787srbVAFEOdI4xogtQM4V0f2+v768HZugWXvRX+IOxKMXCFL1rwKQ
rTMg5xpxaYfMpNi3uaiKjI/mlDw4IIUyYAzoNseYwRBVaFMvTwd72EmOaMv5V6Tv
yGLy/zNwWOptI9BsMf1NLPit4DRr987vPeEpd6Yr2aYYTb0KD5ng/3IvFOIeBRgU
Lwo+savPATeT1eE3OZRP0cv2UBnU7mXSzCUpTTqT5L2eMiALAomPeNZoKzaEvvIA
0FQPZaavGZiT6qYTiKqWr+yf4R34t2lRf9QVedTLhDc+jmgABCOmpjUkxQMjoofW
IgZyjGDIDsTVh4MNvNwcyjNSkASFbf3rr+TxJhU0pKDk+C7sEr9R1xUMCzTQ48w7
CqyAn6m0203qXxov0DwO1I11d/W5iDeMvJLxEd3ZtkAlVQznHqowXFCeOsq95EHF
lgIDB7rHsm7N64LuiKUstQp/zUylByFO5g2FIAvVxpxROP+h0CSkLpZGKskwxKmH
VqaN7xaE22EEw8DAJxizsmBUv9Vvu+qNsMoQPkJSN+k8AjK8ER6DbBaD1F58te2s
SMbYIlImKq+DWgxOJs5PxVFfl4YixKZwgK1sYsqfyaSWwvgrZmflgKyq2U3OtWtW
yNn3Lgs+5C8/mT7f/c/CAD4zaVlA7pQnjMuBVubewwXEd7qUkkUfvxUTMVFiD1q8
OE7SSQ7hiaKp8LO2eXeG6a+Xu7fsNKh72/LKn3iWVedpsHx1Y92g7Z3m7jVK5C+Y
O6tP8ViYs9kb9rvCiE1bjLogyy8qmmhyzucRNvDKDkVTgjkSg4/vQVSqWLXWxiFt
BJ87cHoJ55UHHgTyaLLcYvT4aAofnxVBAEPIILIDDI4L83208rANWOEiuMOhwxun
GvcxOgELBSQUbCAL2Y3bDYEjdT2T7/aeQ1qTjitr8fidXUUJmKjsqOATE10jTg/z
g2g00EVqmD1nhWhltTBb7/IAsYR33MDpOTaE79ldwaWw17pLxmXXKZ8PqX3vjxuU
QcBDP8C/ZydVznv9K9lYdZkCZFATzQ05HqYoqOPXyKLQJMLuFRvzYW2U9fMkoEaB
FdcaFMyNUqC7dEw12AneMXpGTGx9wJYcbPg3MxHAFiigQjWJsA6FGfwqFObArCvh
GfCg7LoNkQgGmDYLNC94Mg==
`protect END_PROTECTED
