`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
M88qSJdwBDnBv1TaA54zAdTqPuGq/PQDm+jkeRMuTI0mgfIqWbxZWnMXouVU6ism
y0JWWBWyp+rSuDkK3Iigl7b6Ur4Bx9LziBdRRGK7UdS9xMScv4sOEFX7OLMmmF6P
Ez/OhPFOgFwgCSJnxngW3qaci9md9D0fL1pND+GbDih2OYonQY4oqzAH9bfQYGWQ
bZd2L7pyae+bkJHlNDJEznYZwKyOPdDs02H+AnnxIMu3uCE1S1eYqpfUUquhCHRb
QHeNiqKbq84UzVGf7RQ6crHEnQfvJB40pszYFqDs27H6Nsc5wB1rwBG3b072v1Hb
jBlxCmhY2Xkv5lRpBwKygCW6xQN/u1TRt69jfeM7WYOn8j7ulI35MQjKl9Acq76d
BQY0vu/TTCzSPK+uW+LdsTC7vqvfmHpid+1cH4LQXfAyw7tXDmO5JcKszTeJely+
`protect END_PROTECTED
