`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
BfrkXtfM22YFxa52gOtVq7a2ohSTdpnuezqHnuEowMNfTkRBZp3NrPmP52lyQDze
9f1YtbnPuiGvqwcwT4XGwi34eYoRqn8vQE1xJSxVQmIKEDSi2XKRHwo8Z1/s71hJ
19KJ4/ESKLPel9Eo8XnLI97sQwgPi4mG+kASv5zQiPk77tLCI/Uo11ktWrzKYTqS
MAVrQfSEFmFhSWM4UI2O+LYTt0EyHcFMByoa7F8SpLtwKTksrwV04s3IXFsLktVk
zCDsp7IpjE1ZmTo4aOiIVpCZS8onQpPfWtm9RsT2xXMy9WFBI9wxB93vRf4NepfK
9De/2vtsSwKh1VMLHAkVNnfGj9h8OccyCZzybIaIEvIwxHcRqXpS9VZ9U8aJDAIQ
yAj6MzhoytI1bk2EhXxzrrAp6QU8vJpO/+cHS3yz/hTBdogOMnwoL6kHcsSQazE0
mw3bIjk7E4iMWmWkCkrdTm5ytSxVrFV9+7jaz4MDogAOu2X516l9c6CurCItIl9O
9vwuHYaRGYwpB4kC4uYpUoApRZI94i+EedWbl8N7o08mZ/G4SBLrLSBQCW4jmTSy
jWLewLBivonC5UTgtN+QjW5mpHzLlc9gMiDJuIv0IQZNcb9Oez/J/VmZ5t4IF0mV
tWuom/qY+PWw/WfYbxUOzetWmTKk0ktZ4TY1cNR0PR/QI7ARLo8sFvFXgYgllcwB
4KdyX/1LSGIm5OgxAmK6MnOTnzR6zTB4w4lCZzmHUVHFJl/SN227nshhuzlI0tOm
Q5cfuzZ6JSAfGF5uxSyqrgtGr2IlS0S3MjMbRhZMIvXX/EBlOpbdRG8YNYY+g9ha
kISYD9a3bAt31syuNacU59JtUyRNo/KOwjWjb9Cfk85tscV3Gwo+cN0I5hN3L6Ba
n3NSuxCOBHWPIduW0axZPk2TgIoPmnVYOP/mJSkLg5q4VSc/3TDyraOyirhP8F8J
Z4PXdx6+nC+T5wpCb0bk4rAXm3HW2OUYlQlN+bjKHA5hqKQoWPHL2LG6nuk5cmiR
xb9oFRmhQZTKivisvkA5e6K4y/2sW+fEyeX//zlApGuMv+yetnbWbmc95KHh3Iqu
K0lGFiYSoriiDojGaKbbiJVbe7MCB27y32ScPuX1MHy9LWWkC8UNBwQHvV6v0IkP
djs/9/yt9zeLRO5ckSBK0/cY8jjgDx83mfS3lGuRG03MOmPECNK+5pAPzyEjj6gA
Ra22cvPI5fnmgw0MKwJb7EVKD6BRgmx8FgCW4QXuFFPJpSc2aSkAIDQdvQXB56WZ
R5CAR3c//fObhk27iwuaNDtsKjpPEGoGs5IS2dOLWolgaTY4KuFYtuUSTbK9E3sN
g0K5etp4bTkgbfbvr+bBXVyxWcJzkFSUdwMqeSP+vGUTYVtlEO7YUlTHj1PEOn2V
tDmwDllCK9ckMisPDOqrK3mYbES6p3pDB90NoLDXCEiX9J+zVNwYH5zO0niLGNyH
rxJsmH1oX/CCN0shwtzZyFOTBVt6L3Am/0O5qllczJjpej3Y6qDNlfRB4rCHwi8a
cQdxt2WGWcyHWiJcjZN14YUbCFOSps2CjeVEk6EWnWS+Ks+nB9mleqPnYEKK80v9
bzpQR66V7cnlm52aH1LVHUBMKxRiT9ecBBZdDZYi2BCxU3cCn+VLXKbr57KlxfR3
HkJvky4edY6Gq0XCfQmyqZLwX+yykOtF2pwTA4sbIsxq8OOnjdk6FHq0+wWbuEsX
4ddckmqoW1PKFwRZW6bCYAATesA2VDHgyLcdXCyHBr27JHp+XRYbuWATU6jhNZ2z
sHYWHeN+G27SjwH4lVsToCvyMaKXtW8P41KRvvr7E97rhvQZLAIu0idPD1iKj8mn
e+F0pCYV3w0hNF1rAfG3ts/f70TbxArotKI947WEB/cqC0Ua858tlZA/8w2w0Njc
1W6UnTXEKzuOV3dugv64JC0eF/jehRXvUU2pS0Aal6nM74DNA3TgfoFbymNYooXx
A7gc5FrDXZ14MPhmHqeLyKdEqtrvv1Y1KNN1HPXq0Rgo8Fh6sgRIcYfBWGHaVc9o
es4ab7H85mLAofhbdyOIqSpnNcTiBQdJlYWJRVBKeFkYxFW91N/KUvrHAugV/JBL
rMQFbHtZ3LZu8Bc+3f8Y1mXYtP7O4zaHdxLpdVnJ3BcWOOJO6nts3G+dDuFxPf15
gVh2HgbO7seH/DdyhyQAPnSLv5Lm+mmru9kEDM/an2/XU1zwjewU+ZxcMXFr+wXu
KGHFD2j+P8k8xgemlydMt+fX6hYRuwYsC131QLrWDIjjIwfGTBl15zn1NxVgpxNj
jmKetLjan+9hBq+CvDzZY6TL5tp8roZnIfIBo5vm+pdWHdQdjscA+qX+fbQOPXug
m6KmTUQkvnPY9iO/Ez2gZeWc8r0rGZyv3ocDXyj007Hu5+OFsgCdJ55hNMrjRvjQ
DHN0IEAvvhpy3P7xZr+THekpnhagidzzgPXPI/k3fovRWbcWqVhdJF/mX9m0/J/k
gUT7sB2oVO2DkVZdYmf2xByLvDgOQmHgRDsxiwoWT5aLCiS+5wm4nfVAIxrJJEL0
wY3jGuGZViPg8VTw5VAaFncprV2ic9Lef0a4QbVGm+niNCGJBx7HefIvfRcvwfGe
vxJcz3kkXyJ/clZ2HvRGMCSyu2lRAEhSZplTcen6kjyDM8r036+EAl4j5rePYEm2
VmufQnVWt2a/FVAvcUx/8K+POY0Ws+fnQYpkc/dc4+fJ+3XOOroeuM6AbEiVBE+9
AwpeWomU2Qy4Cc6YX+88cy6h/2WtKqL45fIaol3gstoVLhUAYFjqb3CdxOfse7SP
zK2hazsxXW/Uw1Xhfi0ChRuLypaxKAHDkmQniAeu25ldR/8GbNhmLxYiCbGDixxi
DIf3DgMdJpq3IklAX5QHVNgHaqFoFTgYnTSIgnQja1NzRNvAS0W6osLlouKc2zj3
VQUpBhPYWRkkqnenOENhCVTyXGG3RVtCV0t+sHgMwo7yYpFFLqgXIbxbkL3m5hNc
2HVkMUKin/r3qq+Gxrt8XyUDsSr3FaqT//YPCXA4WKgtwovEPT6pri3uBgbI7Str
U2vAPHCEKwSaaMTPQaydGS2ViE2AVSiDxN0hZi+lYfpFNkCT+hmkbL2rGqWZFbqX
uhZCbypRz6CWVspLX+GyTJ/Y+/4/ymhn9c5hx+GD+ai5lMJ+4L0rzErYC3G+nmlg
zVJ6iI8OA68xzNtUy3svlO2QPlRSb0w7SG9Vf+Pwsg32UX5qaC7+Zee3VFLk9h8U
6EcQO2Wb3Zq1iFZufyu1s25iyEkld6nlrIP+w/HpfvptnDkY6yKqKS0ZWWoqSuvk
qhAR+B44zsHTqp0e/GkBfM5dXOX205/tCQB/z/2T0+sv6Q/+javZnn/oXlgjnJwV
WiPJjA26ExhQaHWRUzbqbRVF4GDSsqoGkv6jb3vUzzICzZisF4G5+Lb7FEXfR1q+
OzGfLa1HmkX+Y7pCgZD2X32rHXOqL0ZQmaZ4Rf5KNSjHHOGY4LJtWUpumm51uRrT
0bTICC8eDJI8566L53ekxAo3212Dyc2LfqpklwIBI26RTnyL2FsRYPjpqANZ+Yo+
nYS6CDHFnsGGIFbSTAw5Hwn+YqZzPhccZqJvZ5LSIkXHDD76P9izdxMCQyg/5Cr/
u5xLlSaWI2sKasPbTXfFRA==
`protect END_PROTECTED
