`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
2zCYHnoZfpc2CQnjh8y70nvFycZ+mQJh04BQ6Y8L0KPB8YN5/m/9aMHpbYBCUJOi
HBMeRctFw3Zg+3l+Oz/URG3QD2MS+kkDZgQJSV1INIhgCDKpXFrklfUU3KNfnVoo
WIs3N6uhO6ovUl0I23EeQpO3AJGTZcTOvH0Pe15uvWiWV3lOZhbcFIabopJcUC+X
1rZT9Kj+kCKn9XfXLTUNAnmhkOLd1naJqwvn2O9tBEJY17gV3JTLkoryOX9YJO7G
5W7iG7dkXQ41o3LIFmwzA6pwSl0dAJPRcOce6hQFbfhUFEwnU3hg6o2IctVNCvAc
48GYGSptWI92S3AUY7lqvtBTVZydCHxyKRf0Dlan4D8ViMqpM2ivwAuTOc1hudLq
7gSJ9iBnSO+HcEvYdhC46GgNPHVHgKvM6PsvK+BatWH22dXPoU0RHSgQ7PVKIpzz
rifeixCM6rViF9bIk1hVEtcXzSS3/pGkoat+pRbIv4popzuDPc0LPR5ReXgTnwFk
1wCVcQc8+5SGsWa3gicVTQquiGKCXOpfsx+DKQrCLzmME4nsJNHbiwpp7Zqg6EWD
JHBI19EqA2Qg6InKb2T4T06IS1fHXBTTwKjUdQqoKKKOADhXtRUmwjpuaIEKIJex
i5oz3FsWjhJhbw0anRBuWeTENWbIiC4w9iaLF45GvhhbE5ainUaVJyv+vvB77yNR
em0KzB64VsKvUdGrlnFWWEg6URSeXYziHvIuGZsTsxzDge7kEHmESlzGtKo71K9s
LKDmCeEUaf2YaWga8AY1F9+/eRl9vS7qobbMSNcKV+pVs+bnVy8EHuUPMXvEr5CY
`protect END_PROTECTED
