`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
qe2G4w0bVygWGghjjRzp3CBK/7eGowT0A7x+3S7wZo6LFX2ynLM75/VAKVMV9/zv
Y/d61/Y2XLqgHPCbXTBZgZgPjuoDf/iAA22MlJTIHbd0bTcM87kmLSgwERC0V5ES
DVWEIFTjIhnfCmCohP5YrFfN+YV3a+lucExjUB4WXaqqNq5tVeYH6WGp25Yj+b+1
TU73QsQozqa9HcE8Y9TKEhd0Z880sJlLGZwofOlZFG9rS3ksme0YV/6CBFKOg3T4
N/+Y9u0ppuqpDfR+nsU6o1pHB8NhZQJ5bT5y4f0g1lQQliVplo66gBRyU5iNvdOu
4v5Z/+67SwzYwGJZQL3e6mUd/3n7/yH4DVNqapSbGVRF4Q1zMdUpP18bXJ35lIaf
ZQ91xYnPAiW4B74FHMg2Q6EgS1Yp5xroC9El3u3nCPcBNdeFKUWp5fQvvONsy52D
K5kv5eMe+IWWgkP2wzUYZgpQgzBEqLa07QIIiqOdqggacWObOWGGRJ9s33h0cQmo
PBGofC/gp5wpjUs8G1LgjOjZpfEwLqr7f2IQVfdOhZwtk5nk8gXE5ZZMvErP2nJo
BOjlB8m0IrQPLmPdsqRX8CDxodSZXvXo1QPGKPh1wQfZlRP2HOf2iQa3dZKatmOO
YvmfsCaawwFdb49oclj+ulGr1WhK8hYhQjeIlIiI7gi+DwyeWGQtCdOgz1MQgcMz
+i2lxaOwVfDrG3TtUGo60DPL5JJa1S3ItB+sZ6yvcophUkW5SChDdQeNcyKSKSn+
BcdTEOHAA7j7AXThIgsAqDwD+YWP+wVFqdqED00cPZjpE7I5/3YYA4bxh3Ra8Sfn
A4sfTqOGtkrPvO5gOYP+pLvRNwj8kol3x5VNDef2euQZ3RhU0SbFG9xb5crDodU/
q+OKpswTNxJLPSdZTtGwYKr502KxgsoltFMeUPiKPwcoL25GwINJ2JmOVde23nYN
S0Gh27KTm0U8hEpAB1gJo6X8vlQIJB8u1/Yjyci0ALUOkTT1WhVvl0uYzSx/cqOY
cwzSSF09DwQbNobJGM8w2hWatWr2IHhIP5aHk9d3JhkUUbFS/SV06EVKvh340CDd
kqg4Xtv3G8F5dbQudM6ianNERsiz4mz4MMpBRT7vJZF35r3gLLt9/j+NHQh8CIxs
NwhvN3LhWe7g7bxRhWShL970wWbI+4p1bw1sUBjLyMr76/7W/jzEZXVOz5DsHJ5q
JxWW2lfTsQzcPwLI9gZxm71j8XoMZSTUY6mIUt6xzsBZ6+CnFjIFZ4fFrbz06tI3
ObJN4Ujr576kbvhZshaRc/S1WeaalQi/Q1HpdauO2Jkb/SGX14U1Z97fpOAhUNsP
91y4M7mij0dFbhDgzCCkHSpZLryFJcAa3tjSWO3QIwWNhIWwlU30cl6s49/+HCaj
Fl6lkD+HAJ62sHI0bxB0Kzj9kJFcPXm7RN+5Re8c3F13BSfZMiBlIPov566/PmX9
k5FonsN9fxcN692N6RJjLBo+eV+wKrky0sszj1XXCtdgIaTD5egakWfXjFHcWWXs
d+uYeW8MlLcVJVzE/VWwdx7WycDrFxgZ0NJni4G+b4AZWcXOLgVQxv/YSN+R7qVa
KnVmG/ihxYpYFVlH7Jm6ld0/rcMSkE4rqfoX/20UtGCM9PYWXEbujD6PmmJeCd1z
TwRT4Jfcdth+w/g1J3JHARl+S+t7ARXW/EKVWjAAwgmIPrWPyqoH4vB7HHWAKDla
7XAPmqPsNpqURBjCw+1V2GCN2mp02zFABa+jNvtdx/aea3eKW5cZ6i53s8PhBGlD
t7RAV/GsrWFdG45AmsPsNaJ2xq0a6GJs8zPbLpyy6WhBavnAIFzTePHdc3irqKKP
dMQxTbaLqJoT4ITFLQPI3kiO1CaHsUE5qEPhO5NSlhEwyqrOKqt5FugkR1XKwpDp
j/Weu5llKm1Q6h5Tq7lMf6ntusvDex94sP7Jnn5lG2SNJbTWdDEeM0Audkz1YdO+
cC+eWMi6RGUvfxzzYEpREi+mgkajbJR3R9D7EV2h+XsbDL6pyGb1SN826LuQIMsH
JHdO3f0X1qpCpYtRSx1XWMFsEn+SyIIuCJcYwffm4PXfgHSYJ0a4/bqGlTpn+W8u
e1m9dfEH24jDDZZvwqPHHU5Ypa4O4Uvae77vA5asqfpPXFUw4ESyf2MlsrFn97Gr
2XfbJwv9nm6VXPLgsGU0oqQLz/PV5sGsvqWIHs/dk6OFSDEeMuGQcxly15LGoHai
8/eoT7Isp+OpuVi4voxvFhEdUrOxzMpMMSVwhjMxZl8zJFkeTYg9TvG1kYHW9LFd
xys8KQpTlN9+p6PklSiAyb/6HKSSw92ly4kO/tv+jNu0GDxvjHVdlRv0eiZoi9kx
1apus+ePbPeo2Ra595+E7wVDSusmIe2r59YxUoRKoMQU73x7cLfJ7C1oqSRkRRVi
YTIdBhUgE1Ila8kMUPJhqgk5WsbCfftcUsTrnDjZLJrwmdUU5icZIAbIpLcf8vVC
xr/NGRX7E+DlHWAZVZ5Uzyu1f5Cwj8OnUxsQcxREZEiHQ5KFb6XwRplsHMKXOmXV
/uqGBhGgoPVH4KlLAy1WwIxz0C10rfFWBXYvVKf8xyOvdr0Qrn4hzlecbJeXtpY+
pyWhery+ZT2LBOD0sDYe56DxRUT7yos9aecsIhiMEpXlS8YRY3DwrDCQwzzMK88q
u0/QGEzozjxNKeq5coeuMfX5LxhQTNhdLI02BVpPcvDBZO7DmpK0PWVoU3xFhs++
q4fh80gJAvUm9MYSyPfkU0LC5WWaE6drM337n1LzPxlBaxbhxGA6ALycpRs3+jtA
oUmgKixIuPCtqCMdrlmm1FJ4e2HKl/AJGoW2/0KjQykSQsJPqHhu/uB6OA/2ye3t
5EZ49qj91u8RuZuqNb62BY1TAScHx0UBgkizoHQoDBe5NrjIpeAXpN9gVtRl1ith
vmIT3gMeCXObJEl1cKoUNsfVCP2waoEo2DV6qu7IjPU8bijca+9oYpTtu6UPc3Rx
4KvDafIAiBIocym5E6tixPBZ2WaDALeOC+AXvi1DYP3ps/OUdpEyj/DetBrEyle9
r/azYoZvNq8mjCqwD7trM1V6YSHSKd6/nri0qCCv9TYj9/LAKVHfibk+f60O92DG
c3iGULfqg9VLW7uuB4OkSS9NKxmKiLOIYM86dAVq2CRc1zukdxFCIHaX9qMvUc51
N1pBY6I7djwiduFlgyrGdgblI6Ityo35l13wlMN+mt5gV5GdfSEqB30WmhevXJd4
S2P2/er6sUjdVe00/LfrqgWlBKQeNig4WWUq9HHTN+2mtrtBOTlZj8gfMO6O/cFG
64wvDJZ9jlw6HlWXvQfUP4yufhlVf/qIW7Gav2FmJx3CWRr4XAGegrlK0UR0lUtl
4sbhzCPSZ/Irzn5E+dS6qD6qrttPpNv/kiwDm4VYOfuhZqjJ4okopAGGbbPeRiux
Nzp+O+zz1NEpXLSQjBD6OXpz9sN8LSqAt0Dou1Wlq+ub33uDUTNwMaohGO7AscYf
4wj1UrV+2xzMA+uty/7B1gDy+h8zDm1YjLq6O+dyn4TcEQbSCmaJK6a7n6Kl4h0F
d9seV2SqpEgy2zCkR862ETisFguQzHTZxFm7J6UVUqh8yuCsGLwevgwjJIihACWB
6QPVr0n6YLME2fpSpt6rJyJxkgl3HwfUs05G6KbcjCJq1oLfqRPhSiX6qkFeG5Cg
k7eTPoJetRWqVIQzlO/Si7LSLKfGZ1099E7RmSQE2B7chAFBvjQ7Ia2NhLKbUB1p
AQ9NV/auE7KMiGAZaRPKfzgl8VD02uWe0Do09gda9EzjU6giqWdgzGWNq44d9cF8
yVma6vImkbw0MD2/4IpxW/mCi4NE2C2JZ41cpK/r2Bj6vVCiILAXjQZQV4/5UYvf
aSOxw+FWd4aYiRZ7fRn+zEC36Fbmiz6y6smwt98asYaP28dbAl6QUUp32gdb1c7T
307QLcFj/ZURtxli04EwXvqxmBnMu140YFvuzb1o/2NNpmTFmWrJKL0HUgJSFEjv
7tWBac2LQWJPOwE9VheaAF4rhlU47p+ZZ7LK9Sf7g7nIUJzcb3SVIffYQcBbNmIE
hE2Aj6VQeo8BhfvQYlqTBJGK0G8yEaevEJmVCfpOtU1akcMHzdRz3/FN/KnF3G7q
MzCqHexLABp58fYJlDmDoD0iQdFiV6OXJCfyW6U5wB1IGrC979dyCkdvXBRTmz92
/Qmn/T6gYxaswRURo6aOfXkwXATouI5J7cp18LZUquBCzK7Qn2PW1BE0Tm5gQ4kr
FkwxCY8ZhNFM1kq54PDsjZa+ZLD49rSQPu8VlfJKiEnPyV4wrQtUUsAx7QOIneSE
N9vd2HJGow0OOn+qsTmkrmPnotMz32hhYHlhSoGIwE0AMAwMgK1ZvJN2EkvdVpac
TXjl58Lm1+mZJJZ1WDiMF9PwP+SQBgRy1yKBMHt/X+/wbaBS+bF8vjmzptyxiW4R
NjGr/zYAz+Z6DS81LyIfvocxbfQ3HcOq0c65TrcmgrDZHYJ3kOZsoAuTrF4Qhtaa
291R8YmFPHe0MUrr4qQKOUpCzMv6dQwP3Goge3sNrvtUVIHsoLBejAramH+DuGma
eQUgR0wyfmFsrUYymT/sDen7sZBgXhCu8lZVicYKAHV+ziCqzvDMJD4RTt9v+I3l
Hfmv0K+oCHT2vBw8u9/ZSdYAsakqByexPLXT8NKTUQ3KGFjf0EZuduWP5XodUsXV
WSN1F6Vu6MWAOX2v3flH1GppX5szrw51OPymFuaK+115vdH2Rm4Tx2EiHlFd8NM7
/2q+1Zj87n8rxMEXLfwpa64B97Q8ofh3hd6Pqk3CRcgMKUsndpaRUGWmTVkvTHbM
JLH048lTpqF64hg/jFtjgifz7e+MgAATnRe2Bt2xCyFU8qmSxpic3zrfnOuGL4W/
b92ZugxbXopB6RkcoMq1WC1pYAZj9MPrUMlKc0rhCptHr6pu5pQ9P1aXxc0bNKfs
y0yQL+0EBjX33sUP1KZFWBGdGkKkGVRQ+iBI/j7X1pYYuJD1YTfYK+TMLsn+zwLV
s+4NG/X4p7yT1Z8xyXf6jEsNcGP43q85WSjZ2a9dj2lulCp+HKk3/0b4z+Nr8GfQ
OKOhWHKkVs5bHt+pYjd8uYSLm55h2DNLhJubMuDtd3BH9KUrinS8ztZUBVxHhCul
S15JNybCni1L9uuFa7/xkUJZ5zT/Xn5Z0HF5gGPZKmV8nG1XUTTdPMU3sBSazEgN
rM/tmf9l1cNB2869+zVLBsCCQ/g8NraXJyMo+JHpaDAOs0XOhBVVgR0C+TJ0Uid9
IhO4nH7HLg5bq3V6QlC3/ISqgzgfEHj/tcn1QER3UizgZ2arehpv4dZaPj09vMgK
bLPQcTruvfjEP6WbOYgLbL3lRdn/LDG5BXx9VtxOS6Yj8MYcr5uCazeoZShnvDIB
bJ2sLh6/lBubyrUvVCTIEdu45tFTFIsfPu4NB7FXGjKqOzAIc8+QN2SafQVOS6Pd
JGMM6Vetqnlu25SLZDI+lvl2SiKfYpYLHMDCPkaPhdSpMNQQnLxVM6F26K/Un04d
YsKLeMC8yff1F4TVxHcuiC6czbIbl5H05PWN9u7aiecNOUXBwqRlDlxgxQJXVgrw
0n8yd4wD+PgWGnF+2F2IU7ca3GbHv3aUzP+zdXGbqXUbylOhK9JKatPE7OgpwszD
tmfxFozfHODKjsUE6DdVpBk4nNQoXt7/HYo/IejZuNaTLaFOxbLPBde3UQi9dqVV
63t1tPr0WCo51Fj+Gbc/cKiY+jAZEP3z0TdksrUri8X3CjtNzgjkZ7SjOkYwfO5N
CQTBrTkRLZBQorXVKJFBIiygmz9tU9NMmISZ8jHzYVpuWd557Db7apnyOGniJvW/
8RKwRQ83QdsHHxDUjkJWt6DJVznIZeXH52/OLGs+8abUsFgDKNXcCbRfP+XDN5rE
oXT7GnlGgYYhyzJLVfJv29hT1LJ30uW1yT+mIGRsvOVAnINRcfC89sNfo1SgHIxH
x8oubDXBQRzJ61muK1qq5DIjiUBqXSS72argqi0E7DO5FezGabEJTlpYtplUGxp7
qircgZOq5833atlK59DzKLB0II/Mq5sRV0wgKAyV4tt6qq6Lp3Rr4/WpC5VumB7F
4aG+7IjBSny61fqn0lrhIUdnBsWsxRAODC8BRVSKGqL80WPo3C4oeolIgz9kISbu
LOjT/G1LQTaYQTlI069KiySNLYDk2JxBq4Su2KjoYRcH+sw3AcXq0tyHTHK8fEmg
V6Y9ZwMF27P9+fikefYyTHCgXqN8HuIOi+sUUd0wnCiXq7dKc1Oj57Ful0mXasEf
KYHOUsmiGEA7JHEpXuIC1LQSr65jSUvT7GR38Ydr+LoJvMkIu6UMwbRX19mD0Sdv
lKNnSIg+nwl3qC3bDp7UekCDVELeWTN+3rvqFyhQCaDluY9HYplHPODNq72ZHsft
uJnFEr1aDfVMWBPstOKE3RuuwCpVFTpArmJXOcbdhv4aaNgbPrE7FxX3Z6BUR5Xc
i3nhs4oTZ/VNCf/izC3+Ef3/9dn8iyI54B2TmljsEMlKf3BAbhLolCdERb0aAx7k
ZxeHmstFHN7FG+ZMW5tHmhVHo+BsHCMZMHr+klGCBEsSAB8GCx9uwcOgq0/Ssdet
/EXVMJSpqxfFwpKu4euaI8q2SLPUHk6Q2aC6Uwtt0PpyIVSK6Mf//kbMAeOd+GD5
CdVrg89nkd3lFZOyZSjn1umWqxtCqVOsVnak36+eglwqU23Rp780n3CLFQpiP03m
8CFzg5ehkpV0IkX0RuxgamZLCHPYwnEUe+gWgd38zmA4/jhJY0W6LLDF4eA26cMi
CSOhvfBtLTHvCXn28MrZ8sH6afIK2xMPxjAo71sIYZ8b0Ci968+5eucs/DxnLQYb
+6RPuUrVW8CljlRgQ9htOf59aAqRZf4ekeLWWH5Uk1RNVNAaoUV9BqZlMDYPkgWi
Yutey6jJlPSRGWYFQGRxkgtS2oj+Wd1SommOnc5Y8Yjeyz8sd5a1xlz/BYGFc2xt
O/fJeoO23MWMjdajBTsXOBMd3kdtxwHsMJ2bB4bb9jVOK2Lwt/fxrgT/I2JPD8tJ
M3fij5zTPzNRUiGlnsxDx88uB/lZw5sKazQ8D/BVq6yuCmZfTAlIej3TgxzyOCHk
BtEopdhGOgluwFd8doCI5ymfdL7ibKvFqycf9tIpivusNE+Xua1JZvhqbw2Gp2Xo
z3qjZp2zXHF1QlFyvUv2YhZCQmv+zBTHRv/nSpkAvv6Pe3MUKNkApG4kZbtsuCeS
hjZKOvvXEiqz1+uOTP4HdwC0LwutIZfhEDxyqwj6XkvvTLBVCMOvqmEBKRz4j727
uzXErePrfdT08sFo9ziPFHhG+x/iftnYR6wSlJtpgJFHPoGpjur76imj3e0swtN5
f9RDGqF9bRm51t26PU9MXzyjHOfIv5IHyZ/XHlpr7NZ4hFFLRGgdFnK843lz++Rd
awBystOwmdbZkEzZ2PD9DK7ZsqTgk1bAFU67zcLviVmjNhJ6UP1jm4ab2KwLn4IA
nhNcYtgK56uWVNg+N6yWYxx9Q4vlzFOdqcRHIdhjFKhIb+omqHLzZnioh71E50RW
31yFdi/NwbQodFKeV3c3yvveEp8UhTpYeR6zJK0ZaXTuO2wbX+03KrhwudGrblR+
iQn9mCY81EYNqHJp/7sD9Ro6z3ucr9C7eJGnxBrem4i5w0MuWxfW+FJfP4liJkuf
6iptqboor7B878fn/NEjRczH+Fv5gkToP9zlnBX7buFohenneRuld/S2EcsQ+wor
XeeemzwktDmT1eztrhF4tYdWEU87wnG9Gw/jyNfSnkRsIx8sGa5AabfGgG/uUx4x
uNpnZJGtqvWscwUiRSvKJ/PyvGpDtri46jvM3ZVB2+R41yD4t71h+1iRWABh4i3W
Og9uh4ful1+uYrfa3F0yQhn0wuM3S9AIlpO87HQhSDHQBjMASO6geWOje026Ecrw
ajwztRJLQoZjRIhohI3x2saJLpUpPGD253Vj/3I62RkIOqh82E2Iv6yLuoPvi8vM
0MGbWL+9UMZRgq8pJCQRkX5Lf8xFyz9DevLNhdakbAYPKjT45+TBFuGnuWM8l57f
yQd4dQWd2MqRfUxnlWgUkio849yZWtnCGE8fpzPGkF91rXtM2TxLrFx8EMVR/TWT
Kj4wOVUOGEpNCbNHiEFQEwC+uJqfIeuGCFMiqy/7ubn4VxfVVAUdQjy43qdG59TB
+6DAmINpL71ZC2QPL8H6ed/YBhIxgRqzUpM6zHjtQHgAWvSnSsZKSfPioZoSVc93
tmL0WZsULyyBKLAR5Wi6wNwzhiNLjAJtJzRjq3fDcTDm+bWWkH/0FuPYh2FjSmYA
h08xYT9YquOV2Rx0w9l6DSuY7rm+zXWwobAvMhm11GDVXD+gJvYaFEZiuOgYrsSL
ctaMVQpDQ82qFyEzO0adBqj0ib1FF8OT80yfHQgVGw6wX2VtqTbiVtncvhC4snT8
DbJ6c4iP6orok5kkO80TlFvl/dwwbdNkhF6z97aYC1ZJml4/g+V+G+BZYKvzzVBH
LSIM5hHXA+M09mkWqYUdslBerPgS20IOyLFtTiqejgufKrgrDaVzHxr5keH0AF3o
+RbwpWOJk8bfzjGwT7/3Re9cym27lQYWPiZp/UCWRF1wtT19ycZX5jXArBoc3aVY
/FMs6aqqPeNAZnXCNVslop3N1jt060kgr0cn7smEsEXf+/nZDh0y0tYT2mzQ98ep
8fcv4VMcn6KrQj4a8fTLlvsOpwh3m6/ghGnmnSfYK2hGUgijyLr8XZFu3/Sg2nkY
KdesEzbuSgifahSGGGlxVqOTP1c4bE1jci5gwCOZZe0+uV0OjZHLbWFwk85yFrd/
UvH6L52DAsb1Oq8T2dNzuUnlFxCqrwOpMXuUY/MwReURrbCbaZwzfPUuMAGoOpeH
bp8cjXtTXVFzAxg6dceEun6deel60diIEEW73/WvAk2V5L9tI7QX66DAQLUB++jp
SM5r7OPR/g6NZGOZgVBw3UV8H8cIXs5ic2o0G20I4iok+xUZQ0keJh5c57Wzugl+
yfDt30MybDl1YoCHn8yVsgYabFITwhpFR1PKP5foIS9KkXtY1pLUyJrtPSDRdmlz
hzRyn7efBjPYMpWT3ckPX1wuBXJtHR8/kz+kpKQJfRM4Tn5G/9F2e5iEY27tUGXw
KavbJQPW1Xw4wjUF/UbJtK40WPAo24tVI6w2X3sjenhe986swaL/o1H/nsLcgS60
N2rfnab+IDDwQqSJUmCUgWHyY8NG/XJD51CFv3RURc/zT8+DTPMUn0ekiWFj+nYB
AFFr3bpG8WAl7gkuIU5dOMzplouMiZIPW2bCEsB+SYiZ6VOKcc6hW6f50QqlhJDx
FcsmytvIYm9TiJsp10//+vL+JWoMj1QLPH4pK/+0J+8DW+qi6CvX7ESMXffgZ4uP
qA3hd66bVFCGeO0NTeKwU2AA78AJIwhegNPyZ2w9UQzwlzmIzKHLFC7QSitUf7Op
60Lrm2y5KLtR5mifcGxsMZR4LkOLxRUgTO8oG4N3DS65hUynrowpbMQY+vzXLg8R
f7rjx0pcDMrR1hJcAnNd0YFZFYT2YzqSWz9ByMOoh8EY8ZarZrLUzDeNUKB/Bs+X
PHe/9IF3+mr5RJxwMuajf8PkdL5preYtvByFMWU0SKZDTEfCyd7JpR1Tk5GFuzle
6dHqxw2GxwOlU2cEFjkW8s0CRNYPujaa4+Vq1O/RwmXpoDs2ly1SYE2bylgOJQvM
EGFc+u4//MoZNUp9nFRTRYLVT7wy02igeL+e9h9uVGfN1twcDaGcEZPQYV0XFZS8
RvQfVVS6CcoBAC+UBY17K67S3Sjg/b2aFhupeIe/8OP6XDkVjECUyFO0kpFw1n+l
QGqu69C95Ct/1itoGXmugk2xonsb1DvXIXQqnaur4JdFwo7RY0Mt9QPz2CdOmHx/
LprWm6sxnWX/6LGyykL+bgShOk6OGVdgH2257RxKDyp5j8LIGz/3WbZhJHuf1pVH
Nr8kg4GhGB9GUnF6an2PjtUkx0jITNmDZE0amz+cuwb5r0l2YW2RSJ44atH0KFcT
Jad/y8T+meL+UqRI/xNAsOY9gfSk7zsNCv3BHZxYYjE4djULwbcw2dYbCiriEO8S
FUc0w/rv7mItPLPgrfNpa1xatvy3FFi79Y4UmKa9O3zhMua3j8UV+bkhbQfn/eMB
HgRnsUSCiprxM8bGeJ8wIthcFQiF2itM3B6P6rwkgZVa7dkQn8DsFqHD/lZ4aacN
FTagY2654I4Z7E58seZKdIOfpPAQXzgJii94itm3eo+koukpAfwxdyVpSt3H+hYM
fZNkDEhOUbqKnFwKCtpYPgUA4grvR8GJJXUpPdJn3/F2PF2/r8ikLJ7u2xyBJZgn
3YA7vHoAjE+/CBplC646e5psXNcJWDrLOS66t75PuVFp474tlX2iZmNMreall7za
NT30cddqQ7V0AhHsHGKER8Ji2WWYYsVYuFKYWQhVx+d6VdN5sXGH8MenDqyy66hR
ZXsCmgOb0FrZJ2HGqjF6Qii7dsdG0+K4Mzy+mwLTuECMQMqnrfdCyrqTE3El7Uj5
23Ff2yOgMy2Mck7d89peZyV2Gx9VAjt34sin2fjEjypg2QZrDq0N34/gixVT+oCa
7RFCsUA9AiovErttFLqYiL9q6KJckwcfxXxp3FH0le9sFPhoLlyjZaSvWksFDSr8
zGApaIyqSpwxzQyftJ4E7fsX9KRdRoCHz0/MBbNEvHTGnS0lFQtqWlDkVPiSxbW+
FtW4ri8cfyP9cl2Ynnbe29eer3/+A6GFQqyqcsvV46mksNTF8d4ZwmzIFviOr3OY
t/edddoQ4o1dhZm6Ccj6FQDT62MvFH6WmizA5zfjGy2IX5K5s7topf7G1uxQbpkM
XPUOoZuoRb0URgh6mgoK1qomFzdYDzPTnu75XOdg1+GZDz5R+AuhokWw3E2dYhWm
pFLKBV9ZaPgLJ3bh1o05LVA5y72OngARZ2oTHufI55nfSbQf4k3fvScdRPhSDxJg
Z66Rw/UwT3/cYjpmHRKM83rH/Ia5GPstSj9EMooj6iFUNBqKYTR0F7nG3ycLJoDu
kStCt8on/q5RExy21+tV38KBy5ePlyQerNBlOB+jcJEssSdk3KHXdRBcxaBOuuJh
Wrxj0tXJXGoHc+qOJdl8hLQLYceSmVMey2l+lGXrHT/J8EY3SM6x8XEGYlJI4A9f
DC/cpIufsQgOCmNwW/i++Djc2UWJCP/SNLPKZ1uUeA9tS54Cny0iIb6UXyG2Vymw
o6GxovXex5GR7TbyleiEUISjLVwhynNN0Ta9gDhvPxWvVOlA7f0nI0k9ocwUL53R
R8t0m+uDSgnqVz1ZYWtjU7ALHb/Lh4yD20KdfV+OreaLkRDfLEmYmuCimdF8O+ko
OMfyHs0GE9JxAUFaVZ68gnynWpdnriHhDYC9F6aRGIXey6PDt6MwVcLoLMuEAhnc
PDY5CwWdK1ft+6fARdC/BoWNxqoRE8sSsqazkclszQ9jYf0kZHadec0t1ZLItjCQ
+t+O5c0GcQf/5X4/czMQUVDjidcb4c2jzQRbXLM7cYq8nnwfUcttV9czbbSCfxBT
UOraVNBrDU3ecftM+ZVa7seZgazf9ftTrJfvDGMaExldFXAdvwVp6RUwBXact403
qaJKzwxgh5tMU867ADp3LICjdMfHB4p32dsTrH9UYXsAN8iRmwk1GdIsQjf9N0Wi
RPB3TP/iDVN+vOK8GxE/FFLJZyHOi1MaPeULCkOVPVXbZBEETCoOd/c41cH70ILX
CFH2CPoVGVbY9ccv4i1xCvckgZi4rhnOzvIHOTlO8bWjvJgpOU4KCywt9FOsZWGU
EHMbVgkSJUA6nzQQEt6R/PNAttM4ThO+vATpFjyYSwM++pq+yBL8H3ru2uYI58ww
GnCyLDw0nxNGHnP//Kuf1ORZYum104kB+v9UlyfUlJ28JQQSk5X7wwwl40d7fhRZ
kKFWxZ/XBGUpZcdRm0AC8hwV5kPVBFEjJzsDS7EaZ9FfDBzlBGF0Mj71V6RrT56c
cMK8u7Xk0m3MF5P6UyZoLIWA1765bx/mWHu0UAB94IoPxwJnR5n0P/lYeLglsoI/
+7uB1R/e77VZOEVnbSrxRxKad1Ep6q7ji74tRLYfYc6hIgqL30akuhy+rxOHk+jE
8I7r+TMuSIN54IwirtlG4ko9r2MQnzITeNUZc4DHVvie8FV2q57NsNUCh2hjQMBJ
64M9Gr6+ykYoRvROiTNBAMbHwUTDVpXzUQn6TDIeTkgMWiAPMkXLcWhd65q3U/s8
1Lk39S+UQVsnmGYihVl7ea8XvesNygcF4NaRy5g7PNWCQsJ1dLnGVOnLWZJyx8lz
yjsTIqMIVBhEHoCzYx8sVszZRRaXHUlBqbXVAbCf1z+OD8bd6Jmu8JOgWxiiKxSq
u4/T6t2NQ2wLQ+mAaQs9uh7CR9cY+D3TXav0zGvAqdjUxoa5UsPRrDCXnuu0zApz
miOHCLSNolLLTxNP3y1QwmbhDtI9s1vkXxpawVicRAnK1wXglAsC5W1BF29wxD6S
QSBgaWlAq/w2PqKpeTONDYMLrc/hSASTu2p0qi1nLTT68AZzR/MRsWq0vz73uMZb
VzaoZXWY9AqO67+iQKu/QHbB17r8uGTrZgMykqI7wGwKWDa+EEdcFtWOpR1Ug+4Z
YoQIjw1U0sg5qgjykpV8nlaHw1fqPv2mOO09e987Ox5zXa4geYOzELPHVxaRmzGF
QdplqXDuntdqenbRDSb3MaoXukJBVkqXg+qdjHAU/WqD28g2tOhMFFPvHLRJ8bX6
DQAXvf7myaJM2bD9l66jYIyZ/xJG7mnlgFxxaWIIeyUFUzfR46bAaRhwxvsPzYrz
dUEdcQdpJQ7wAaKpo546LjS+u/F92EA09CxJIbhFVqoHPhCB4nhXD8/1M7yvW2Tl
Ymnm3Y6Zc0W8RVeDccf1lgkLfTjwgAjBIJCNHIyS+oCI7qgeHGcVwlxerjMDT2Vp
FbxZzdxbrGwHDlJQMUYvMeV7Y31wzb8GW7N+Vv6fCJFtCKSbJPgfSvvLGmcWITxF
vsJtF/emAY04j7ta+eV8J8yMmfRffmfESMaTO87wCaZa0fQH9WEkWNRZID2F3oPn
7a88xDYPFrUCbt7mhxh4PtUQ/GiGaT8DkUKpn2N3l7n4FWi0j3FmCzRG94yUmo/F
K0W0rJMgTIZdBHQoO3jsLZiQQOiMvTEk/6NyMK1MpmGA7TBuIbnS6eWiBpJRqW8A
EpFa57hI8s9mc5Bh6RdTKw==
`protect END_PROTECTED
