`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
MHFdF8qAxoP5KqWrdukTHRr7a0oWCpImU67rOyeV4MACPAew9mDjujSy1FsdC7lX
5EqUyUja2oUS9f4mwf1GrlJ5CVhbff/pbibKj9INMkjrDhgEnFBztm07Z56BJtzN
fGx57XbPtU+Sq42g9c8GFa339dsxkFI9zsjWqLcCt7T4BZZbmcAS+MaWBiZiMETc
lGi8VNC4yyhsi8jMqIyzJrUAxwJTtehdLwRy205u8DVzUh/DIndIi7bUGW7d/9W4
/8vsnrrW0Mz6KapgtUSfOhC5Ov0s1ar9IgeLMHqgJNjmSmEzZqXS8ppldzKgVu/N
rqM4/7y05tf6epcKlUg8LDbQPAcG3lYqrzsqvd3mCQ/JDyuX4QokOGZeLeMdUtju
hhxEFQB+trbQ6Ci6lIXABZWo6evs+sav+4VU3ZNON6iNSa3FH32f4yUd7XoglUIk
F0TKl1fcVuxwTPGqYALZq6BwMS2AjbRw+z/q9wBjK9DBcowLmy5oQ6FL1QXY8azH
VmiVdfUnjE0SdJfT9XZxCChjnASeL9zkxBVgXxGH4uMffkrMDipv/oeC241r+RUZ
a1SSVI9iFkMlbKwPkx0K/mmOL6ovmY5+xMphSWDyn1V9z5WEvEgmWLQ96pel3adt
ahpH04k+34ccYatbUaqgbJG9WxTaXynR04vu3ECAV39afJ3VS8n2yofJUGWri5/m
u83rTVvOltkpZJsqiYY2qAa+jJ/8+js20gChgNei9mMBlLiNKZic9amCwtl4bp+t
OZYRJ03SuFki4BhnpB0Y45iViloKcdsA/fE4YaiI8/1ufvtuIYjdS9kTB/bcE2Yu
IU2D7P3R9vNk9bYuw6PWsFAkTwlY2yd/fT/OWjAfmepw9Ti3PpmCO71fFDdw51sX
7XoHuG2tXrGxPC62yVNux++IZhh4m0rGtOwRQfMeuB2E6k3mbzZgjwiOj22nfg4B
u3TYz78Ig44/Wd1prRumVOS5CtUaCD1Kt/aOF57HuJ4HNN/LFNLNQr4AonsBPybx
FM57FRaXdmDGWSNFr05HhSh73KzRTaD6KMxAG2A2RY+OVEIpo+VNUhFNVfF/4k8P
SHjVBfx1E9WO9H3RPXnHulcWpEi9cFtLgT1+rSH2DO9fLOEFs73m2pXjWiKCWJT0
6x/Qkt8Qfz0kGq9t0TvJ+M6NTN/dngJcdh0iFDNUuaT16pgkTR78yklXMmUFv60z
uCfKtw2Ma4HQy8N5Bi1qqExCTxEqTdDlOSykRzpq185bMZkG/x24XV2PNJ9zaX64
VRW2XHGKq0rVfB5x28I17Yv8fvneXAh9UXEawoonyFboV80GcKLbbRoQyC4M5v+t
ypx6ErvFw8G0fxBUDrErlPPUrKHZy6diRccl69il17Li4lwbl0xwMBuv4cv2dC5c
cR6cLdA4/KN9KTyzS4Ya5Hge0C0EVB1HPp+lEenS1NgTvqAxFldPahHcigHQbFLG
APWlzOB6QCwTrG6uEO/49dnN3DsIjEosUG3QdW4IpvDHifFXD5qFjfUQTjKTkkxb
lw2QYZ8T10dS3TWlz4jLuAFJKrS/x5/xaGX/v//SnBU=
`protect END_PROTECTED
