`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dKsKiQg3gMFncEQhWsWjIqFouZMdCdV9qkWbhSykq4PrM9RyMNT3QvbZV/CrtgpG
X3I8YknoRoN6Jq863YLLJWOyCY69Mm3WlhzwYKgRVWlgMcPNuOhLrEq7kCaQp2WM
YILE0rcUONe1bCUcdTUVs8ngsSNZv6XU8JpzDFjDAg0uojWIH18U5YydD9FAQ8QH
zv/jHWbasAUtXz4WsHTMoZ5QBDthLm6PmqADVk6qjrYmDdd3RZp2eF109/AkRF1L
usl3HmoT4NZJ0FV4TnrWqvhoDy42f8lXUOkJRkzaVIkVQHkZdhJVLwXH94Jb0Q7v
OnOgjnNL7Sxbl1TeZ7a3qU/xnxV7PjVrk/VkAnfnpr65TtneRUCNEmMIiXo1SXCm
N1CW4Mf3ygEzhY1HPQwk4LOmZjxVbZcJD3xKjeHVWF8VGCxUJxJL8QQ7rFfi2LCt
Cq59JJEnROkGmt1uC2/SAkwx0bUeFD/fTEvpIl+Ve2sR59umEkNCSMNUZwQQ262+
S0ZHkugFKF3jqg35/2ljeNs0c5fVA7AppYokZ5a2D2FpUmiwc07W/HDzodlb/QRC
v9JwA3T7laIpnRKLNei3/JGLuyHHYmE4BxkRrtrhO+xtIrP+wM2HJIiDWlXrnYWB
/4Ql3f+uAVHYzL/8yDboehRQIEQKfWiNFJsOaXaYPXQ8dcnI2kkvdSWJ0+uSB4Hi
jJmWXgDjpYI6ZJg+/V0ECS6vqAJIPz++8qVvUdXzymK8yzjh4xQ1F6H1kpDQooF/
Tv9vd4JXZL09pzuALszaz4H1xgyh/xBT4m2C0Krzx9u4H+m+dcZbQFB3FWvXa189
zy3jcCYIA/jbUiC0RyL34MGZILVYM5fJZDP5N1bM2qU=
`protect END_PROTECTED
