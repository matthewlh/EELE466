`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
4e2Mx4O59WmH4EPt1V95kjLw+X1eGjb4hmj7HRN0HKk3a0Xl8195HcltNSvaKn2a
5pXO7PR4r7477KptjWckNLUjY2kv2l2husk7zA0jR/jN0jrnwJ6FwcgYb1lC2hXH
HX9UEktEekG9cqIHIk8SVhEtwPHKRKiZbOI7XdXNuDkWftU4Nt4F5g/NnLmTIKyH
lZ5hlvHB3ZwKfvFMkGPmRh/SiLo9KlO6Y95Hz2ftt8jnZKTgeQ4HhRfrYKYhKpaC
QZ6BgPCEVNp59uZF6pwT06eYsqXCNvq3S0lJNJ19+YTRkeCbNbVk+ZuMOjkUtM3H
yMHYmzZAyU7GJVmHk4SOIR54d+JOYOJ0yH5+2FSzQ8Vr9UIckmgIQ/jfkU19Pcwf
puhSdkVEktAQMA0QZzWT2epQMuOB90pyISnZJWijOJNk8nQ1SCEkXsno1B3P0WAH
51mwTg1QIfCvWkp2lKrXK2elOf1XBQEYomGXE4XUXStRAUryhUuO54bf4qy5RYuD
hH8Fhu3uus6pBiNcYf+VRIqO6+M0odITfskssXG1k2xD3VHHh2O3bWto0ekSXp2Q
rnelbNc0DR3h/thn1DiZnm+TYk6d+8ute/A5j4j2dMcwtbUwIY+WBcILlcoC9P2a
1XW4+QFw+QcqrokBVlszSVZ5gpzETgSp8gDqaZqYjmF8XQjIpclbwHzzY/zG6ToH
x4ejl4zZ2onC7VnSODpApdtJkPx4j7ShaVzeGJthZYJ0UwgeenV8wSizN1v2jQ/B
4aCICk+UitZ2aAmOOZO/zhLcgavFEpfhvW6RaPknA81d9W14einlwsv6cCFqxPwv
3N36WafO6BOIrgJo9ZOCuMwLrLqo2W3Dn/1a9tVmULlfmqMjzmde1nCmTHnq8Mji
A0QJDN5o8TQPmlIudFZCryMiFoBFmISn0NjVrBSF+SrE+o+maQwvGSsZvwax03kk
WyV7S22ywgHinEvLqfesBElIp/nAipti/8DRRWALxCnlzhOaWYd3jjxeYsDF3jdk
76tF8B2BrVb0tIk1+A2qQ5NUEzpWgRnT5512I30htzSKXStiduVxDMjSciwhbAZR
IcZ9iVPoZOWYkOtiKnV5tOmSIDECAcsaUTtdEowJ6Hpwov3Qqh3cC1PoNeh/UEc5
siXp03kDAcfjchzGzAjWtSScfRt+UsvOTEossreog9hxhsjtjCvQolZU+LNZWpTq
zl/+PVR2OmVyCdq0O2mc0znJPOo6S2W9Kpy1CDTSaTSz3g+iRtkPz3GhJ38rGSjr
iyOk6g34QZXktyqklg4Rl51Jbf//7Jpw8wyE9/00O+w23QFSjzEBjVdOfMLMTPAj
PgqQiB30Imuzsw83lMYYmuIv/aLRbQbmXH2YqlbhWS1+7kMkfBwabcItMdQIzhiZ
chaguYSNR8DmnDUTngR/u82LgG2xWXy1VXquqbA3b6I11vpP6pMw03/El2DE5b6I
osF/lDt3W/gwQPRGUlnwtdqAUSsNIg7cTZcpYg87N6/JtOC37j1hw18nyTCZ+3Jz
l4SiA61STBui7NjfZgCCrX+6pV1EQs76uzcFcElw7LcBABUrwRGU89jYcpDQPr1N
m1VbiOSZqp/HVoFlhtWbcrWW39H49qjk/obY9KDMZXck45ldzqZU9waFQFlqpMEJ
vHQxcmW9C0jZVtcB7XRCW9nGSY8t5nrJDwCkHydmYn3VL0L7J4ACOChOywiSwbiD
6iidu3dxAcXMv9KouDd+tr81Pe0hjpnpg1sHcroohcGxWLecRQzDRqPU3S3BeCGW
B8PsffN82hhmvIXH3KBsDOfvMcjG24UAxI14+OjTEsBHcYCcg1djNN4j3c0D+ekO
4uXYRp4ENpEZBPJyce9ZNXI8/dLJHROYhHEdVg+zQi9VQIdQYzBiU3B+yaprFJ0C
iH/cBVG9S9ZpPkmzlshuYocvmBpPMq3cGBPxCETVy4I+4Oyro7lX+V1vFY4BxgUN
8Ql13vVn2XNaBlwjLaM9NyuKTTjmwQOYenokI+jwwjUSK95L84Z576efAcHmMaAI
xF62s+dImJcUV0alXMArneIEKm3ZSL9AKa5sqnbIg7g26oWjNyzOrDkWdGJNEYTC
5FDNeElt9+eaBeYcTyUPLoFCrB+nd71sxBbvgyjgtLUyD8c/VhamzTmCeMQL6Z/f
wNeCElBGlM5gfBT1p7hgDw98IH3jC7f7BJ0N9GbIk4ICoWkzOQEqCTlNbTYEv3Sv
inHh4rn0PTzCOwGZ6uI7eS4Ovzrn77M1wvIfXAG7afQDzxLxr1ky1AnMf0q9ewxS
dfPRxKSCcSd7uXQGguy4YR0glVlsUpOZQ2onHnzvT1tlE2LZ2yZpGr6MOrMH6hhZ
Oln2QJqt+eth649Wbb9+lnIfWwIi9twrzN9NvFLwPNfpg2RO7Nei5nkipG0Mpnck
b2M2/DcgaQhy0qOdgvvuo3y0gyVpLquw7D+AtMSyQ9T5IMEARZdOpvjUeflgeLZ5
er6/EO80ivO8kZIKzzi2jv3gDQj1IEWd8NR1DtN/gEWNg+Sd0i1hC0ln4olRMjwx
oUSH33mTad6YlQWHfl3uyUO7NMmLz2DTgeBWOBmN+IcASLbejQi77IO88Dgmnri/
mUr5Y9K8s4D0uX6YGwkMQWkyCrVKl113ID4kI8DMA5IsfNytp01z6VxH6Hic9A1A
7wwCuCGqaqy5BrIhL759YYPmXCMh72rJBcuS/rKhcUmV+BAF4oaYuY6VuQDj7ptx
25Zqo6DcjKW08IjL6Z5WVGlmJ3670CNdbgUS3DIaJtspcKq1hpAp/MaHH5eFRRXi
5onkINKkHuo9ADib5hOtJN0J99xk/KXv8oGCeOGh5FJoZS9g+WqAjmDugem5Pt0Q
6zj1EyDjQe/0twDm1Z/zy6d/M7eGwr3538ZgOlCowraBMfDOJt39YtzVC03PxDq2
ijt6k2/B4QlzX8doSwEte7qP4PqWdYaVp0ssOZw8OdoMhgFgTgsVLaIqGGa14uZP
K/ecGJfRKgCki711kqVx2hTdrD7a0FtpoiUsh+O0PU034qIiikFRSfG9DlYICsYL
k46IcjokZwBqQP50UtxKX6ZeNTOr/xNUlxETpp/pYD5H33d1aLO2NgL2yMfwkjWC
UqcB0YnWDE+uQkcfBUQQzE6rh1zkJvint/LZxs6v/THlg6EK8uPvu8b0yDuhZC2X
jPlmLi+at3Mz+fkbYgy9MTZsynZDFaypt1sFv3V/ZPZlgezj1f7ryYlPbY1C4dFE
egG0Z3KrqSFGoBV7JDt0cWQRc3ECR/bY74jvYsoKymGnTu8EoLQxWV9KljymNj7E
JfhjXiBud2Lw2EzjFtMwr41DYEK9IArkhuYj4SHE/e0NZBB4A6kow7QSj0ZGmw+Q
/iIiyjiqM4j7tiUjxNDouv3rcWA/2jkXneEvAuZoNykNXwG2tg2cq8Wc38k9Ukvk
jFi+VXsOh9CCGg/Om8yMwv30JXeGiKiEkwFA17SEcmSi/b6gljlC2chsoCyHfwuc
GewessS7ieStyoAG4CCPzS7b5dAFdCISAsaVvy/vULPR8QA82VgLgXJ/2GZu1Jde
WeChonSAo6Y/S/2UAdeZ5mUOuwns/5cIvlx94lu/R81gfH3wGxqcmWRlXwkkJBwl
9QIsKaoihZ2jJjElI3rSVmOtg2hX3wafk7qpPpX2TS4e5yfB9MKoWjyMMPOLStlt
aUWOAviEY31OWxu8TvYEEuq8NWpefSPbyGGi2JnTVNXf0h9kV+Tyk+fGs1xWzwfq
gFLNsh28gvZvHX7XznQLy9B9da1ISICnhuEmf2upxfEIaR/PV+pua+OdvI9f2SdC
16p8YUUY7UK47t66W+ZB452hJslwHg7qu6tSH5RVvvLnO7kEIyqDS/VwAgUC9aKE
RrsX7N3frWq+H10SnREz79X7fHTxSYR+1yTP6uysgR7b7Ixk+/hOGzCrpI698DJ8
D6zBoJtwDDUVzgYl4iPNI2/SMnck8tAzh5dh/u9Yuo4AV9tr5G+yg8+oPF18TK8n
tk6O5wXTATNqvhKnM/TPJnU8XkJmkr5TF/BKrLiFHJu3/kzIAX8vIK8NmOEaJD4G
SkSRqgQkDjgZNTU9NpVquDn/Xw8iJW4RQ+9XE0yDHo/5hGNlLHht0ytUzrFFiPJl
F+zSaa7zhDhM+4zXVoAzlfenXq+qyyr998z3RuzYmXjb5RZJXwX3jKFumL3ETGYf
iPDQoCDq09s4qNIdkGYActPd3WRJidWwg3DwTg/GBWowYkM1dwUHM7KsxgdtNI31
X6yCcElsgPF919EoQSSmAsjrS6skEbWRZzq+bc2DprGNxjM9do8id9Ff4WM4ds5X
bytNZZnwr0PCsnhwHymcjQm4WvcJz2b2AYMQqcDB+v9hgDsUOdLt8XFEZbDGS8mT
BaMEjSLAh8uGS9S+Bib+Iwa7b94IwemldODYW4KgCs+8hr8ZrzDXgfh8NZ0QedCx
dt9pzFd+JpRJlyVGGZHO0427BmxHwvLVoRg8a7XhkAZAsCOGSjbDETPTrAq9WJbN
ylvrsjGWawzc6U1SSg+P0l/0nKNYCtSB7GF9taW8xktT4nh4GOz+7ALx9TUOci9N
GujWD/W/arDGR9Ep037LaExBkTT+1q/srQ4z5xxz1+PGOfon7LQVrO/J6bhz8Kau
o6Gcc0utm03/SVefCHkJYFtCA2e4ehLEkgoozktuib6xvfqMRGOYtuaeM/V72216
J44C7JgqDyGdI5mTKyz7Gu7jtkaoArTSD2DrhfIZvtul1740SydG59VRGg/zEvw5
Oq7aOBin0ptfXqGVvq2EwRljqELNPbeT1S/h983WsA2Zdj4EXWoLemZPn6ffpe10
bNVNJ9h0G0ddgj6LmYrGBlVbayusf2cnk673HHGOvZDSVbr0QczYs28kiB6Qg6kj
rb2rQB358YUb4O4uRHjwuKe2KA6/eGrktchSS4Y91kccr6b7sZ7oHnV9xUd1eqko
70jeJwPYEWRThk1mjTiJeQTN/8xV8hLJQqa0IrnZdXmYnVbRLgjH6woKYG6Z+TxQ
5cL3rIAsgoBV1Xv5v96vqyaiqhYCooMBaLL+PBU4f4s3DTqoH43qlbHfXZ2tRTxj
HNe019ZSdt9TZqxpWyaUyfuf/a17H6fGMOwRbjaqgDICGpl8LXb/CERPyfwQrJ+3
oTO0YckgiZqU51RUnyPrgh+W41bdxx4FrR0Ad8oOvG5raRnDragz8tbh2kwLPMWu
uZT7Gs90QksHjI2AQiv/yeE9JpouW1e4x1ZJOWzJSMN6oQtN1gx0AvZugqOMciY0
KoFx2mRjQ0+N7H30kNTtnW7CeDgZH2vDt1MS252mS82ZochSTp+drMuAOCy5jke0
2P4PBq6kO3rE+8SuZ6TS65Fw4Vd4tD1xeWcOsbkWHw1drsle81E0JnyCH3trFYiN
VXC/2TW+UuFRzJrArFRhSuHIHIrKvDHpUwMig4yDnpf6sng9iocJYoMRNkrz98cZ
VuPdiN0/cFMsExjGUfJJooLrLJKs6hVRcCNZYOVNEl3g2lWoePZS4oVTE4sdAWo4
lrK9VAtjEli2xr7PNGnLRbQk+N1VlJuaGjmMzagH+BboWK66qk/ep0HgnkPUDaMD
yL8fESJ1zmeIo8T7ivP5EeubCjCtXuPD65ysyPTZJO9pJO7CMPco0UXh30v//GrT
vCzX0kW3Tm1V11W4tnrSak2qxRplxXgtWzBdRfDEROhmTVkznX+viesVNTxw1u0f
LfxnTyjq6rZ54sGtCqSr/I3o2Je/C1QTmf9PMeVVHwDZP8mpDOxzUUmcKG2mB+kQ
dALj+DkgQ8YN5fNn8oP3batQudUZkN/hs8ZDFjEQwTS+b1zxw80XUs7HjLOfxF38
Snkbx9EFLoGZaqvuQjwuM0rsQDDDnlfwl6FtvjPRRK0GuI1A3F2+8w4bTxV+Q23J
ASYwIFZTB/v2ZRJRSZgrLtk8HDz145jn4APqwyh/mC+jTJkfCptQlAc/6eC0g9K7
6w5U2DovPAQKdbztPKq3xK40jfGBAtttUCTAUnndUb6GJfs3B/5BIdDoBYMYVRHh
OkQXExl8OvjyVlyjqAReH+aTrPKpDD/Qa9KfDg/X18rIY4FzJXMdKZ3AhsNHaqdW
MtgQJ+YmXfjkhwE9ybmMb4sh61A27coc8uiS8642yWuO/G/oCWv+6xEDatSwkWh7
WmMO554zcDA2EqDyKbnyVjgB25tFqoYgoCcTvAV7B1bwtmnGJsxFMYgp8MB/EP6k
/GBSdelPJ7rnldgRVS/7mxCuc0RUBgS3DZery5NYbMkPYT6YK7Chnw5LliWJBMFH
gyIyOZli5lrlXQ3HXFrqt4dn6D0zyqJFfle9zh+QfZchg+ZD9c0+vt+rGLXJ/cc2
P8a07/g7jDIihi33KWGwsd9V3bk2uvIplAc321zyBCGiZpyTpaeQc4GuVNeKKlsR
2/WMwQIj/vST5JE+1FDLirTxC8EpaEyg5S9ZoueC7c5otEwJHDjoE/b/jFVFHCnn
FY4ubJNVJ1tzbaAEU0hyZXfUQHBNFQEIEWvO5Rdqx1OR65Vz3bbfSqBsCEW9mDs3
0eCfozSqNBGVG+45dDnI/9wSIe1JYFPTKP21JN3J9+V2X1aHTtYLZDDnEBa7qKMv
Irrpv71r2a+rVywRSEH9UieUGQs2cQ1qdoGpJnOG/nZ0yfG3SEn1XJ2XZmEQbhI1
xZzobdivfWvSUAE7eLMO4Tau6cDZKvnh1QXq1FisHihclPLvzpp6peFqsZAfi9il
lKgKlsq/f+x3F0MJZ6/lZnLuF7FF+L2HMxrfNzPud+Ie2fiBE2gODAOoMQI9OXDu
mFG0F5Ipi1NWYcYf9SZM5YfOkYHn58mKLI1qac06xho03LR5p/hwwCM3PiXbywhO
1a1TehvSICfOOrx3+TdYdnd1cOrMm79zvFU3C0m2xJxqiUeBfzYC/2lRBRBBm8ID
Gx1nbK9FVTDtUMQecTYw/QS6oJRzYWImV6AjzOnwhU1hS6P8AhKGwN6aMkO8+Hpy
mfK4apBIBfW7ghtyC+g1g7T4nkpoLiQaxyZSu4yrzPrXw3UcNuoNlnZOHn4bfFft
raiiDcLjvhFMgTlAOF7QMo1IvtEdjJ3kVHw9MrFLba3Cuv19fByV065dEIB8cU3a
dOmmVodtQfo8oaZ6ySqz2iTjhIGoOhvDXHrVF5ZHq3sDPIrdY4WX9WExQbZ92yrm
K3VDZPTXJ2SqWqRsjTFN2KBoYsr4PE0PTouBj3dboBqP60AAG41iQ9Xisct/fFOz
B5p9vbd0ncxIy1UhgcwaZFLZGwL926lps1NL4X3Bik/suYMaDd1+8VmE8Vf5g78Y
SWuPsb07pjDXik/IG1fvD7iJOo2/H65aGVTmCzoOnPK7NgGbNYm16tsFSgIIehTM
s0a6ggsP45d8dbQfg77Sxez1s+fqBjfsEDXdn8r7OEQ1ntwHlZu8lctL1Eoi+9UR
/dkRhEj5wxpqT7OTXUsGIqUv1Z1251inr+xM/pxwZmLLwjrZj582o0UBQl04lIWd
YSF8N8i9XWvb7OfOwsxXdUL4COTPKO8appgvR0aCPX7S7QK8E/JhTjC5Qsyj3O3o
qHA3m6SYwXzYKyzFDQuN7vUtSohnt6gWDNq4KieaPz/D+Kd49fmo67FArlsY41v2
qQbDKEt5nzTCKLObhDlblAHM385WXyHxfsWC2Lzcoxp+8bwgUZZVkidzd7L3AWyy
ZTqDNhWv0o5o/9zuugeMn/W7YfRtrglPNeTSJvilCnFC/wpIg1v0KrrSkZp1Y/i2
+OWJn+K327JnwZQosdOwJyijTmSayABDzmpPdzM2RH7wrnguVcCGGcRKce08CCUx
1i9Ai/rEQBOy7zOxC5qQrS/fszZ3z2xJ5zgvEBb6+m/JCVYmTrkypuAOPyhhpNlk
azbAlvFXvwF/Kgj8w3EIZ6SqQPvPE0lh/hZTYWWTIMfrelL8l0lF1SVM5A+MwTv6
+w/7ySEnR1hWnIs91RluFgDz4J52GRiErdlI/ApvQ0EpbKu5ZBwDbRcJHXoovKn4
Erj+fha+XlujG4icAMmWOpFNV655BSYEYuH/V3KBoV8RC8kt3rOj5f30zKhSTuWb
WlPZR20H56wn42CMiKp6rOduTcAt9pQyvz5GGwNm+BQdXfew6J4CUH5HvzFpHwnx
j4kO8sjx8lEWNENuk7SBdgqHz4ER/MnPpgbMM8DFYD8KF8XVvxeOvqp12M/XCOMh
VTyN+BZK7xlyHERLDFlLsnEC4xbz/EvB4gWdoCh+6vkG8iV5hP4o650qPq7uy/Hk
6y4kYOQjn/ibHa0Ec86xu7DNEAe0A/Q2wy73EyfO0GNaOlDy+UcUE+Sj+PaqTzVH
Z1aJWhP9Znjret5qGyFJDhlT1DS6rNsxC4S6cuZdgWgY7elHVT9npQ70nWI0hX9c
r2GLq70fd2ERR3An8C1KD6ou/lZvYjxLZWirWdLBJNqLQJ5N8IuwK8qL8tvfRsav
d7vjMLi+mhuBd28LPpGegw+DPbFhtl0TwjaNRpYyfbilAHjZw1jiIRB+9of/NRJS
C/mR4mg+BmweFeq0YCOK2omuw9zLQVME/zNbkkjJ6bBSWxBfLs+2alBMJ/jwwUHO
SYVzQFnlnpOIMyUec6ZcxEtzsaeRXQWWHWYXgzy5Cgmi9leo5Dac/lDw7332FbST
e/yQj8FRkLNosH9Sk7aiMhBUMtk+7I2LjjZ1NaKz4OqUn6ZT4w85U9XqAplqOimm
jVkUXbxXu4ZORMlxJqUxcSNzq/1t1xXiOFsmlvd8kQbisXYJYGO6m2eElGZC4Hq8
Kbm6FyKZUdiJ7Qosd/fXzuiQndTPFr3Gi2Yu/BdGKsoaGHjpqUIXf1QRz4r2Uh66
kbIM8mZevv+UCaC59blC85eZwM/Ynz0nfZHmcSvwc8OH0ubs9LWya7o73qjvgYcc
SFBbNsNOCc+YlAi0KwLpakOPmYeWehq5Z37zvNhhvhNEwpIO2oteb7dCovJSKOrd
VerdHiNH6ycEwjfaAo9/pyDb9X0sST2IhErA9g+80IFjEEWJtG4/f1oD7/KczYvH
VnV2hdeJLlzLUnBrk4cVssxSn4QZz34SuLg4wJOhz3jidPoJD+LBY4LfJ6moPeHv
eHPOkMRzmBD54cLvohIr8EraSZUYb2pfvN6jfxaHT5UF6IT3Ub2Von8TBTdun6m9
u34ZmvENsmpPghNa5uwGtLdOwIkVT9dhWK/Pm5N+DA3pY833q9icl9lT2iZoxJQE
5aDAvECJRhR3G8OGJn2PYBIsOBtkJYdROv5CCGiU0BItAiciiU8n/ffWioVaLJcd
k99z7u0bP4gbMB3t2AWZxNydFuFIUoDMpDK5KL/pJnUv51Ism+6eNzmlVhXAc+jz
/6uq0V+uc8XaqGzaak79c2INq4nBJmwChO/oKMv2VwwjywpE3GyJop/BtW1XJ65b
16uACWWEbGfneR+gitfUDkWHJaw0X5eRPClMEaEcUl3shsxorqIgoOZixjObgnUy
q03G74H/ZkHMN8BYFQTIUlWc+wQOmZx+JYGbx0ypHaBybjmbjTB737NM8hqdYIF3
Dcu81an+vfGVKK+xx8J3QSoWyYr0tVA5pRLuVGiXGp+YX5C7b9dxPKjwz5p3HmeG
fidcaVdiPKME4V95I3PdBqlSsv6MJYlNaUyz6yR2IZfEyp0lHxnLWo4j7POuMXBg
indnCIEXYedX1mrdvlrg5VNS4Cek2DWN6SH2RChgWEE7uBSTzeLBMQ/ccjRcHx2x
ZHH0AQ+V+s0p3CdlKEzUHqy+ju+m7Xu4HXxQ/4yM2e5epuL2Yz6UufcJGKI5qyCM
sAuTehOrJYuSenKbOCD8QJoeChWnrNL8V2x7W6bnG+VdrC5/AqAuHI1sIfK5b2CC
xHzBktpRCz+sZBI8mcIihYlXGOt5DR1aY6vMcISvCQB1gpS5Hb9DKMnW599iAZUR
IVY2/GAJUUx/IY4OAADTlzDEUsQLLlMxKUYWYFQGIcMkvtBeBZ0AlXJ1OfXJa9gC
oyTRBf0gE74/w2RLAqxvYwmMuCzAMbC3Hnr7msDs2KhqaQFKHu6csXMBSlkewN9H
oKFYQWZvNQhfG0cIdNBbSbQAwCReGPML7qpqx2ZdxkZXggAA8Pu/vchv3uw3ufgo
gSH47jdklBU6yOx7k7mLJPdjj3leh3nYct2IQ5FR5OdHzxlhw8Qskm2d0dk6iaoL
EPZSObLG7nx01ve/ROKVo/xrFSc24eXJOEGOHU63lHzXFt9phEHv4ENstbmUPQI/
zT5WToVDe8NoudKNk6jCBAe8OQuq7hEUlFskkQ7aq5ZVlgPyHbP+FMGaCW9MWaWU
UtcXSA8Wz43W7+ZKus7UDc0wwE1zQ3muHZ92s43ytXRGnN5/cVS9DN5cIbInqwsb
Iueg7itr7va9mtZh/r4jot0LAjDPaZJkKp2L36dlFu+NiThCMPQV387usyukQn1h
guPBYFlG4Q9mSBVLCJn423+y3deprawCp1ns0+M7JCRkZdiwegoa52LadLF336in
vszmY3PBiwOGiLIV72+I5Id/TAGwnxFkDoIsBHLRiaIulRknoxrY4Yk/hGteY5D3
CcxGUFBPXGn3NmeuEcH0h3q1GvMGcZnUsua+q3Y5RVwcXlyaGH0f80tp75eR/okE
8FS2jdE6MWvPcby9SvdgtFeQN9Os1vn+GrOSWqS7pH0h3SpRPoxfh221IbWCTBjY
xVp1Y/u8nKrNICvL7A4FpbAxm6AqIgtDXnfI24551caQcM9idPJoD8DmvgSmNLjC
WG4wsCGetzhbRJJBFqq0F6yAdu1iTKKGd0a9tQHRmAMSlN8tKztxSO2ic4yQv5yg
tC2kz/BqHlTO08c13ScJjSZD3JH9p1VWONPvVEk9Ub9BTk0N7TRSyfIZ643CQNAe
DXZYLlEeUPf3sbUd8EnYnOQQMnmJxSl1Kh62QEX8wGA0g7Aq+7KqojnvI1+O51a9
H/hnbQueuq/ynB2A9OqtNuA7+9K/r27xEH1WLKCgfymAf7rS422MrQsXckJsM54b
C9mL7iAT4aHuZN7cZI7zBokrjxcUVqMcqhrquBJIZFpDTC548Rd9p/wcrrRIDha0
xUpCDUIQ6dzsVsYumkqslbSfQVg/onFOG+98skXD8mFKchCbcjKDKz6l8B+EN3ie
BTc7efLJwDIWKb5VChCZ3I1wwgLD6igbikGt2ev7yRmwKw0vOUQose+YVxeNegru
nRWbj6cl4Id1hE9ozXBYWb/S5AdAi3+G6umA883JOXP8H03JqJCa4MWoFc7GWN17
p7YoWZiqNIMZijH5rRoWf+/ZpeUUeYXbICigqQbkuxH27tzpzibjWA3N+0lzP74N
v6/k4IFGerR8MbMxzfQzboAzTCaC4Nz39AmPE6IjwWmZV0MtpeTuAdhlfeNixQxE
L5YUyMEyV7qguT104os+MF3z+ySvILarNyjECNjOOwQ+3rPh/JeCg+v2WiwHBnm0
bP2mB3O9DYDsSTcSnN5b59fi3TI2/tWMoIPpwF9H45ZnYuaP/VqMmFtidHoedkNG
R32TFJzYzOZCyFVMeNPzL/7/aowjskN+EC4xofc0cHgJCP8+inxokm/l58wvzEJq
yVxXzq1QkL1aInQ+SLF4TGbkB5EaU+apRvKbVH9RxCi6WzRWVzpnKOH9sGh4mHtS
MsljPeHO9Z0Zt0i5zZL10D45I3s+WncY1Yqm3U/SJpyGKHRK+ccTXIpKtOh228nK
SZX9Uj8vEhEVKUxHNaXG800WMo9ZnkpPXJUCRKh0BIdXL+r+RmN4B3J7w5tpGdoJ
yeSlMhS00Cpkwcolcky6cM12dXnlVCwLwH90MEot6D2BwweENrU6hxoRdcsa5gBL
4LjFl+9FbFsjr+JP1E4Er2a6rxiaQbZQCdSFLv4M+V9oe50wOUsTpTJZcBd3YT99
rK9OWc9v67Moac7RARpKXBuB0OSf4NWQ8uzFBYfX/v4UcugVeCRLJ94NVn1QxgjG
0H14+5WqM3aHdHnZKhzyA/EM5u5lvm9FoUBeSxHKwLpONd06Mt0d6Lb7qwzzm1d+
WeBCEWakYvUUMeVKOBDhervxtgpH+idOnA7tDdRyhVuLsW65pViOmyE2utzdOq+x
fnTYF8V0/Lkz78epOovPkRPBXO+ByAkKoQscRHNmK/jlWa363MEZNyq6OJ8+5vZ9
RafQ1LUomc2URdZnz0RcDTgCvQjJrbI42kp5UoYJv7EEIsmflsNd+rG5cK09FsZF
JZXz0tVceURxIGa81XB5qyol8Qbe52RL7LK6jWOymEeIO/S/yHQAb4fETAq0Jd9u
NTYyN5iRzrZP8+bRNc9fBS1oJNVP84N1DCKnA7ThQ51YFtg7DsL/YAXUxiq9gBGN
x/Kel00TQxnYXwJ5oxmTC/Ka7qQQzqdt5P3hcBi2q/hGlJJsCOce/7Sp4IY30tBX
6KtPBFufbYZFkNazNfc1OFXaKcyAcUN14DE8NZDnrsCawMKQSI9/UIjpJs2rOCQ9
kMkswtB3Mscqp9eRqbWYayQkLLA86q2d+WLjzEbD3SR1yLBHLu2gHy5DXyCyCIl5
FtKSI6f9vJRCdIn3I5KRaVGNWKiC2u+LPdfEkoYNXYuCKJ1HTiqdeM3g6B6FvWPd
kBTb9Alk+evd6NBvhfNjldNI3MdOhoO03CqqMXUrCB1d9Jlc/zv3WNiA0AFkaOOP
N7aDSU7eB7rHeigSKqgXt8poWuS2D5sbnDmM6GW7ooHcljymQMOwiZ9lm68ebr9M
EVUjCp/8LZeBDAn+pncVHKx2v3LqJk6RqE4X/YnCrYxoyd0MeC/8ppM8Upn2lj3i
ucRrqQO6MsVdWsInhHMMqSH/lNWg43HQR718h+9elwzf5yd92P30mk0ZYvgZ7u+7
mLK0sGzOzf0UycEDIAU3k7t6LnkD3itK0b3bIx6Wp95eJvAt+XKW6uUww9qy2GgV
bOwsuaLUI9TXnR0p86va/fIBw7RcNhRkG8tMklATCgSj7rWDgLHYX1o6qMzIXqrW
Odqun4WqoUIVonZptzJ2TCxNSwpmjDYxm6C9aHY/px4+nr4E1UgFtMvfa4v8Oav3
6KYY0FX6Wvfizp6ofxR/MGe33PKM6X9+++GN72CfiWR2/fn9v0qqZ6GqGPLtssK7
bHze+fc3svZEmiBWfRmMOiRXM115Lsw82jtMhvaE7QWHvWw0gLHKvI88WTy+nFfP
B+r9AnCJjsjzq6flxc31m7Aq3GMuUlFuLHbfvOuhd5eqMcPDLflP2XSVIY2+Js37
DWszSqdXyYDRMyo023Pky1te29JvrVPRyrrphgcojS0wfqcBZZ1KD9nO9TuQYxIU
3XsYnTlvRV0w53w5HayuLrnDhTpfH0ls4Brbm6133PAqMiIzq/3eJ/kOMLOnLL1i
0VbKnbosv5bc5hf9uK31cdzQh4aVZbqXYRNcNJr0/pp3DKT/MFI7q+WuUL2GIhRQ
u/gCcf5x3d08ok0P3MgXbMbYQEMLZX1DgomsQcLFZKzN+bfeCao89aB6gohmGR7d
q+rQSWDYbvMUWZSrXLWElkyzcJq5kEUJyz8U8xoWtLAm9LEGrMg3xNTf9vg8xIOm
KjjJ/l20IPRC4DUAQLEQhhZjsGfMVzTsRSI0Nr4lkZVLNfMbT9YRSL6vrk2G3k8g
bX5PyLxYkEycOS5dH1+yz5XH+oleEVC/YgvMKoHrC1RVIk3pKhVSst9mSZH2FOkW
dhxfNTFLLf4QFT75vxT2OE4SVaxwEL/iIGEaLQr31N0ZHnsKD09kS2+0pt36ZF6N
n+d0gqtxuNTmzDCLGynoOadFen+kWGsRxWy/HzqYkpmoPvSdULVSkIDkrHBGFuWH
vU+d1/ah/bi/RuE+WM/xz8RlGx0M+N4+QFMZsI4F+9HwhW3WCAq4BL54oL9lf7Yr
ha8jSvF8QtuwIT/BWfE8Vg+oOsdAtbvpBQti7JVDxs0duC97J8YI5wWOJvxv9TeY
oiPy842Dxh1GACoj9o6smDjpPwm+ufDtZ63pbOwgdC8QQLOY+x90Er6iqUiZmYSm
DZZonW322wL879OWSeIU6ORBBOR1fVAFno65srV1EWCFkTKV83YgKzpkHRyanSBp
NJ6lhBTjfcYI1anb93MAGMn1ZEC2ewznCU2538ZTtNqzp9DosOxEw8cZYPeU6IWv
s73ws7F0vGG1r3jRlEboxKflMQPwgyEyWpPFbRJfgt4zOXrORmy4GmM6Kbunq1GG
kgdZTPLUjb60JNDVVYMgfP1voEQgToQqtH3LqhPMHq3+4MMTIV8aKNFT6clr8k1T
rUaspL3roS3MycibEQT85hlUCbfotb4RtpARi0bevWbv3le3hO6cOZOamVic/z6u
yRDYXlQ5eJW620OTcYnFrwLl+Q9fMHs0lTucDAsArqAD7N/Ll12IEBNNVTen20sM
pLg4XQcFKWNfeFvp8u5Ds6XqqxvBY4VvKnWt/Q3nM8zHF8f9cSnlDdFtwUBpVhnf
wvzWGJEfiktaln99DZ/aWGj3VoKOvCa065Vigpi4Bxpx3YcErBru4Ld66axujh46
BrS+JR8/ELOdZlsSdnlm8scEeGuu73j/faWDfucpyJsVz5sfGeMT2zUwx8GJVzqh
3HCRgMBcPyBuJloPhGF8vS8HcJDNseE3o/RGoTP9b1FiL9SU9ax4RWttqOoFCxZF
xsi7/NJMxnBVoWdMS8vRJH0CUEGaWjkYdLkXqMJ5CMz+Gd6djntwUSyVL0JimTSW
6pZVlmEpvPR7erKA8npPkRo977DdzXFpITTVinY5I76+TOE3gp6ajTrReBl+c/S2
uv02733qYJZ2GinoPADnK0BpX2nId4/UfiMuAbJ0Rk6gXC3hIBCFZ75fmz33ss+j
jqF0relrrSSlvBmyyyZudBhe2Lp3YXZIy4vkGOgOIgcOhsrZPbSVSBTJXUgh2yRr
qRNVrET3poSqahM6h3m8/oICb+koRYOZhYmp4YemRonN0J7KlFCR9a4UqiixxVRW
WLlQAHXunnAUET3geg85fWHX8bYAC/DZEbdzy7CXFqoK2ICfnLgJ9aUJEOww8QuE
5q2W9qTfnpPLVK8bmMYD7vFy/n8A8dZGbkPqu4fYAWb3DYzEt+ygjV2ZSVO+rQNj
Evs5eAMB2VuYwykecjS2sMhDtz5f4WWTTlDsXQbaQ6lXFwhhD1Flx2UQrpQaZ5uL
eAGUPaVjyeqSu/pa+xOpEf+cYflmaUUtaAtZkSdyGDFQZJXvkPHAyc1F96h2faRU
z36i8TRESGj0GBbWyumLi9QGLWK6eeb0Vdaw5ndbanKlHdJ4YA8z5f7GNI7tTtVb
BOBnBIustL6RKBhsjCdPWKlcJzQooC3D6nP8m5xyDfKlPTDuMk+Vo4KKN/adCYGG
+ilLSqZX1jP3/G6gIxP3KsihpmSfrhdZDgF8fTDfE3G7m57k7KIdpX0cxdcAbYZo
jMk5zF6FspsFI8RFJPzyn26dIvB09D0ZPUPxoT4XRqr+j9kjh7GWtBdg7iy47EV+
k8FVZrq5meif8q8xd4E2gv9uHj5mXTqMCz3tiZD9nDnKSeeUtFGqchUFIGI9Rs0S
rUOkF2PWJMflGM9sUKLXpD0nfJZiDx4yXQNlk9VQsvIf0ZMdnOC2YTb+ap42gOyx
i1LLsZFikWl1i7puXqZGLmt2w0AsfIdOCT0iIJJYIOMEi73J8jAN4cmR7GkD7KNv
SDhs1HSCOGwTdHV2RWFKgTrk8pwhz9/CWCH+jwKsrfiICqvMYbUfghowHdxqLRqd
i+qIqR5bCez6lgXmuNssC4bV30V3rT6ZeRs90EuLwZQJVnJDIRnNYoS8DNeSGr/g
SyRFICYQflI6KiKZjs75R22nOPw/993bZM3mmBBN+y4QWJaZTrA5Xgt0mPYP/Y3f
Z6aA2hwDMMRS/55PJQ0rboTZ/yw5tWaoVen2M6mdjBsdknWnAgHokRA8cJZx42HW
seDMKik3kCpw5SScdZCFZMFaBhoHIDjv9Fwdp5vz9bNGXBIRJGB4ZJpJuSLuLUwC
wg8eELtVrbPeEk0O+AWmrxIvtX6G+BcwRmOvtFxnwwMZbGUKzGLKdrO5JfOkg5KG
97JV2SM88hmtZr3O6ch7fPerma/70/tD6RV4gMMaC9QzCA68AyYh+Q+dfaanwhYb
QqQFK8leg1e+aiFvl9ARn0Y7/Bp3fUJlt5iYe1JaVjKJRco44Thwj4HmDKTIb2Wy
CFw/1XUsadeK24vLSgqrAdh62f77q6AGSuM1PA3rcNRz1gFNgLJ3nrm80RZr91vP
JQ8FyJgMcu9CuuKr5zGloFoOsVCRk1HPOJTOryQLJEwFyVB1Lgp0GmVKf4DL1qC6
kVg2sCf1jV8VcutcNfu+y9mikKcWReuSwVYGTEX7YvFWu/XBfO7B3ZixTK7SyFZn
RCXBY0+b3d8byMUimCFjcRRzhK4SCahCVMsf2f0K6e5abrFfdZt767v9kVfLDQYb
DjJa3/P0+ubkgZd+I1F3RGwHJHrQ/98+PIT2Jsc2o9DgvpZznnojCyaM2CWKJb3v
dWAeaQryQlSAYQHX4A10aAlBcxByf9rstxHouUmT0YaMgCklTnKeY1d8YPkQg9va
Tco6+FDG0EC9oImPPJVNXa/qW4M2GkAV1VanISzMGgya+yIzQfAOuoYYqYXzqntI
/lWQWTKzn6bR/GY3gOF7+1jAu/Xuw6Nh48hkITpfVMhzdnpS/QtzVJpDowxwVrJH
048uB9yu6hQoCdtkrKTbqcHfJirUF++LIJjBc2LuFF6COxsimTyxDF3GKf6tKD1o
vMaF2Y2syeQ6P7qtoy0V3xhgnGnEl6rXkyhiK+jd7K8dKZuNmCntrTNw4W4TjZcl
BUCQ3u2XWaITVd4oS5/rsa6Ec3rqroF9Hi/qH22PUKsQOTVy9cRRcclK+PCZvzda
MeAJJHsUx4hV9KVHFIhYHoMYEdL/r7eZ89uQ2DVEwWGrzGaydgN6rNhlz745htP+
wCbV3/eaDj+8TQSLgl4zv4Yx2JQ1G5DxQis//L+nPU6vjWKBRRWReYobBgDdDk50
pXtMfQhYF6QPL8ynK9sYQJFAwtzYd3nkkMbjBnFWQgdrzoXqMJIgxaaou1duYj9f
BwurVG5w+jewEKtZRJCz7/a8hkATznXOFdU1zccANX6SanToQGsAptce3ZGR6mtq
wcsofif5JkoY1aPIEp8DyKUHGOROPrqno+L1r0963U3NC/3W3xJkeGikfdE9fjLk
QVpsIMxjtRUEnYmydJkuu8cwuxO4g09AAQuT6FOeMm2t3TWi6CZ3DZdcQsH2W96o
6Uc6fR7yI8mkwZjJjhErY5OJCnm6G4Km4fuRcpHcrqeb63m8Fqp8LEg1KdkWXHZj
JHJoYpnTqg7Eg+kBk+6k/JYQcJaU7+s60Nl12Z6u61CLW3L1HNl3aALtCjGNIRtH
oxqKPfpOXRbGUzHZyhsX2n0Gh1TYhje1K7TjkpRHUc9y66q+/mYL+k1ZBkhIib3l
4DEcaoyNwgNlmsRK73q+vlHFVjWrB7UOxOPA+Cjx1gL2ShXbsuIE3vNiuFUj/QZG
DmR6t1jdkmARDGroaFfu+R1C9KhDP4ydK0AidnQYuDHnGqcG3pTktqy+aZuSlip1
qe6LqGrFv+P773Nbk7RK7MkgHoHYxXOdeGsHRrmzaHtFmEt4nJSCAkM4+EGLFEMj
Ydp01MYoFVveOzzMzV6voB+NwYj4WKGxSdMbAPcN5FvTBmY8UQ6KZKiUE9zx3hXW
8/j/xbix3kh9Y/Px5dkrgB22jyjlh7ybYTRu4pQDLCmg+Dhm9MwqvhVfnW0k+amI
w2gmwST4ev5EmsuRZkT37WZuCgJZxK6+z1FIkayAiXftJKfxqQUgoLHG9uUGbZZH
oLvZS1xMmjFKt2Ud4NGvXiOt6BIed7BmABBwkXF8xJsqPnPy0yQwAXXHbd4Bl8Ry
3UhfVit/Tahg55Czau9d6lB83bmRuFT2CHcTIf98KXSn1VGDD1nLdV4vbxuGo3MF
XgCwyjBEpzOyFa3go2afQOK9fx60TlgQwed/NmFDWw6fHgtShnPwLoHKhNN8otsq
nJ0y+00wLIYph3NAtswbtXMtsQNVpk2bOKpQ+GPO3x+CdAIh5cyEPbDgGiM5991z
KsA154YA+ImG5IGUtMSh6qfV1DaS9qgrKua6Z7mTtpZBtjydAw+adfnuxyr5OfZM
vVPyqXfXAN4FjtE7PKU2Hbi/rkupJCFl39wEkSRSt9ddFC87ORhwuta4GQAL3/8W
IezJp55EhQ4420O48q5cKltHshidWD7XbwW2VsjO74DHT2AO1fsBqrDLaswvRn3U
OKh74O56pNDXr5X6sQ1n7V+HkTdElFEFTSmjP7wvDbYGWltOrBjANbyqJDSGYWYJ
hah4lbd0LmbLmNSOwAN8LU/ZfFkkWD1u1papH+HwwpEENfdwAhSkHNEFQ3pVcJom
p6/NqCiYhRXqR935QJLHxjUGrNCzZC+HPpSM2WCeoUJo574IKkLOcnqV1KlyQLzI
xZA/67ASUFu+DiLzL6K4LjSE1kKkHWgbPYHaDfBGH1XI00CuJI2ISv1Wo2MlBI/7
j6UA84EQ44Mvf7NjUmzQRmWWIGVSY+ng5K0R3ib3QhSHmSjkNZxT0ddNgfiKmLJv
8pjnAfcV+20f5YJ1BCfDc/coCbJnOhUIvWGgVebnGhWisaES42KCjCHMAf9SDYXK
xdifmMSRxwl6Nxfu4pu3bUhSb/yUwjr+8Jy9v9YRhyhaB1ewJHyuwurlE7Sq6iS1
Y/sLMrjfMyahLd9CiXhOgLpdknEP6r7q9JjGAgPjPoNMbEccjavT3Nd+k+6G9dBG
Vmy8pJ7kIULqFk8YW6nwj+WCiSTI45z/Gicg+mTUtEEqEplQvwmrbk9MZARC6/gz
CoDggw93sibAG2vup+O/zSGtTQASbo6T6qMdDVUZr+VuhyeDUxIWFP7w/KcmDVzN
9mYr0P0gzOmoIrvCchVB2ySlipx9b9VR5sdODqzd/NOJBWXCzGD8PUbeCK+oOMHK
10OzEejMJsuKfg51X1NZhMkAqgT35Vo7khJEjKSeZvuQ2KvNaJ8MyglM6LqOCkAq
3EueBV+FTC71sfbvEevzlYV33Fk0s2jQ3E69YoZOHXHJgXrrpOqA3f8frMpLE+xc
u/OUfCPaFr4b5bJGRQ1hKF0cnyG5ktquyf+nrbOYfL3LIWUNpEPcF4VvLfASrPcK
JYGkFcMCN532mGZiWKeRarhSAxfV6+rQxikP4slJI2ppoNmOEI+FfiKByi7eTK50
0Fdq6Ncod7v9xdGLRx9JsjT6kbs7UjeHaJQ9eRVnno5oWBIqHf46uJ0NsqceAnv1
xxXq/cfx4V3o7jM5ZID7svkvDOH02uO4TBAUiE0Ky09AILVmzAXdVwCaSLuGtkcT
LeeiTNPu4I0vqnf1gvLcf1FDLE1z4rvVtjXWuRR/BDbl4Hwqurt79LagwjftatIO
A1J2PFSQv4Xf6c6niTfv0LZLD+ZXBUed8dXP5Zciw0jdrM/ZjwB0+3vDEo5G/+qy
I3R/VWekg2CwfuEvva2RcHhHDD3q7YWi40W9DVuY5rXA1J/7uiVeQ0kNm+zbT33U
sFPoVM8re8XP4pJiv0YMh4zyqDjJ2xLCG0Z3+t7segLmQWA17eylWAlpEwVrcKsD
3rkT7dv9DkImkR89uVlx3XOhu1OEeI+mAXMLnRtpMFbDarJNRad3OwQ5XSl13SsX
J3ddcdqdvzO0mXEEmRv9OLMqfO7FYUuHJHtt34OSwXKWMspAc11UE/XjMNUe6MkA
T7q4o7m3VdC/QvbbuF5XhvFCyh1qpSwD5RMSXekHkIZyqk2c1591fDCT9gjKnEfw
jtqD8VRMxMjeJX4JM6fO4xqusrBIxaG/ooXyTCSL5zDSEgesTQZ2sg4EWqvFGc9+
ceGKas1aeJ5u83nCN8JtVkjA+9oqutDNDTIX3hh4QtrbnmY7d+XHylyhtA4VufyB
2SDKK6/zD0OeJNps30FYpmlyDKG4OmuJPZvvA+Nl5ytPTmpNo0KELOSuzqOMReWm
6uBqxVhI1NkzLcy/qSK64sZaqlIYr5PA+I1UVLvroB2ycJbH0mpFNBTHlr7Z9dol
iVf+Hz4HUvOSMSlhXVdki487lV6/JEOluflBuUVK/eOKNrXVeqYpf9RhTZWZqmZG
MSe5L21/wpAy+00DmYM5SE1/nxG/eHiuwUz71065vLWUZTYtVYhaIk4ScbfHgsEw
kaBhxRDVTzYOoNYrmVtACBkyYVRTJ8Tl51zY3k+91IrutHa/aaNHaxuBY3Vmd61E
Pd1euXyex79vY25xZqF6tOmknB/EJ8htwtfyZA2g7gZC/kgWr7LzyuC7INo6KlJ3
q3IZlvcaWhfRebDPMnn3jRMXtzAHMLn82Yk18I0OiFyqg0rgZbt4WxToEXNPDRw6
a/JBfbm5pCEX4oy1uVOjIhEtAdYQg6OuOLY1bS8VrbZZp5BpCgzh8Bn8bj0RkPZ2
yaoGZu0rUvDURfgCxNLpX6PsbeyEd/UfHPfFkp5PWVoyVN2N4L0OD1bYLVdK91Sv
3uC6oyPb0mmUZA2Tw91FmqF5CCwAkV3WlSnAZvZlbXw6tsdzUwIvGf1r4LCoPAWD
PM3DKO3OT++1aAnF2Mj6J4vaNU99Zrol3w5zNzdlCUqAfJpZTib2o9fTf5/eHyjm
UUIAfgzOIX37xoCb4jCbl39Q6/HJKv7O4o/a1s8OXREPzLdPJOH/pcCzh1nQesZL
ZBMAuL+MBbeT9cmLxAHpvmBxLs33Nbon3tvh+VkNhMwE4sb7VMSAnyGgSnRejuh7
6OMpwBPpRuR0hajpAPPAKY8xrSfSfw49t4zQ+uzpWaDMpNsCp+wGcKIE7Z5MDItv
hBWTDjLW8mT2nps3YP2LhQ9WCquKJH4JqMkFmS/IrCPfnDFW4xx3lME6sJVxHRdu
lJPQN2mlN0uFSLxlXbyOjT/DyclpEO1yFx4bmmHSTJJVxxsfSEolnWBonX4ptvoG
M8ELud0d+peDv6BRuYpGJH28qSU2chRLaauo1JhfFtAT2wcaz5AZqB8rs4fqHT00
xYXW3nd1XpyJjwZG7F49ZpH/eaDTbXSDyaMn2UNFEyvguQlexLDnySVo/uIWw/XK
2IZLl9TO1FVMAa9NVAr4CGH1B8wPHz1jTeMiUpYTAqa7jEzqpRDEMzLABCAM+hLb
McXqdZ4+ZXzMiw2cWaPRcpCD2dUX9hCH7+EBnvMq9p4KrVTIZQHA6rfblcv5wJ8I
Gru38ZgvOT11Fhdxfwc/7xuI3i5+JGbdsNvV7/c68OcY2nXsCCS/2dnOUhqxjX03
HA0MEocx0ltmj+0F6aYfQtgAGOHCAEon89vAHGxPSMPPyKIvt/OyC0dqGWZT/rGn
yyS41z7GRpKDfCeU4Ddy7JQWHb55KuZEWbRoCvefuEQ72sQ1YyzO3OhFO8uXtIQ3
q2GOEJYzqd4mqwk62jdwUDK5+mKnzhJ+v1PWTr8rBmOGm5IroSShKx9pILzMqw/r
aP5qMDtCmzhxqPP7KLwnIWuCyx8PIlZfk9P+CxKNVb2SEiAIJqQ48AQ7xRFIBKlW
msJeF7eM0HGho3NTd/v70HAz9f0VsmF0UykpqkCVfMuTAZ5QQgTc1eSOhBQJP2Nw
KptTHF3pn5IBM8g/d+OFbh/wp91CKMtphTdKGgrCXtROuGmujjXhN4HSr3sPttCV
ZvgdMOCTXQNKRLmu3xPznYEjvJP/8WDWiLSso9jh67XM482r3lJCs3EctpNKtuTE
b64z/NJCm5lInME8LoyUVZnWMDdFuU2tHcoFN0pzxHzJfbg8OGXELpgmPnjgf/mh
qC7fWDFh4FO1J/16+YFuMWfdesr3SLbr+VraE7BlOMfXh21uKDF25cGJDeP3g24l
/haxa1WGtKYYVjGVJBBpQCo9h1q35qiAU3SjMAq2A1scA8SGppwgXMvKGPyJjHbP
5sUeT/Lwy6G6rHiPijLTG/8zRitUdG4MVx/ycnwJClMmFSd+TxL1bUyt+MgFZpfd
FcV/sIf5AeSui5anqw2LFHwavdfjl++/bZRKH4CpMDJOSzPGT9iYqbWtFCEgmPXj
J0xp6R/6rNcYI5zzPeSCU1PlgaCdBS4zNzWm7AkKePB1pxbOA2iXhLzCRTtToH7U
00CxbvnNZQkYr1mbYlZ0nOLgipuqVtsaijJDib2MMDx0iLghShX95DmoVIVacHeQ
YcktJJBQVwaM73DL3c9BFTH9fawk8TUzEMirbR7m/yWn0Jg6rGvQb1vNAbnokS7j
eChfWy6SswOkYFWWGDbi2F69mgMDnq5MSJwck6E2J90d1MwsQb5iTmLBmR1Fl0gq
1eulP0nqqi/E60I+lW3+bjKpRCjF4tZ82G3OcGtOLD/RrXr4FACY4xxwTmtKPMej
QcWJt3T77wbwClhSuAsXU/SC/+Rb8xAIh2eguW7Yn4Lx2vxksMauaUiqACheulTi
srAcGiKAigeKduoRPuel0JiVuhtJXTQu8dBs/7gx+fdlJdu0pC+5BpV3J0tzMuwM
oQ0YpYtwc1OEiyJDOxLUzqsm4CsXKwq8Iu9VccMURW4wvkS9j47e+YhKaM8Bja42
MHfMTh1u52LFUTwRfqWsEtKUC7j4JcZf8s9uOfS1TWy0yUSwTQJliMg9VplCzs7D
5skWyHozFVVmbGA7JbMCXh25ySgZpHqEpxQMkkhkTGlx0HjZatEDdu0VtRZLEBgN
wgENCjS6U70RLe4ZeJHFEwWOOEs5+mmi5qosnNT4hjE2+iy4UGIf24znZBFdV0vw
0f3e6BDkmFBGQtPycXxC79Vs9WD5ju88RhFfHNc56r+RnjgPcazzd9XQrg+If3Oy
iKBzVk4w5SjDkXVVTKgDbAwKN+Qlo7JpR2Rtr34JgPc0cqTAU1mBiI1nsqgKRDzo
4/6nl4nLtwyStUMW0T5Po8X40h+7NZTOmaNsxQqC62Oxa4068qbI0difZPEXzLoh
SqnRbMDy1M5SpNKFR4vcszLwZQ3CfgJ/Awiu49kx06jGqXHn25pG0+ulliGxupf9
E1JvZJWi+jXrRKOAxStuxm6ohpeoNgCEgOiEsktLIHeE8axXLrg7piga7G+QF+B7
owe2pZW/i2tLpQ3CCriDrujr2VNePxVi159HbyEzJyXtUKzdxmPCBuNUeDMBeMH5
JxsvPETFxGSjx01Xjx+hGEK0QMe09Cm6dqkVbAffxgvf3NdMaxVviPH4sNrj3z8M
g5PqWopp6CZlKkBk4oyS7GTg2jScjf6Yog+Ruq4Gx2ovBslc50K2EtzXFivcE5CK
988JYYbqn7TAEXO7s5YIpL3XFOBCjd8iCIijys7fcIFtoLsRYJ5sEWojxq0cpL1R
ou4OcaR6me5uxxh+cLqUOb/q5CXhIElr+RJa1uyy1yw18aZXW5MBeKLB89grWXez
rX8ip9AnuwjX1MumPEMesr/49Uv3hP5pKGZn+DJIhG+3lG3Krlikq1VZw4siG4H4
O/rtysKkzyUrqxoVxIRViLMnuiay9nw7czzwVlyKzwEKcm/mQ8hfEYPzklRdPtVm
squvf7qKFVMLUzydDLB6ZCQ5L1OFe5DJmifN+XAg8s2PrJ0uu0YvEvAoAAqMeV5c
7a/unuKqWK7ZTKt3UstH9e08TA3VppQo2VD/Da7N/itvtwhlq7JeUt1nVg6zhTRN
K7SiL3rIVHGLDM5mRjLZ2GCA6yIhfpT3+X6SXCDcx3IwoVoe3Zxz+Rj3DILkSeiL
myvgtVb0ViGe86BvIbBqODtgPTlyxtN3FWW5jUPBvtprx/2gCvns4Q+u8YqUkC31
PMn4JYkHLoQJdedt2St+E9+zGCH9SYabaIpS2Z8IYj0+yx/Qx7ALG0RTgUATCOIn
M0LGwEXoimsvvF4CzBm5x5uAWUoGpxmtSLV/KYjna2Z/68xk8YZg/fb+JeyAlyj+
4hmEN44aK7IQ8eBhnxvg8EX5fa67RGX+BpBKza7ULV3tVSq1uhX4YFgWK9EWgvKf
LtOumJdt6vTZ+2Rf//xIsBXpO7A5ILR/fSezZTDCymA6JVeyqcTSc637g5EbrL7V
7Ek7ycf+Ai9hBEvqDwa9a2i3rxJ8Wzj4LhzQVNkN9LiNlXYOLUhZIAhfYSIqF5+r
v9GeYFkoagPTYfE/8H5EoH2cHOSf/OHQxLulPSBMc2qtf1l8lLGXaNpiXPuApjaw
aGBiyv1Az1xCZMUsY1hflWNxvkjWAfI4ieBcrepKm3dHZioPpvgg+2NQ90uEFiv3
vtqqXkkbJMnAbjTaOZUjMDSVqDewwjBB+V6j5oTT0Z9FQ3+OmdD2RJnbOUM/SC4s
cc0ZjluvlHVDiJj/WQvGie5aTHIc86ZHOp0fUeWIciTywfKhst+LzMuVpQ3xakQ/
hSVPVcLBYZwMRlB2pkxAz/2zy10SfpY+7X9aGbYzx4wGg7rJC7xQGQKMu7FKGTu6
xGZP4L15fOT5X9qCWvxFC6DLuqY+r4lNdRvNqHvqODM0CB6m6Ir5Rh7Eaq7c+/Xv
k0bvFxbx0rPecv78u/Up93b9DLO/rTvUIKoBcitTr2AT/ueo762kUuR6yzbsRfnN
ANiBjq7+9xxpmysv5veX9kOdA/b7Y2LWOnKvghy7KObr20+Fk1GuGtXdsds+723C
7jZenSJ3/c78+XF6rEl4diNprgJvtSFlX7xPLA7wnEU3tutKSL9jjH0sCo3NVi1u
EYX271BLHc1ELdyVNeBTYwInsu97gD70Oaw7g3Q7o20Q83bf22SHkiDhJ6Bvqh2G
WwbKpCS/3UBRONMS0mPhhTv89jhnrz+Fbo21sW2/T9UqB7GwKnU7v15ZBfN+sZzm
iWTEO6VTGj1czG4eMm8iVOH3r7o/HsOmg0aHlo+N7shhmcJyRrAb5CxSCBT/1VnW
YLGMFERcfdORmkc0sO8CXdIiyhKNw1kkYtmGmuVko+QEYaejMZB9/ifuyLoOHpK/
7Ow4OmJ9LOmJF3RLqsK2wpQhiQiEDSqrv0O4d6DD0SxpnjseUiV114nO5ZLOEmOx
5DrBlICtpCLXBhqDXbtPAAkEsA7Xjy1hFfIksfFeTmT1DYomj9rGFUR68zaHORU2
Ruj4oVM/Pf6JPQvb4kHtLKNVjVyxH0yx+YAoh2+/DeLN68l7YGxiOuK+J8hCW7+F
ZvbjUuCyrXMss+rlOjysqhdI4P9LAmkd/CLRYRc++exGHYxE1Mw1cAsH3YQ2BM1Q
OMXT/lLLwHzVx/+tXsvYUPDT+xv0DB3yqZKqsZeanaKfOa9St89BBxShfZZZW3H+
WK/eZAw+Xrp08ccei3XcCEfXSWKXMNhgdgshrpPdvod3oCx/l4kx5Vcnd1iH3E+V
LzIi2EIjgYzMvMIBBggnEUOqIeGHXrSWD2dzVDR3GB1z9CE91w5PiL6+2UwyN2/e
7bQo6FA78yc0h40zjvLgSHOoNJmc+T2VFstMcf1osQ/NB9897AdiALHmXFSs29Ga
w4LLJRMoN2nFLKekxQlsH0Ix9ZEky5QO1rT0xFi/wXhRnB+heW22U52bPDXgzv8K
sBxjQJfmrIMnVfw4+WIAhKR681qRQDpEwNQe577ayVAM/IHtGNNRzzprcgwPMjxT
X0tdGS+N2dqgEruc8D9nW+fOmJKObP1hES4/63XCZp60spDJLrtUOyfieLSq/WT3
Qy+9df2Pmsjw7Bfa/AYB/rlCcUcT5Ydh3n7tU2fn9re9hkUm1frlCJdKZYQO/rFQ
Y7NH6tR7Hj42BAjIrCzhZrdxYpDj1w4y2s9mil9ByVbSa6O9LUBl9qQHDtVC5c/e
C4rTCXnwForl3wWFNPz8EPWz00wT8ndawakliMf/xmGtGPPyNMqD6f3V2290F24v
UrUCG/6Fs4ltPUv8ACsI4JoN/2WRgEVjXcchSyEcS11opwM1AiNn34quBSukL95H
0A2lnnbvJQutexC5mOxyALeoU93W/CS0wFmp9sVUelADG6xYDqmtn6eSpv6HuEnD
Cd0zU4DpjmdPfQ1C/HP2d8X2dNTZqDjgxDZymPieLndOzZvaFjd4fTba3CAkhsGg
A+nxtgjTMBQcqhxEHB8t0z9wyBAgmqlvEiAUHtzKQ99exFXVSM2eAenqR9ZGYwGc
eZV61E/c9w6zRCZzPbP226Q3f6hgFYiAcQL7yp3dJfXsh00wtPrtsDVa+XVrDYOC
aR7tOXKBNZOGTMTNsLoviVjYTbsUImm0Ga/a0M7BeHPPoWYBU84AOy1VduVM1dCu
j9O8lKxSx2Cv+WmTylGiOJb2wuXRHLSioU/KXwk7Ibon86BruJkYf/jZuVW8zNyX
ZB2lvnvqDHCKP6Gf1I7iDvELFwY22y3VWsJz30YlkEFeUjuv/n52hhtZLT/O+J1T
fUQUFzzbCs5IHy3sWD6Gg39ZndakiCv89uSi7ZVyfzSjUcD1kwHw1KYNVY9WFpSo
8SivH47kNWCfYNAme5zAv9kUIQsrwjtZRAuJJ5/eW1cB6XYjptVaT0UGSFqjbuKu
vh17zGX6SmYH7PqYHZT8uYQWcdHXrKxCkHk8ZLPgjtKswlOezrvGrqgLrxW0UcLX
RwDspsH0S/RNEttFrPOOHErM8LV0y24oPgUORBKb+pFC+lL9GHQ0er9iia4rvMrP
vGPMLhXf8R611tOwJBlE3/eyU0sO7xek9SPQHHwU7kdVC0KjK+eKkuWqiup1R5Ny
rwj2FU2l5JDgHzt7TiPtx+qKMJEhorTZMV7fKrQ1m8XCnSgXaAy2J5VYi1Mo761L
h5OHqg8o8smG6yjlxBz+iTI6yAYusy1tK8/EPjZ0CDFfE3j5YzpX355OHetSAcNa
rG18rPSiFeAFNZ69uIRnSfVj8Oa0J2K9Iq3nNvMcFKqdFLrdh+SY74J039Ox6WoW
oDt3MyBJaRIRRJrdokXuJwaUXwAH0rfOmNN0xv8+Tj1Eytq3+/2lbPI+vkuq4evN
sohUUSpNSRSfTEBVGfWZrjPrKSF20ZMns98D/HajV87K+z/dXWqyqK2ytvJsPe5+
QVnpt0iqk7fOQ9mny1hNwMjXvZ9nKli6qeuO8VdPgtwqM9P6vTPxq5E/qqptvETc
NHUpO9ku1JifmqIL0Kl5hm64tlR3t6J7MTrc9lOAC9FWo0RITnk8b7x6WL2RlJfV
JlIuSXLUQ35Of1O/JUneztbcp0mUqJpDqJtLBFs/k4T07O4pSfUo/M20laIr6P5q
Yh2/lO96NH2t55cgBXKd0eupkKG3hkJWMFEhoVQpUWJ/ExVF2+uNSeo3oGDr/gC4
S1PFTWSQ/71en8LYhnAsRUft6il9acDer1nQT7Hoa40fCjyv1JwDbHJFjmVIff2D
WCFLo9t6T2wVyAZyNBDPd439Ooyr71H6qQ0cYFZe8TaPUkgjX5Y/0f9pyO/neezq
fXOL7yScKJEMsXSd+5MxzhLLoLxEKOMi4TmsV0DvkeNPOvjrlCMtzCHo3c9VoNFM
fvzL5cWEzX1plfIH5enxW0Mh4SZi1bfbR62hs7lNVGAsU5QU9ASnbbnrb3UaolNm
Z1gQyKsJV8iA+zggkHFXCWg/OW8fiO3PXCqjN8UIj7TTqhkZJAs2Bj9Tdmk77vUr
fREgSOzSqDSbPH6eFwkpDhdrK1idhwRnH7xBoGoYGzGd0dkY6aYdbUBzdI3blGZi
r6g5r1Lk8AS0COTI3XqCyIpy/pOBhiVt2zauf9hw+1BCXWp4pBscHTnXpRi3dxCz
9Ay5iwGoOFOunvZd5Aaz74qGNXtY98YaaM1VAWyQJ2+oJW4jaj1s0w/lky27G1b7
o+mTA6/BUMWjThYgrGTAp1bWW+Y1DvFmjwds/fjdPpjkP7K1aW4G/QNT502XVeof
+HtjQYkLiiplo2F0YA5Mmc/jaMCZ4Feo/vs+JYpoCgdlHbKLDixPg+LOnsPt4uLs
PUCfZlfM9pts2yUEiJqAVQ8FRwIm3gECjvCRb3HKVyDWDFKbyUzqAd/NihmYuqnM
f9VkMdiXI0Pmsngeyj3WQZ7qvnbD0Fmgyv3NvFLeFsSl4jdRjyW8P7Q0+O3jsVcU
wfOEEo4mhD+gRQLow6ThTJTsWE3RDKsezpH3VrTVDZuaUPJJrMcv2wJSXZ78rGZc
OVhslntYf7lS8Go7ijbjRnMKqq/mHyDORC0ti9SlkfInyGHvRCHCOqP9b0+MU1XG
sn7vYNiH+LfH5M5vnG+esZrEVOfrtCB48msOocItmqXzrx4TuuqcQ5T6pSQ272eS
JgjwDUrMPOzbNYqzBMmxmjoKaFpr+nxXwDRfm8S4Rqwyo++VKZuvMg+QsB2Ote6e
9XQSrbZLU/U08qLwUaNLBoSDaFrZup06dYgKPIp1DBHkR1Vp63zzrg//uxIcLdTh
tkBysw1Tr3zP5Td0uc5OFB412naXhJhlNGDcm6Jp2PxrFSD4cwYbCVPKv0r50Ka0
EJFyqf/HoMyKbNf/NX0QuToebWhlAMGUyXzoK2ajHrKD+nb7IYshpwkM3oxCjyQk
/9bLQoGB1sLfful2ml1fuxk6Ecz/xhNWB6w0HU1w/PCJEizop2DYudZha+yZLydR
SOX+6/Jhwjzt1G5n5T38lTdQDYQGEMRamX1UmEIrdG/T6CeJX6IQvaURGniRzNB3
5G/ylJEQ2A/sNBoN3b/vt+8BDAQoTStNwVKH/Kmn1QIL8Gaw+cQ3wlrsa4FSWRyL
IpzIa90fNDMIqgqpzSHIZp9rQm6TLG0o+o2ksIALwUiuinPk4ysCop0Z4xhGrWHm
MdxWydieumyXOO2VdZqQtdaZsxt44qmV/Ahw06EWF4OzEcGBF0wOaXr9jW47fsQc
rJQgV/g07f52o0+hEecb+lqCME2/rR2PdwXcdM1RS3YJB3nSm7rqt4r+T7gbdrTu
c0Xwx9YrGML0RQlenxjfFFR2h6ouoAIQzCNVK/v7tCcg66aFMHzpyQklIrg0SMP7
c/lZkfobcj0hdI7v3JQgMnopIAZh/v9vuTnzllhAzGCae7kTHDfQFTu5G7WdIErb
TCeHiOZgqm98rq3b35jjIap1XmsOLQfVTyQzVZ6yy59uVn66VdOyGhjqqBfwVfT0
NkLPdRUBfolso8P1wVvDH7ScRl/d06hoDK743Ju5FlVs+/YtpQPPm0Llev2Hbzqj
OspKkIei9J+P2qkYT9lirwsq0zdtkTpLZxROt587m1gaJrf01sr4EgR7ZUoQxfL3
BYO4f2Q7ixYQox+qan4zg0QsMM06h8ULCSM2mdwlgn3XaKgak4DfuFCuq2uTTJtW
rni/veYBy+xLddX+xTT2UwR95k7UeoBJhuZ39enmNepVw2EF8Pwjye87KmgUJblW
YPPGYTq/vNbOk69WS4uMgpGnmh71qcsXqE+Hfi9cFWEC4af7e7JGB3awhbtsamw2
rdho7vNCITK8JbBGRhDVFK7jy8aq+LxQy2scsgxJgcmFxZN3m01ZglFrokXJ74VI
Rhug9QKJzZYPtQzhiTHyPuuMTKNwGXSVEc4rlU3RvXXBKNKo6hvANCpIJmuuNwmo
fghEy6+13xyWlnuK2Xf0O6YCp86MwL+uG2Y3WB46v5r6NsCoFKvB70PFrOr28f7o
1OkxW3Wt229p51pvUpNxQlD6LIiSlDOxg3O8HXdTfSh5okQdJBF3prNJPCyVr/eG
G5guWM1abqbd0hoKVdumMekNIIEv4srMl4A56b/aJklBzLYLO+F0O6nwgi8mFQfw
MIEHZPj4Ke+DmpEZ+eTJMvZrMyRVcghPrAlHdZwDlASVfYCpBOMsmqYMSk3hUgOk
Pz1KTNo/pvg0xniic0GJ4PXnNzSGzdDreATKts+LZOpkY8O2sv+689O2pU0GpHRn
mU9QdtcF2VFmEXXftLtd/ZkvORh5oIfDQ0EHVwfPXtvG3xJcZ+i0mHdYl8jkFmm4
JUWfe74jukHVU6W6ZtACYD3oy8sgFvDQ6fyRUIFiQBJEuUjKJfXVs+KQ/iH4AU2S
T+ispD4KGLFM0zQZzBdjRCX9mM1j0UWGOlJ/0ugH8zSuKFBmQuZK5fe2FUDmbRiV
QHpKt1iAXTcQ/hL53ziR9d6Bqj6gWhG9xxiXxMrYojAd4X+tWN3ZnESEdyuzgS8J
PzozVgCU67XFHY/BufGuzt/S6sEh7kgNcKuzXGg6g0giS2XPHoBD4HnWrh+bk9ya
iLmpeqlLQGml+XZMQ3NBh/+XTBGLeSF3d782Kij0idkcbt8hb9mz6i84HpmO0qeQ
ihcwjbOMAPv1Zbkd7HE5b5zQllCsWTHbAaO6JvhTKGTMqUPwYpvulOG2ZRoF09Q7
AX4ibiLT4HQhep+fIbwDxJl2ij7Fd83F+PFpRqYANDYh0uwE9jghLHgCCn+2szas
/RvQsguRxjgrjUfRExWG2xrUgOtxOCEzYTnOJvanfwn+xvR4/XGyyJTLcxgVer26
vdkDdkLHmrvfPJMX2pxVq2+/H98rSd05FR+qUCuCj8ZiZBktitUr4tyZ4luXF4hH
KaDV1uVY4tHmhF+En6HUM+10brWKcT6jfMcmm/hytLryWUuOgZE8ug9g8ZOKd18N
kZ6AYJe5gg78YhWw0R8ia8U67ENVpFiIJu1C1I+LuPUCNU8+7wG5St4cWFwG2uSw
uPdwlDERO11puBiAo/PEPaC3Cy3Xomu6PNpnUtWXSCiNSfAAV22UXzIMzGb6PFJ2
vIe/l2XnYWVs+yeWq9JcOofHPtMTpKoLZ52lctJfJ8LDG/aGFnWNPHR11RERXG41
ed8IkBt6PYdr6Oudeh87V2PIvGtkOA3Bm8UCH8+otazsTksGAtPILUcTbP5iNl5+
bH+kxbsoyGnlebLlS/m8P43SdPoaRFOTfYLeK5VJfDl0Td1fzJ1Zw4frxpJgtmKa
mB5cwmqSX53sE7mwmwVJ7y3aItVwJaTv2/sBY1+HtHPVbHi+fwTZl9fBd6/DDoJE
g9/hEEKwE1k6wIppLyOzmhV4eExoCkfJ9LTaqxAQtC6RWv1D7UJWBYeUMGwLWCOR
VZu4PkzbB6PTQm4xBdCOCVghA0PTjLMY1kHWDlT78AHPgWU1BmqrlOwjZ4M4ACPZ
nuxZhWPlcpJ3FGlolNQXUNbHyzsoeWv9JSeO8Twue15sLOUnAm2vzAhuFr0eUYFU
JPl2v9xpM+/WVSjAOIRnKn0/7tuQLBEjSw/teoKw8oTdm7maA3ZXqDWkQRHmlRlV
6f1vS7p6T1vu/RJ5OctI/C4u509oLxceKIULS29JbBp19KH/8U9LY0aQQNznctY/
m4zu8QNljfZDkW8CYOrtpMQ7vZKBXOpsW7ZNUC1nnoy3tRyiUhHKMRYQbIPiOLpw
bX2p7kppoqaHjsdBoU0qeJoF38BScAEZh7xsuDfXgjyEFr6u1cItyY4i1q735a8u
31o6hJxE2b6+sdHc9u9Yn22127Ls2VQx6SoOheJGcORFjTGt/iyuDj3389b89xl4
t5/3pvMdhjs04otvNJNYONiUiaQTay3nPR5m+6svEiL0ZImUYsvRais4ryXr9WJm
2FJxnhvAU2ObSrRM2hj45rWxmc9lyvRKAqg7tosKTrDcTf5ZEp5oxlJi9EuqBPOS
esTjWcTl6yt+5ulMh1fxcs9IqeN7i08cjnhPDhwY7SAzZKw3XVcnSVUDuiB0svI8
ORW7ydRxoLdbwlCUhprIa7H5YFPzfxwJvZSoTu69fE3wzaNshpEOJZijiAicHNAx
qHuGVGppPDqxg6BFjEy3aA9qpbsjaH8WvDX3n01ot8Vasf/OhzjO+GaG6JTcn35y
/KEVS3Tuw9yvNJH08yHNeToFaXU4MmbyU+HNcgwap1wz7eKy33UFKapKf1P+XKlf
sMCt7735NZweoBli7OxUGUcBUJRfrhlM8kJrq69KM1VF1znNhufzAi3CWDDEHmuv
2Y6rx+5npjzpZhe48exMkMRSdrvTIsp5A8Y37suDjjirol0p0uyoOyhypmXWsLTz
Y+VgEZB05UnYL3+9mXksizxN2PkAYjkwEeAXLwXeM+mqLk7I84fQe0wegGI7dB8Y
f3XvEfqBLzbn94D//X4vruQzptHDeixiPkQueyNUWzFr1Gu/RBkIJuBAxR2plSNH
i0WtVlsIzm75DOlHYN80H0+hX+iu1sF+ereI18CVT1+MXK9Dz6/0pSVcmiM48RbG
OlqezMYP9pcTut4MEGVSQnXucUMXpjNkJfIrjNpPo7satXyj60zz6cI8vLWRXVKS
cUGXEZHqm0c//xMwqDHgRl2VpM3vAlrBTPtkuOaB5DK9dVWW2N2dVmM6WEIIvCfx
lRy/eBn93tyDJVcpds2ZsC4siw7uXFAmVZMaBHR5mnr2YyUd98SVSLpMvV+Eja97
vPg5F/GvXOYeruq9KnHAeJwMZwE3aK7e57RVyImVo2dyAivyZ+QFc4XjWLuMttLH
JtgKOLe4mTx1Sf+s2RW7/6VxRkNihCc3pwW2Hw05XOxgbjrGco2/FHpKzci8Lfsd
JMFRwksihNpqGjMhm3dxSXs+0QzmhQzjqCQawMPMs7MZAZshrPZ6m1RwKgxe6Q8N
SEfaADCwO0E7/FEnWJq/dt0bs87yJQ2JAAGU5EfGyEw1rCyaualDNqJTfTpz8ADd
YiG7l+qek5GXzrVEZxC4VCp75L0H3Kes4py6hbBd8RDezK6Wcw8OnwCy1DlUIWR1
6WLoQ/9gENBmcV6o8DtxCUQB3J1ODnw9CWtfSKoxm89rUr6eNH3oh21ZaNkCFFhb
xs/YBLnQbcMKV1B0U9qMnU9HWdiHdmiMblo1MLYR5kvzB8UeBw1qf3TV7jm6AAyq
GKfI9beKn+XbY8/MzkvpgFsYFlE6mOtFua7/UcpEZFciOmNn/GRgPjGYF+TNN6gl
BFQc5yzzSV6njD5Va1G1duZc40Oz3QF8pWZ1wA+eVmv9r/1HTwTPkuQ438xEQovw
JIC/ieW82PQYyrgpRm51r0GVc3R1etW/ruQbto3Y58QSyJSLRrzXv9lgw4mrNteO
LItjKuQAhGyAYPTj56jQCrz5FCaBCMh/6s0hXMyzOHKe8u+ar8bAQh08NkO6mhMn
xB8STq1Esng0eLxcfX30i30YwbUFFdArvcJmRMne8JB0PKm1YPwOx4c5M0gni0qE
2kx5xjI/1PWp1WbgLQ6F1wCBkdglyQjMkZ78pvKCSG//Ob8KNsXPCAqJA0xXAY9L
bLVxsPpDAmX1Rhkyt3+pWmhEV80SkaPPxIcZaX3ZEXabdapGgM1vcxiouKmF31qw
PEh0QSVBFXpr22rtvLRxtskEDAT9R99R5zDclNLMHFjzqYhyUcKbMZcgWqIdjk59
Nw/r45pHX3CPq5XNB1p40kaq+GFAPb8+u4KSNtA5ynxH1FzdjCybvj2S7hllerbw
iwfSZ/iCmn+tjrvibg7R/Q4H8AeLODY4ovRrF3NpEe5Z2Vyjrxxu3ycaD+AfjodF
0dNYEWNHU86Z+Eyyf2DT/X4OSPdfcuQiyT0hw4qEcSP+/X47qz4CWdJRyXqOnla8
YkqD/ycR4f3N1FGrPwEC23Nb7jap0FheMQVonxNvHLc+Jr8VsIv3iPXIDnUWFdwY
rSDTLK93gLXoPmuD239HcjlaA2ZD049A42/YH8pbgfiohB/tx1TttTgVqPjnQSOP
lCHhJxhlBIkp1XTOl42XXcH34gvxfApsnJniHBok6C04kjfPR4GkMC9uoeuFnutG
iGDzQb9TIAVwjDyyy8G5Ig5lbG/Zy1bjt6ow8IlPJcz4cxqfCnx/fPCVyLDSm9dl
0FvkzaX3YvLJm4IrHFeNKw/6QvX671OBv6OE0j+dQfbEM8/gT2bh0yTnCSAYCVdC
s0CriVpOx23DZzdhwXttMQfiw7CEN1NHx4XwRhYZRAME69zl1SisRnP3/ptw9s7d
pyRHklGoG7YunD0Ot3t6Jkp5B5ojKbvwn+kqY7vlTFc6e+K/S9ZPZswlVORBDDRn
XRK8RutHlc8DQiuwH3y/HPU88wu4NQkOQPCsHfY2BRccqHA1aXejLnDdcwcrAYAg
VZ4MWW/YnRPdCxOwQd2Q6SOCvgHT/jXWKBpvBgq9TPkl54PsgXwJ8mgyAomTTjGL
jXi/O7fGP5MEBZXJzqF6KmQC5J/Yb+9U5tAfZkDcTK7fJ09xW4Y8zxy/kUWOUwlC
/hGlv83RyI3YUV2BIAUtMfRl0WrOGiZ7zHh5W8YBFKwf9Eh2S9lpbqlU8y8CXVoy
P+2PLJIERrFAYslvbfkBIbNiYxqspYoEkLza1RLJy8d9pY9g6H3moVjY63lMLS+K
8TzaDVf37MgI6VpRYZd6RQgpLwRVpeEUi1v51auAXOjgLB7x6jRhCcIqCo0g+NgD
a7jI7U3RwFAGlptzN1X2vwQqtY2f5a2atUWizd/V6WD7YnXokiPg+p1gSE8MjC9A
SDE/SWKlQ1xtwf/BUYAe4WPCBZtU2+Sn4BFYT+S/EBt7jGg8kv1tQ5GiNAWYoLga
7+IrCTaw/c0PUTTGDv0iVF0vgWznTYADhZmpcfn3RnTOIyEwCP8F6im0A+m+A2lF
ANsu+q1F+GeJWrDYsjx2hxymISgLcL5xqAq1E/+XY8WK9zopHNOGxHh47tv3JUde
jrbWENqcrLTNnHk7hvYWUQt9gKoEf4x1ZEPnOICgrPuAsfiPAhUbT1EBcA2lzp+M
7rsZtGHYKN3GOHPFqMNjk4xfUAqe3mUPDxxv2pVzXXXqjLV9rQu6S4pCl2pGGpHf
zcV5evTBbaqu5qzXr4JCw06EH00XC+j9ytDtzqlenhY09CylU9u0IOeKG/T7/8zm
+7TSI/FrT6qhbruivVGzbsXO6JfuHAIWUjw5Y1bHDe7QHpGTC70h5vPYki2KuzD8
bsNj67czcjSVDUkf2LCDkhH9V+97c4L4tAu9+SAR/9fe6SHkxu8lMw6vyLbiIftP
e7Ru0B+pLSfQ+YK0IfQABvHev+0435uAHSEkunUsABh+Vy24WrX6x1KZ60mKiZZZ
whTnKurMbmCBIvivvNyy3Pqy79QF2a/CGU1OJVyII45Hcpqre0v3hCI0qmkqZMmQ
0yDNXmCkqZnTld3qXLuxhtGPE5D55vfj8xj0064K+R41P6QkNJfvpy0Tjqpy/Ogd
rJvTgceDZggxki5mf6DPTA/hQJa1v+TWvxu+F8nwN+WPEk1+sgohQ5xEs7uqC6Hp
eU3RQR48Y8fgc1IUUWffb9cmFl9tkdO9ZyO6i6dz+hCN8fHL6ED2LXAf/L1KSmmN
YcXTY4mriIMP3KHmImWbhVsHZD4rC3+fa1v1YV0Q1yo0gcVmZH8B0Ac0gC3zY9+1
+dyKhKy73Ho5g9+lyHVUGg0esuCLyi4Q2qDgogVmP+WgpbEWMMaGG77+dBcXOGMz
Me1wQzmwZtDGkZdPFcESEVOT2USWSBcXbKgse6AeVb9Se71QjG5VbVwczeTk2HIX
meliSvZ1uA3C5FBHRlL6oWMCGv01R1uQ2SWUkMpioiiAohUtb/7F34oIzOD30tzG
qm7eNC1LXpy/ARa55BJgXYVEcx7RvozhbSD918BzybgwI+QxxXWRchLkQFeQqdCD
Q0k2nl3yCjcuBfyuYHs4ozirBcYvWUFn/VKVRx7B3liyvBQFzxlOJSRgPUaJeWvo
UPIWlenFBR6GOBwSP0h1rJrBAWZ66+p4sk+qS53soyMdEPs0nf6hU6RkJAGcwVFD
iorrc0QDWtRVzBE42b26CKiEZkD9CTAuel3/UhM0Sq3g942V+NA9bXk4MuqIsmNq
TEoBCgBNC7LJrd8DaYyH+KErIHs2lR6bgppCqG+OpgcCWMlB9nEy7IG0+eVvzClR
jg+qlkdCVlkKG+GFrTIcoIDB1wzIsDBTC4RAsrJurF8PK++kvePy5MD8tXTYPCL2
2OdGEOTP+GgkYiuKVo6jV+8ppR8aLmuWiUbcAys0yZaaXErbb5E1DBQBYYnAhRR+
AsdTMWFCHicAKT0iO3tnryrmjUJ1lA+kKT6ozL1vYcbVbcISem3QBb3Rf/itWVok
3QvJVwp7egBnBu1Mj8KU3RhMjNEe6noaX0RLXn2j8/27/r0l9Z+Ge5I8YQwzKcMK
RRHVataZrn6/pgSBQgevO97FiLUuJH1YXvTJQLUVvb6NDcGmi15aKRLFhKUBo+yo
WHZixYtd4o/YdlIsItoFfFykGUmV5lOujDEn16KwjjgXCNC1TqQZ1C+IjBC12Q02
pUfdiKjrEtT2b4vnx/96nI2fgY8wtdhDJ7SnfblvLXfACeOIOdpxmfyiC23y8+4w
Cjc7oM0w26UW9c9NEY18rI3Xl6V6uXoA5AfJdClSR6gGuraU6nUvk0mhO7EFls/M
gHDmkhu7mEb3RKuWYk2dgngEDnY3IPyRf7z1Caejboqr59mGlQf75T1hkMaeDxqS
u6RxZvqFqoAaQluEePgKXi/35PgGZxhpje1yw90pw/E1nDK8tEXY+vuGqAjEp3Gw
1hoE/UNSa233+GZyo0d0zS+kNmVPmvpw+ErtfP+KWOwZ5HFnKkBNEQb0KF92d+dd
lUyc4exIbItcAestD+zfMrPAPxnjKXBnT1PluP6Lx3/N96Ex5YSUWF+Bmc8I5ZfF
brZ6LHfVQROD1M72r+2wJ7GrFSE2iNiIZK+wi6Q20cCwRK8ZPapCYLqw2rYTaB2C
au4ooGbJ2KCTvV/vA12x/AiApvxvaVQ4y9iUToVVuyspCH3BjJIgdGAo3eMuBntq
7C9Vm8rB1BFD8ZnANOzEb8rPpi5s3LT1mi2CS/Yd89Cjwlh7PvuXX568fpPUa2xW
aOMyVqDEpQfjsRYsSygkcKeXjPZtOrKkkATyQ2N3UjqhX18HYrKEmvvzr993/gOB
Q7DfyeC2V8lRqhhF029pOpqRqfAhm/1wwY/13zPv7wFavzD542+2XiDioS20r9xr
iKG+Svq6qI9A25ymc5x5NPHneo/C8uk6fRzdpsFzFlQNAcp8U2MYqZk2tptdMz+O
V87XkcgjeD0bUKwc2NkZw4L+yZx1X/juWr1kBs1ZbnNxf1i+oKj9j2sS7IJ0GCDc
zHu3xkGdiNSGNDuRgiobT87pmeA6a7ASJIs50A+iaqMN5AM0wj6lVA34+iJ9THB8
07U159H6wrY/neSpZbJac3PMVKwJnJrg0NIPrYlPpPHIz/j1GxMAfDrab8vcojJy
WGYnJwyoN+qhUcJs92QlivMArM87MrGq7LeidzgRhCNlGWlG2zcrz9r18STCqPtM
zxHYzNgUIhLYkrgtklmm4xiK2zXWl+6YWq8cvaPLvu4t5zD7PBZsZ4uNB9t2fBRE
nUeNWtn3fyIvIiW8pD+BuJZ+ZKCJhRGMk7pb8p9XLlI4zWBieCHl1uPJ1TCWqOOw
o+vx3LZlqf95OWKLQ8SSsO9XvMrtKU5FNa015/wg9qnmUZqkyc95cFKd1IbSdci0
rHtJyKQgQ4zUthB/Ws5sxCTNmagJBYCVd2a2T723jePP3pe8BhepM4mGMpLlJcX7
rarZVPgTwpTO+zMK0EbPSM44Pdg7h+EnD/MIW481woBjx0E/x7Pyfy5gEDPRDcIo
+R9q2Iet4CXsUsrcdOYh0g4CaT9fOQPnAHxS+Ut1IpEu45HEpTEkE+p28sf8Dgze
afEev+5vZVipBZSy8GaRPySFLddaPcP3tsv2q5D7ANKeAxUiyRF0xO5MEL+jsDdJ
lcCAzyYZpZzA6DhG4hNCqrI4Eof1wjKJ8zSURtGpmpSb3B79VrjsxaF81oWdtsCp
I+ruyXUK+77wg57klmldfyHT3EHSmQ99dUQWYV6JdVibVYE/GbujrirS8NPqlDW9
H02pEXSFzuUOF4oNbxKumo2gjzsNjqQKfUYLL6Toi0VcneoW2STJmbDwC5A9VtJ0
Ao9KEiBv/+w+KHknc/Y8qvuj0uozmYO59g+Q3QFWSeFZHEh3bw+uQQXS7lCt7WeA
86FLwIELcoUn7CjrgnnILdePwM6cR7B1gEfpIYVEL/Zd35mKq3xzI3ILsNN5Y9x6
MtfGAtmkaV2g76inu4f25uBbeCHAQYGl1dyUXfxjTw3zilCNfmeHpDW0vkhGWfOQ
YLSPJfedbzgToOw2WzY9KJHdZj9Z6paN7L3r6BmOoeooNAWIuEMYoQRsbyw9DyNB
Cehc0ACcRP5I0AhCMPDNVdiycGwiWYNmrPum2xCWzpGOXw8EMQV8budydTmmuyn6
OQX/Cz5hdsuMBNfP3PZhwuH3HS0Lza4Uf2HmTBd/opScWXyblWQewM0dFO4nxGxc
UZ+hTGiqH3Fv5yqL/zA0kBZAqyv1ucqhNqkRbfNlJdEL7fySN6kyr4RB4lFjMjCH
hPDOC1NhY+se1p4EIpXIzPl0sJZfd8zhqNjO2VJob+ORg7CWbPcTdqot1/qm3jYz
tbMCDYTL6ihHBYD4VSNrX0wqRVBkldmUTofIeiCMFgAb1zFjRbd/HN19NcY4ATHw
RazrBF9R0H1wbsc9ZcdohEXn1g05F7lQ2A9xz35HPElmIox8coWCltsdGv0aXbfl
fzl1/wPz1xgbIv0k10wKnO+Ftr7UuH3v6P94T8gxsPcK0eK0vBRB/yzG60UfHgfj
MF5+rQ/f6xLlTAosupqn2paqYMFnXd+rqujBKKasMy4+f5QFty81SEWzPPlshYJ9
/eRNsTrziD26X9lsyEV5c9dAIhndoryAQpDxJKk7RenT5TzBxi+F4OBPPWDBytJA
b0qGkFHCfEx5TIJ4OQ5orXCsubJ8+44MLOyWs1XVRmLo+8SVE+I+kAizHQOZ7IDB
i5dHtqGFT4ApQ0I8kD9i8a7BsFctvgjquKZPqtGeIevbALmYrnTduBfMV1K7rKoN
+OAHSMT9/JLeXVYilxbTy+Mh0P2U1m2BF/evqfJEChUMUXypJM3+39Of4kGPqg1g
hN2TIRLqQaMMfZxxHktlh3hW1FrriUmWUrml03pY0WoSZkJ1axUPHQGXnaoCgwu2
b7/t30myhw8MdsT6ZcVVHF7C+VsBeHI4cxJalkb8NOBKbI+uHMUy9OlBmmghptn+
COdwyJ1UL6rqmV7PyE6RfwtFq4QvkaSTzIsrNp+wQBGmFDadd6XlN4WtsnmFXD5X
OlBBBUN8/Un6bR3fv7Z6CCrwPQQmLrdQf6JEcF8M9UyAJiylu97x1lFVQK2FL2yB
Q1V6wbaq4ps8OpYrC8novKXVoJpqvtNz7n4mQROUfW58dKvnUNH+jistiMK66iRw
K7BH2j5OfCW5tRB4U40gcCBah+pc7ofCctap8uKyap6//X/IZYTrgy2dSL7w9bYz
NsvoFZDVUHNaoNvpEwIqVboZLSTOZx+gYOjiVN8A+vroAk0+HBm+oqL8nZ8WBIOR
GLdjcJrnhkPyGMbukF8HQeA0fL6BbBVIAoCAoqAwDiyO0sxkQmDoEYPEQ/d1rc44
J4sqImhNYTlYLMI44Z0aO4k68if9ezEhR0TAg1JX/KU9ls0m8N5liu9mIC/+A6/7
Fzu/VpK4N13cil+vSrd0H0tQmQuIFvXHHO5JiXWz+9OUPLWo5YEP3OoxHkVW2O0W
FlnLzygXseG3+PDI51OeP0JeFUgpOQu37WtwhAKRjo0slqOCuvsGqEv+GxaKwbbZ
EW0qbkpPyu7z7AVdHSeiIN8fTUbuP5IhWPGwv+9eCpyUoL8QM3Nz7YAJyM9d4fih
aD3ZBK89VVIW5Vzz5fBr5+Vd6bBd0jBPhFPRygzybQV9XjiWXAIyWPRmWLoMTjAH
UqLVCeTaKx/AJ8Reh5/qRZNyaFigf0SnSKqI150HbcQz/nhL3wco0mjtZETOZPML
nk5VR4dAlsCudaGRBkgOZEwfvLTToBoCeuPJnAjWgd3cqHV6K6VHYvyoJXVDIJ0k
u4FjEk5G8pChUq49q7qufMHbB3agwv1PV5Ma5yZOWWcIVUmFGL7hwmcqN1uejCiV
d+AzQURlJDSCT48hesEvtNc6ydApyPHtLRRWi/5kj+3Fz93EbCG3IJCyZZg4zehj
ELhO6bLKUX7mZ5kq0gXLn1FzsfU5nj6nrJ2ogF8PdWCsTUCGXDRbf0JqCmlmgtu7
GDeZ2y/Nd/u6bGLHET0KYit9NUTsjQE7YxAp7ht5Iyy+7ENZq/mE9UX5yTHG0N51
hTBybd+I7G/HqvueUbT883k2cUTbSLPvj5CGltifqMlLl2UWrqh43LguL702qglx
H/9SHwLtwi/68mtObHwnh49GAn4P3ZMwicUpFivEPveXrR7alwVXUKJQLT+WqfA5
gGvhvSLOXm2VvZKFxzXneAYs2WIkxyhW9Oc4VH3wQIslAtFtX6p4MSGYqHcW09Mb
f86Nt2cb93CnBXQXwB9/KMG1/Y4WVdZmyOl/PD8RO2+weyeY6dFoXICf+H547Pum
QZLwL5TV1eJZMtU3f8mHXggrjX1pAD8/EjWq/9OzQ7UmPmKM6qPZ6MomLNjOW+5G
btQ/XS5ipfpN7KLaf3wOaGgkn0/RUh3G87K4gT+t4F7LP5nMa8hFd7BosbwBgnK4
l9uY/gho9aWXzhKUMSDvGy63IQS4BnRRmv6Zv1FwcwrnEl+ObsvAJZrB2HaMIeKg
Rc82f9IvyPkAhkNAXEuPKIP143y8EjtxYACWTQiHe1qUoxZuX4J2E7SgSEO/HRlI
Ljse0L4ybJuKhCG4sv2eBPDEtFiXQLrxkeNM+FqlQEVjAzQCmBsyi5bQLCh+gc8b
sr0dJkshFzeR46iGClm7XKVzyGlHlsrEIW2M4fxRcwG5Kuv7nnFthkOeI+/I3Knk
UyVodBiccz0ujlppvM/fpm+GI5UTu5Me+wvZrkyJ0MukpgKAncpt5HsET91JUyKI
i9ZinX/b4gpx/q05VVPN1FfiIneb7tzUWQ/1W6D057dg1OEE/8Fa5VJmR3xDIePk
6db5vjXDnhjFtGf9egYdzojHRl2Rj7uAHhA3O6l04xBwvYufIVLnYrrZpaeM+6g2
i2FVFvrhasIpIoj/obixpgio0Xt3P+mJeQFIdZCCGzH4LzxfK7u+m8Y5L4e7C6fZ
hgLJgNhFdx+/mTjvz6anXbR539S0dSdGvUVSO02y3POdrmlVaLd9ca1yrkzW/dtS
ZnKFXPy3BYlVjBtvAiw5no0B+UDzoWG2/Z7ZaYPx82QKyK+VWVurx+9Uo7bgSjq5
0AFoin+s9prIju9G1kZ4kFKR6y1oOGfc8u5WVNhU5UHbhMZDJrJD0vYUTwK5LrbT
/0Ex0lV3tnH+pLsJnf6DgVAiuh8AI9XyMk0cSEGWXWs2VqeU8lpFVBLLh9slbc6B
Tiy9BG32x/BrGe6iui9j6V3kcq27+qBqwkCy9NTiKub3b9t4Fo18Um99GQiUe3ai
x+rL4cnrY3JUC3+Y0FTDkhd8yxc2Lzn6ecm7BlctVDwnMfe4UPo68GDqg9GQfM7X
cC/W2Q94bMFFB0eZrlNg45a7JS8/tlwJqiV9uwg0IdSybSurBXDZzU370OHczy3k
CYqCCTPWh/8KDkosilQCTwpXLbQw1vEgL5SRksCikkFhjW2f9KkfvEEjI7wIy7ES
0o8QTlObymVsPux2KClcBK/F1szF1dnPgJASRceUtOoXOwvVDJegu6OQXK+XKsnb
veZel8PcQoKo0EIkPwaTZxi/xgnJNlECWi5v/PQ8XmDadh5BzKamJymqWAPb1oR+
LNKR7n52TZT1RY/iXdMXtx8VSx+F5bFrLz0HL8H2NHK7Lt7XfCh6L8oxdMaS45Tt
pQxScD41rZYOMF1xseS/3NWaGiYe2duXumsQtzRQdy/0ygN2lwx1mXldsJqkmRaB
lvLn2X8NFjJZbwHzLhuTEQVLbvoFYnxZYPfzvDlI6G+Dy9tVyuNJyrJ1gKMKz9q2
f7mBgRWZl3aG6IalHoPT/PeTSF1w6uIPfp9rY+4D8uIZhimBAqViIFV3lrNa11UA
t7NfOmo7FKU/YMZfW8I/7fMaoAdR96UHCYm5O8SRfkTCgSjdnGhJBZYSurLDqun2
ZIWtoc+AC8cxdDfk918NGwRms8Fx1deqBg4bYyhT7o98hhEfILVCrsg7REqWXWqi
4mz9nxXV7oaFdwrygYWGXcA+nzW3/Dv9csuMgjx9bvP2kuZjUZMVWsEL3PThxTS0
0lZQP6T4AZ5vNuGYGOkOZABz3UkmE0/WS5OteqCIgOVOkb6Pf4QZu27iVRwzCjSX
YRVjZl+tKCNKn2sZnfzCpvjU23pGbWacitFNEB8wLPaQzuv7BVS0CKYMYzYYypUR
/CtUUqLw3uaizyQRoeU+L5SVqzcqHIMMKoCX+K/kQG1K6iN3FiZh8uapxSEDD6NN
o7LDdjsiTl15LBCGyq0VQI/vra9rsAr4RsfmY0B8+ihlymLv87Rd1dmJb2lh5Ouo
00kjG3hFnJdFjLE+A6E5a6zZyzITBLnHbBmqY/FejafEDgLZjtlmeL6Clpi7zNwd
n4djHkvYv7MY2XRIcbc7pbvTnbDM7vBWhIPlHmyMvZJ1ShU4rejoiiW1ZHQfGajo
K3yXFPcIfQycHwe/54xUYpGEno1ZGuQ2hC6RbEVJ4+SGQf8jnp58YzA3szdnwMLJ
y5WiJn5JFsd3yrgDR+ZaCBa6z0E9HuEEhKoeHImlx042nzU2omKyRPFho+rOysHt
D0+fRwED+xL1UOUwjSDBR5xWh2tIQYZuOn/ulStSRoXFynQu+ZpDCmOJs/xjwtPJ
5FAxwA8TKleINq466iB29r65P3oDTqCrYAiypogQSK6zJQwiUA5L7JnulrToODrz
3ztP1hvdlDW8QwzRb97mKLjmp4JY/CLqooDVGUeoXXwzwFXDLnE1hrcnzHklhJpG
N7xnozaoVa7oy2zWc0s/cXDI8hQBpPllvh7x3UgOMPMSz6JFSGzyZbWxgwL3PFG6
HkFSKyr7w9RMr4wZWMwBmTfHc0BdSO1sPfhBrHyE51+jkZcMjGbc4zlbAwu/AG9m
zVoOdE0H1ECOmwrap5Zy0VGvvJt0ES1rtE3JuhqMgWvwSM/Lde5wFe5Uu8mdqy2y
hU/Jhu1cWNL1BL47HKIGznwRa6biXUXdyhWEZwhB20NlQHSecWRov7OStRzgJ2tS
eOLjUBIOUoOe+6KsiIjlvwEqKvXurj7SMdvIbfCFWby04xFWqZXULiP3PPJoYIs/
oIilGJs/1y/3AnpNqV6Z3rtO0eeANcO6+9xLPw1qXsTAmuOoJUpQmVia/0gkBHnt
g/tbH6h1/SCotcMd6fCZG8kshlJa1ALPFXVAB0dnCZBpPTy/h7cUsKQg4zFYI2mH
Bnw2Ki8OCwSTo0qrgAO8G06b+VJs7KINWRvmObCNwfyel4TqAqHJnQfEhsr35vWQ
RFnn46kMTdOoCazfsEE3UIwjECJZ5UzaZsM618fur50C9tzS6IIwGSeLdr0joYlV
YEJ5XaGvsqZxBZSo3Sfaubt+BdJMGAwBhj+MMu6LcFIAeZ+7f3wwtmTrsYkPCisu
PtmH+WmAkRjItIWEqpksQqIPHRh73ZboGUdf+jvyLB2SjCksRgd4D9dWIMOydLET
TACu0faE+dwuIpYPZwms/yktQtfh01k8dy0lCt2VCEN6khWcFWw82D0GeBAT6FP7
DDA7A4jIb6pLO2X9D9tFy+LB5HjjnD1OWWivotJNdRyQ6x+JWVOGRQwsmL2Ve3wE
DcpCbxcLFZy2khYg3D19n9Ngqydju9K6QvxTX1yKAAzD4bYRSYCZ2hTSB90ks4o3
lxBVUvxSDXFBhhsOYRIe0zLOMuQPWfRm85bTA6mBZKTyw1vI0KDyeonhbfiu1kN8
zJL5r5nFS3P/QmATGmOmVq6pkbv+Huy4S03jVbjP7Y8uAsu0yFjAcZlB27EtGcIy
jMZXEmS043kYTwyQzzylWFxJbU0I1y39H8MAXgNl7GbQvyHx+4wVVAkdUMHK4AvS
hRpWEg4zncFddipJFUtAfMF6+a6nwkBagU2Pd85SIN2kgqm3ENwImokQNmsa3XYy
Sxn/CqnrRGAOhbh0n3U/ZrTH8Qz8tLYzaPZLvjLBqJ3+Veh6WU9cSw3cmOBxuaHE
5yGNtmlUmzR1fvj5lMUwIO2kcAvcEifQkBPRZ1hUhL5cmOO9TlInTy0VanBLyp1X
z2XIM3MJJ8Ba//U/8/InCZFyGi0Z3Bmv/h+sgxf6AbW1Ll5B4PjyKvUfBeVnjkhN
LmleILZrc9d/io6N2X25Tp6JlkQx3F3wSpqDQVJ5TCZRMvOzoJ7eQmXZDJHzGDfZ
PuCyaANo0WTTKo2mFJ42yTkwt6pGChDrqCNbAnGOHvLdEuSOKMnrRaKAQ52T4oYA
TwfdlNv2AEpHUyib7A7tBdkjwdYseIOvUclgH6TS2M2FfS56XJ1oqypoZyJKKW8v
JqS01tbjkcqxLbWC/tgn0kvIjy4Cy1j8NUi9uU9WzzggAz9PgzwwYiucueaVhiX6
DoUY9Oq8TrnmZ1HPlzc3Ip4dydzHBhJ7bXWihyaFrmaMO/WyunETv7zBqmTobs1e
Dvt7Idm4Av8MNW4wfz412x+Er1+TX8M0eBs9pd7GrJx2WK9DXW/m6Sda1UN4ZxTk
fTwrrHY9X2om9cKcYQ2y/pkShwEUCnkzUjArobxY33TPIUz3qIjqIT9BfpoZzAfG
784btzCxgjyD10hzmem9rcJUPc3rbN154WWWn5vbv8QlsWsOy373qKIcozv68/FS
9xA09y7gOWiFlamKIHOVPfb+ikDgyz+1LQtM6HdWkErC1PH1DGz2NzLdEUGrGQBi
B6/OT8xiUDRla6m1UfO984eXO1v4/V7M3OrwaeRsPTv/olUirA57O7S7PEHS7lXP
SeF9Kyt2JwRrzUoq1wjKowIvNATDIxq45eUaVhcA+VZk3DC58F6+fmqGCq+z2VEK
faj97P2pW7gwrTdRFRdZDSKECC9H3NdrjaV7Y/XCYj6/nNy62/ZCmc6AzO4KvA8L
lrNtlu0HaEgLTdDA9OFIVtIIt7cVg1w1MUAH+rjuE9+B/iIQgGnmeLlYpFZVr880
bmpMuv02lF70fBfQzM68eP/DPWjVJ7gHE6AyquSyrTJ2u0Hb8LlkMm5d2QqkG3gd
x1/go8F//gojJA9rh3lxZVHz33ga7OQw1Ac6LkMdDe4f8VkfgjJfrE7wFTXkIWN2
gqu303Gw5cLvaM+2g2lUPH5tBpsKkXCssTIFITlxQAKzFTkmcF3kH3rjr/D8b4QI
OWjzZkpHWxdlytrU9ceQnj+ZSp2SDO4pj5o2w8PRAP3eUchvtcgqm4jxlOu0FyKe
a5wKEgi5VBEbxcrhp+j0Dwix/ueBGVV2nmHDJrHiebxJcaURUZ59u18SpFTNM1VS
E2Slw6P8b4hc+eLEhK8e1LoOiTxUtzQGedgwQtMd3iIjcZMk0L26zuTJ0SFKJw0f
tL1LjxW4DC/WmmZSpTXM5/wfBrexakTXeNeebMgXUtdBCECUYm/gRJh0A1hcsycW
7jOWoVQSTVyeRI4HvhMfnlOZ+7IqbVL924idS5zDSGR8mkbl/4VYmYOljH0PpC3B
wYA0YHr5fBvBu8GUI6uHp/Xk2faisVCcqVrA/2p6xsZHeFDTm3v08ix3Rsh5HF5B
237FAptTMwwd0M05dnwojy+pSzR7ARR35Dd+bDtFZtU3KFFB3Mjb11o0x4uPD4Ow
mEAuPWtFNt0embP4hLFAqAM8gcDcN1KxDk2sF5N/XN3RJ7LNKLkgWgAE+JCYzu41
7acQq01M2YCv/JBkyBVBVs407ZOP5HTKK0AkF+yVykVLwHpxQTvNEeO7wQVzbQwg
3JiYOoyjWpD5nufBxR3yKJwqQedET5ybVoWWaXj6vOhk5D0UpXCb4rGVHVU13jUj
W3ryCTsXtnCx7L5dLCbxHmP3VmiubYa1RWgllDFzGJFSeTQuMWmhd4HHXw05VgK0
NCZQi/5iOg/ZrAqBOX25Byk4WI4aN39LRpHljzA6TEDKzsUv6YMgLv0ImaGEcWv6
t3cvFL3ctBRNqXe2NIr3Mz28LejlA9hInlmnMl48jr0D2q0CdxEIay0qMyx7nICP
V3dRIwYs7VN+Y8pKhECHQm2QwqOT5dzGNBuU0g1IcuKT9/0HEqYUqeXsxVw4n4hW
8DL9caIuBpQjbacsPpZbqW/Hi2eERqA9SobG82nKvIqfxzlfjqCldHyV/KykdvXe
mwVoq6MGeMrC6hyoAJ8uD1Wp859BPtVsR+JCs+LiqUBfuLM+FQ9j6fFTYGrbUMK/
lD5jRT49teWI9OQE+hMM0cytzh4IqZWoP/l3Jvozo7AEPrjctkPMHPw28sEeTGGp
DOrW+oiWSJeHvsKarvJARcVI5Ip/146K+53/typzE9ryqWzRvNn6PepTbSLE/Vqy
vscSG3ookMeDQACqwo7r0lRkwTqwOgVqYZSj7P3ECmT5D53+d44fXd3yNrJHTMYk
tG3wSaJjtjcKxPOEdWNC3ymt0pWUsXXPCzaigzMQRJyfHEu5Upj94W+I/ZrHfya0
epzz0s8lZn+DAuXHfDr2msnCTnC5Q9MVIKZtFzemLlrT/CAsmyyh96pJMDHcTrVg
ah/dZ1EtIwFN6NpsgRBm0K8Z22z8i2azjShKL4Bpe09pAEL1nMsX9RvcQP/svC+u
w0+jmGYUfSBl+ZHWBNp6AF4W2hRLEIpiK8aX7C6/KrG+myEWkkXpnIKnB7L2vRFd
zM7TomTuuOzM6/2oN3/d9dyPaWGSVK+VAAHYEFU9sYcx/j5ppT6+XUe+HwfYCDOk
FGZHmtRnt3ivD556RR7lJVPGeDS6LgjUe1EOw/Jgo4/oDUpoQF4XMJSxVBPS8LQl
2/JqCYOe7pdQC5gNMHW7iW7DifFHbxxzabc948B8hjlLqO+c81JedUA4+BwSx1TL
h7NFi3Og0kdKHGc5RjkfJSUz+KAdSQ2bu9UDIbuSJmint3c+Oi3TB63i6b1We8Ta
K5E+Jwk/7by7ut3R29klwYKNdZYFogv8oPEyeUgm14yfqkYR0Z65w5FSwCZm09ka
SaL0YLJInE/+Qb9/hPECHbyVstB2VUhzBOtQunKKAFssrmpPPVYL/NHTsd/skdyE
0ntnL3AdSL9/djvSh7PPXClJ/P1nx+jgCoLG1+mS2pR7AmMrBK1TAfyHkZfX9b8j
OrFjSjB3b1VU9uN0mwL2x1nasftz5vhcP2t41EFlGWitzXynJWxC3g2DWFgBDIbP
lp4sFvlIEltYxkV/wgfDWrDVgQvfHIoXm7gDjgM6Tl8jmKVNaUqXNLLQM9loRAFi
lHUSShQIG/hSptWRs904PRvzkg3qcnob/sifOsEmULFP7vVfaoElTDNVbiKTosOr
3atiDrRZ588BnljQK4FkdhzycxsPDFzZUgiO0NPUlU4sJ+FzoDcbIsdp0ALqeDAk
3milaDpImHf6hEtByWo3+QjJY/C8mO2CW0wZiEyyOeKGKjmIP6rc5r+aIPfCZ/WV
CK+RPsogJ1FqDRkWgpmnYE0BAY9gFZQz9QRwEFb4hMUgiVEOywjuiRfSA6Uqy0rL
vvBUf8LK044zZnas6uM6yirp7AydkJx/8HdFuZPWjilqyy97gNYO+XKqA+mYpVVG
1UDIcphw/l1BUu3Cs0NMHcPsAfoAeCLqG+rKE0ZgFHCGR8WMywIxWxfkjYiqE7PC
LN20tgaGzIa92SBLta+lxsyk7sQ2wEVIVs6Tk9yA5E9BhAwQ5Rlirrlpw36kPUGv
KU3CqyqmgAnrUQRV+wrRSEWgNAec3LtgQCeDMFzjSBJNVH8GKIJ24yieO8Hah8c3
Whgg8o2+Nvg4k2rJ5plwKDcKRRtEODkzt4MYyAtR8V3CtAzPVZzW6x/Nyu92UOO+
Ym5UnbCNLPWlugGcl1oIi1tjoTXDElBLPWqTwa5lZwtUO/Zv17un6DPhlTrcdiKi
kYSTtgbZbJai3k/HlL85ckVa0ZQWrXNbHTH9Q3lJ9HEmoOGvqaHCXk74VeBQZf25
L94dXupJBtuqSFPEB7b4ZQXTF/7NVu5Jc9VLDPCc/T7qK79qRB1m6P3dpjntZCv+
xQYvC2edC5kA+QLCC7afGerK3eJG09CY0qMOQhnkt0IOEo5UeS8nEZUh4mmE1miP
vlmrQDIWGtVvgv4ZBOnPIDH0egDTnMHrFj9INTMJ/ARLFUkq7lKNukJD7K3JalD5
aqkuDs8hhwn+vFSxF9lUiCkBLFTrrhPRcgcKqvBGH7jWh2RTTwZXungegC7b1OIG
AJ+UHsEwn2HCCzNtbdxi2crqwJLz0PQQ3NsN79rjaJHwoWZnJpOeS8uX66pG0lLS
hvVB30BsnT/EUUzM7U+dJ35HOZfY9KZHgaYzrsltzuYihEAD7enGQjUyAxYzyf1o
7eEkX7UCAeagoKm4LqsWnoI9p+AAZIL00qa0iPxbuEaMIg+EovTvNgWjjZjjlrCn
djsAtDiX7hh9AIY7FV/1829jRvBqn1xMWqSyc886zEMp/yxCwQCzCcnpdE9oszRP
i4JzbYqxL7feHRiX9C7sqn4oaueYTRtChLzAhdH5zs8eiyrSvXyNwSAIZeObItZv
xknMXCO6eHm41931lSHpGNM30xNoFTiartddxzdECmPXoDfThTMonrQVrtU8jr9B
dDI2+j+p/snlaBBkaDpOrwn0D9TaZEZHNc/t/KAcWFcWngYZvVHyBo8Owo7ZOHEQ
kBnt9N087wmJ88QvvX1qgWyXIy7c0vdsJx+7Mxt5J3QFAIH9fmaDEV2If5rrDedO
jf3vAewxG73F+QG+8sv6omoSyhCGPqY1DjBmJXwsNraXCvfcZGaP2sRKaeQ2bvIJ
hcGHOvZ+VpaPZPN6eLptx/a4Beo0MHzeaBnDehGSPvvnxTR2OHvbVKyXcWcdxSFX
ksN1yf99DmKSOsjQ1SDfD+0xGlVh1vAKxhXS9Ry0ePnEWVFAO2YTedbgS1ii3aHq
92hEmTX4z1ELTwRIuYzg/1KN5wrkIittL+ZrePNck45neHseX1lrO8AWTIaJSBMm
LWkxP5uQuIEstWQvMUpa6qYijAfReRH8j02/rY1D3LUv2Ub7wAuEYedrvHFKdaEl
zpXbbfvx2FUQJqaTaFoDFpG1TfykdMJnOMhxYHKCirzOu4EmzxYMoPp3Un44jXfO
HrPU/t7JCZ3exOGxiLqx5LI70le1ZX9+N5c3h/0iuJRMBiP7uGl/AByABMJhHX0X
NZKZ3dcWhqOyaNjStOicYzytE6iuOIA95+WiUYesNXftWLBHPUDFCeL22Q8bVrYq
SMRpj7i3H9RjgfpLXqyFbDQAAIoYofJYhuo911yzTkjdz5WjDsOLRjHKz74S5HUn
XoeytsLwKclonozDS8RDOjXeU37+9bVmZTTTy/JR4ftTDOwPwnK00EjLOY+rufTR
4QannWrEm8m0G8FkQ+H4Tdz9PlSL0wxJ2aWfSWuHRvx9qNz10sJlSChdfNXaXLVd
HaL8yTe40yJ9PAmCZP+VFOsa6qRNqgm8T6KNeJ+XKVfikhU+x7vHG9nBhw3Uwrlx
e6ZAN/tVt6ywDPFNXm8MIGyXucQfps6kG07g3kL/Uj3MGxDawVJ884x+MUB03DvZ
BgrWoPo/rFOs3UTVqpZhN0za1RNd5fBIrkI6vyOfQtmE+iGh4gLqK4fUNvG4NdXq
3XYx5neihr9BhEAGFjsvv2anYyGCIHHJe1TZamg0eF86C/GxjGvcHnHl6IWdAjCN
9by4f6zATTfdnoTdWUNYDNz5fRYcbktluLmDqJjImgSbL5JAYLw4lNvtYP7oc/wb
ZFlv9z+ky3GJ6f5cUl32o571s7oZLfLwclMVwB50bWVDrOhNTL0IKvSwJWX/hKkJ
nouvNsYqATE3E5vFXfWviEwUJTO+Fd5tA9ipNe9GVR+/0hHxNIW5U+pECJOAh4eh
Pgz3/4m5FNfbTRmrCY02MIclfn69RP0WwoOJAyhEduNSAVXr4rjYrHv5iIX1j+UO
X2SKAn7GrsZjutn56nakfF9PzKEizXHq7+1Qo7jqcsQMwffC0HkprNkZ+NPRpBzv
9pR8saGz+Bk812F2IKmQdSopiOqMdzkBG/s93TbViIND0d1tXfLoaSjFC3WIL2CO
E9OG33FWkHGUwLUCSKpRsi0Dtxrh/xHx0DuSMXHzIXFjYABnrvl2IwVBkQoM880A
Sb77ycHq/tDjR29qMp2J7p8v6I3ABcsnKEj4n0rk0zXkI7z/6ixNP1Vm3+GzriPU
mucSXlhsmgUSna86/j78iqPteJvYeS3JSwPUT5J6EkTQ5OVXOSMjBy52n17onoMG
dfP97mYRespzu1H8qMBAVBUnOuPZWSyA4pvyyl5zdzRCMuq9JBZ3CS/0v40YzgvV
s6Mi/6QcKJ3DkN/lHiCy/y8UzaC9VtgTy4HEyB1o6/xxle/HtUUe2R0UQZ9B2s/w
7b354YqxeFAK6TWLgPiy4GVijkb5yoQzildB89qLd2S89QldhA8TJj38nbiQ7E1v
J1YKjNu0DuErJJGUfwjFCCJs9dndzCMOoYbLTEQuSyOXb2qWLjF0SLn0T+oMsTAw
3erPLSq69HTXLJrLS9r+CftRFBocYIhj+yDrAc6IT9cx7NeoGNoQywcYnj+eiGDe
uBsAb2XTcKXCvapSiRRicQGLbq3s/FHVfh1s/z+pRnSJiL7/zGlmJpgDbOFDVdQS
vkLxFeGfhuUsLNSNmDm1usee98o07upY05z3WCwiaRU=
`protect END_PROTECTED
