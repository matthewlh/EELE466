`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Iniqmkxu1I7Z7BhfXd1aDxPOjvsS3u0qy/xoS7aEQb1u2jx7rf3UWhw/SvA3w3oj
4tGaRgP4zdcf7RZ8fNjc7yHm0mwWs45wK1KvgmNAV/C4PsYmiTaDwNLoQLBLp3Ro
f1rGhSviSQYS3swEidnIHtZViWrALjaQ73LaXDUl5/4=
`protect END_PROTECTED
