`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
eeVxPkcIZowSxI+E9I27blpWK1lxlryMHXS5By3bgeJynk+t6z6cdhuzh0XJwwm3
Ahnioqtii+I5gZxuX/owt5jZWGKBwY0CM25Y7bOY4THP+xkqiq6oVdunN9R7G/h1
oOqBMBdxfE9Pb67tAhwFf7llla/f8xh7XZ3Gi2DjvxCEV0FM8ywzU1lcg3xk8uh8
gNcrcqdCUMafL6++C82wpFHY+dtRnLrY5jeWZT7YobWoKi+IqiB+miYLJY2RP8be
YZwDCfrvhi1QFfqIihbi8D0iJav3LjsZ2xnoVmnEAkSRTZ2BrMqdfGxTgGl5Y2Jx
AUx4AQisv6JiOCoQhp1nFLSU4J6htOlHsS5EOaRweqI13tdANIXPEJJtdxwA0Ss7
9e4fhT+GosdZQdaCvJZ0xzo57hM5uBvNXzIkRNieloD+iIB5LLEMJAUEdMP3s44N
scCY7m+kUq7Vjo7mSzjkO2h0dVR2En5a9T9ojBdf05irj2/+wg/+Ik5xuV84RXra
OmREpcvFpd6WCiPdjsR19escBAg6E4oToSLJ4rLD7pqO89+HiP6xN8mGC274VDmr
2Q/eND106nQW/gOzSQqY9vXRs2wav7NMtpajtx7nJ5cAeUpKrmhG0mX1TLQAC4vz
2FZwIV9ySqXTIdWIf3ystUBlLjGUdTOgQ/YsunH3YnOlluq0yVZC1PI9lv5cC5aq
PQ1IMXPwfi11HAuKX2HApUXbWf3q88TtE0G77PZOinrJFb59N9dVLJsZ1bxNfU4b
kyg0sKPLUX+87uAS8DlkbbpcSZ4tfp+G+XaJV0h4AA7p+RmlNdUPVvYcuc5o26Q3
FB7Mi/UMaQscc0G0dCJPCdR4joPHjXoaP7FSnvb6h6ZZXqfACBYns1z2LdIpJ4WA
A19J3i6AjKrhfazoHTpoGHV5HbQsZ7igH41xbOMUsc99QiPgLHCM7e19KDiChX40
9NmzemVEUD3bLyQh5OSOSaDZNhCUZYTfWr56ii/C0wUSo62XmOn/eGokOgrWIC5q
hnaehlCzCXAOx41irD0FffVt/mWUwxqChfIL2jcDfYyAjiAJgPpSqQScMfgTsrEz
3Lp4+GOV5Md5kh/ajs0O+BKMux/Glx+OejxQXBdEvKbSqgD+GFYsq7S9dqow8vkc
obDfNAAIPHJ1QMksR87FBuzObRxfIqFVBVLWL12ljEOEZiUvdMBF+kFKkWSv4QEC
icM5jTCgRBEb7SKpFCjnglDt2QX2DU9GbOdndVps0T/MHQJgEQ9pRB0rFAEQEc41
tW0ncGMY/7vA06ANVuFkziPwM7wNg+5k9u2hdBe0WN0fZ/OOGXorXKNbU17Lvfg+
pFuH+vgk2f53n2wL88mrFzZiiKlfDRQzeQRioyxl9EqeHzpZmcTOxl93++1T5XJd
z5mf+SDb1JYyKDHV+x8/RPruQCmI85dQGkoL0sE4MkknVSp9FhyR1QhI3Gwkh1xG
iPA3+A4HEE1CynlAEb5kdtxnuzyVWvT8vFQ0vCtFcTn0MOpW1iXZ5qOKJxXDYs8Q
D86eoMwqHLe/tijqGmn2Tad2HJCflZ8C3MKWws3mETOwNxg2aumf7s6o33ix0qDm
KBi4D+y43CWaDMPfPmKTVNc0eKiJ7GTKag97X/aLdL4iC/rxMCxERcMQ7THh2XWs
horeTAc9zOURpVBgU0wICzkPP8HlsP8y5/clvSd00TpjtBYo+d8ZtWXYdpdPznzG
7WMaxSZwNKb10aKQ8eVB5K9Q+ontRrGerRjcrRCBL7/jp13a93oiy7X3roozKUce
Ew2W4z0zfjrgfZ6vc6mtE49pD95trSOsdhBV8eXYlsn6srzXxKdYgs3t9GV0ywCz
sfXfM+XUEKeaAiwhxScj9Cdg5T9v9fv2jNQuFK9piN7jfDpDqq9zFpv/RhyDZ492
cWLR2slNDdQPhWUhgFvfXmRjsxQefgYA9ZUKa5B7qaKGGQDefctTCWi0YLH97gTP
YWSBJwyeJ39o5ZZ5700l623MFYELBQe145h6v0qLtufVIx77rK4DsfWEwfjpewSM
mRwi827RPYmvvZZVEVOmjmwvm9YsDvbvmlLguHBnPjiETjlIw2StwinKUZpgaTcF
hwiQH/ChfEwAdrTQhFqIdx7qw12iEht52wtworbH1IE81KJso3GaJhO7lkM7Jfh8
aYo7OW2EFWF3lJ66//+acAiV+D7jRDTYT0S+q1HrRYuXjdmrYYWOlxq3nvgsAhfL
qYDN8JVbrtUZfQwq2jAyKvcyaRqppSwbdJiCsraLoEAe50ma54n626lGEyJq5Dw8
79AUyCUb+DyN3lZzQhb1K5w+0icE4CwuCpngaRx5xAocxlaxMqN8kcZW6U69Qngr
GiL3QZm+Z5GL6wmUSMI3g4DPwsRanlSuyMsjm9Mb8UNdEk80p8Zv7BcYXTTc2thp
N/1cPKiWaLkz5Nft9GI4Uvf/Yy0OpxhKYzjmnRDZZt3lGUakqZ5YU8MobFMHORLw
uI8IP3jhR0FS3zhPBNVzEs78qEFKASc7d843Lu6Vre6i5Z3d5QbQfFjolNqe18vr
H6rODwPQhyx7RtY6tH6sEO8Oj4vUBxBabc7sAtKwfpm0Rz9QMiQ6RtJIzQuj6dZH
ERldgD9MVzqf65szZezjMzVMDZeHK/H8mFFI4IWlVcgdAoTTCvTmSWSBLf/Ch3Zm
bd15Q1hh/UzWzZUasEMdYmdO67u/cwIvW2B6w3cz806gY+GIF2lMzgMXlrBXZx3C
A0BgQMbqdyJ2q5ZTYGFLnLJRDJwJBcb3EAkdzcicj4ZXSyctQU7smJ3q93Isq0UN
ah/MSf2LbQmkJiHcgXuqNiK5zuR4LaLK7vo2ScQvrVknEhbJz5JOwNfwBrZnotVn
a5RTEep4k0ZiW4PbY1LC26neT0XKcJq4toVMTlCUqHJlNmITY4aU48taOnHJ5bH9
ocD7tX8LzKGqaIEuxTzp1lGYnhfcrrh05GjBNuba3pQ0iPvgXPuVj4rWOie9/A9r
+2hChHMYn07NfsOYx3yhMuW4iilu/9lhOa8w2/ObG9tcY0UrMyShCnxpWik/Wxr/
N7Dl8ekGvcS0ldwTIgKVwgVTt/TGyUntuOJvpE2C6E1ylDj7z1NgyFd6KYcPE4GZ
iTw+nW1I6rVsC6kHzdOk26flWQzrAfHr+NfO1lqt7f4OC24cgTJY0s3zOOzupsHW
trJ5gk5dtq5/ce1dKeRmQtJwJwCWr6v4AjwWWoiOeVgPI/QUDasx6ArWTKYC+5BK
8cyu0ydCsDKEbRcPBpof9pCg2PgrMj5g9i4YARRBduFxGkqCY/V8XmB/TKQ1sHUx
Ro8/NVotJ0UExkLp8G3SPse833bx7eF8U0luLDMXmNm8x6A8RyQuloud3g6vgyqo
adeM0VLVbwZf5HTHZPoK0KgcKZ1wYWdj2LA8quyPg7cq7cxbelP9IkWjpFwKDGIY
Lwipc/RpEVGaGWV/RTwrKi0U07Xu+dLWTF4O66pleYQhhKsuuSnm0R1Cq9b8uniY
aXhKmpqm61FgmYFxl0LFJProJAl/ckCShogY8PxXSsrAZ5bCKUTndeN/XGvg49Y+
q1+76LbrhcbrXgz2XUoh9wEw3HhkNL7tL77wblP9fSxsPhfXe7VTsVrH3hY1yR8o
mx6K9eyvWgJfyrCNsVdpKe/zRfF8W2xlssZQVD+86xy5EN/vD72+250AArKwsmJ/
AV3qx2ZGlP3ve57akDqXHdUydCRmGRomTiyLpeUQvtQEG48oYzlxHutepNzClIUi
9oFa9P8sNPz4Gh1tWvOKe1Irx5mcrUu2w40cd1eQTTsqh2bec9D7c1IZ3UWI6IIG
ZSCIzc32BLoeV2xjdI7Oqw5xqrB4gSMUhh5PbbzbsQWm/4HXDScmozT5iz9JMfNh
OJU3HUO4XQuDxzMtFNgK40lmRwhGNlANiYAGvFhc6r8bpnecmYntWTx+9Q/WHMtv
ma1ELmBahQ7h9bxajSnfyGgMAHcXKoCLD+c+vRze0j+szL3+7KpnvBQSAOZk8+O8
Fau5vCbGtno4FYJNyZF3Y4eKk0R71pSIysdiHBoIBLZ5w4rvMqHPbNZZa/O0R5EB
WG0ZSNUB1mgEeeJ/gYqBW1nG16A5OWFscAY17/SamSuH/Jqd57eQUnGfsX4yZR8r
EbXcGXMyw258OAP1jtd32jUhhPmR7oQ4zSccgcR9rBo88JpRzdP4vNGUZ92eJ/He
YDvHpLlIxfzA6sRe/22eWIZ/xNKeP8p7GC2P2VLQkESoylILvnk+F8WPHJxn8cAm
fJWjMHckamfPmhwkGaAaHeK8ND2TyzmZSzmHVDxZRLzVSrkJDdv6k5fT9RK5vKhx
+mnvYkdzt9mrbvJvXPGhggsxc5p/qC9HSL9zlBaCH5Ab8ehKveKpvU0RlaDzqVwm
hVKArSrB3095mLy0t/QRdoXpPDB5BWzG//Qxr0J+aYeCD8jmrayd/NUjC/TYByml
rJtghyFZoMH9UF98/Uj4j8RaFztrma+0K39V2E7WXgRsDa2TZTdHF4z/94hGl3/j
q9e+TEtTXl7foKKVucpa3DJ5ZQ9PL302AAa8yJTx9QRIihUQrVF81JzVUu0phHbc
mIiRPaFSj/8JUTZEqU2K+cNco6ZDvL1dW9aGI8fnSYW87NFQpJI7i6D+xfkWMPwT
F3vk6B/We04DUAp4CNjeK0HrQp2EK+VkX4CnTouJwa3GNwc1m1TK+T6lbVzZCDuj
44phLxI4jd2gLCRP2HWj3y238e62uDxzBo/UBRvnGbRKEuCFeEI4upo4pQnjYWrr
AL0ltaf4LsYw9t9W5UcaFipuG3/lTe6z/Gaub+JDVAvEzkUu8vzXukDzC0Wxg+Kj
c2hGTfJ+jEH+WhWTrPZPLVrotNQs0gC5XVrdN36j9O3MuAnxLFL9ci+ssEpI9VIG
I55cy4+JK9YA9oBLWGO2pZxvAGDRSiHC8y23/UFKOurDPMsRUy7dM561ZAv9JNWm
PxjE+NaGEPMBZjnrRfrw/FixDIACr6zAKZk0JhdFQdr+E2VUOxrdBQvB53eCzuoA
V1AdCymn+TgU9QkWXZ5HH/PNqf/sQpDhWB4OuYHghpwW76unSCp1SS5RIdIoKw8q
IBceQgECPxouyNQZxgi6WQCuT9ezNngKG6deB64Db8dyWg5do0fjiu5w1apnBHnk
ivNQHkB7S5k928+VVlhTSkIzk5M4R0siZj3cWSltv9b0bNkxjxTX7rPmGP4Ty05H
O5sPqkxNmS8Mykqz78z/QLycUXjg9zgLL7kHtinhlwBQAflRrt5lpG92B7U6bXiB
7CuYyes1JaIVOpcXXHdB7DqXTkomDF05m0uAxxmByNeIhzlv0SvxTAU7Yfrimx7k
fCPGYCdjaG9+46Dwz3cfnudVzmtrb6OVsdA/pC+EBOx4WMugbBBYT9yKsK1aQs50
eWKop1TEYX33x/jqNttA+fkQ/MHRzvmTnLDm/xLNm1jPxdFBlNxeTcrN/LfhZ4rc
uPByRp9p2B98B6PkobvHxjTMPsEBPKGkqAZFsIJGfKm6j+bM5wFz3aJWeXcyCgGY
BJ5ZeGo9+7035B8glYgesEUTOeDU8itdkxZHaJToxvwi52CS9c9ZWr4E1IaqPy4x
6yFWYgum3UhVO9I75sfq5Gu/QhAeSMnOaIlLTR1T9swfaidJYvSvbUrdhZSNjJ2J
yb1sEMfaZDw3uGxSjt0svPKvE9DNkUyVp8S5VhyGXsQ6WeOpUapvkl1JzZhXE5Eh
HMq3IxoKMCkLmnDvOm8nxOZn3JXDlMjYnSE3oWVIO3HJmmJOQGEVKA67pXj5WhQi
BB7jkDO/pfR3Ntj1B9WOvbfbL3g+yF6Dj3G4Zo3sLz7TfYkPtaPvXPcF1NHJOqHF
hbj2yEcwcyMvKAQDx+GSvoXWkj+MftTjUM/4tvsPdUz8x1Z9zB572h2xO4ZlNCsV
3vhODqkhpiA75H/Pot0bn+/3jFiH771hWXoYxFE5vMU4CuYmtrMeqYxuG5XOKp9C
RQhnxrvD3dFBS2UoEweeR3vYgHfq6qL8TYZELJFnaOtuRAnX6mR3CRRGbpc9fSt1
ZxeLYB+ePZQcG1J2FBPwIbWuCaY+8slaSs1vsqcqhpt1FecnCHrwOyKIvJvKArVI
F/Prk7VboJPUmHQ1UAOm5V8Jp5WRCjxg0Rm4FHNh+gymc7Jv1igfx+7s4Ibd66Eh
JkZLOAV8UlogUKEBIKrsCQC+ahbyUXiNwcHyYsuoaoxvajsQL9WdgJVO8hQV2FuN
UBHZ3mLiSohEo/iOXM17bEJ6FTrvp64QU0ilxuOv0Gs08k1NWTQaipV2HxZ7eJwd
qGupeJcAv+p6+9bw/2lZsrpfGDQAVNniY+ehF3o6WgCMRUqMXXOB88HNdQ2u5cta
Tats3n/gev6zx+GMQaIk1KYKyAEPehEv7WvCdD0RkM5ecvdsdQQ/gnEjA/sdviC6
thBH2gSL8FnW3O7j6miTO0EeYNHYqJbtecqBs8aKOxbVZGPZmg8q+pxriI0qGeS0
nx8qt5MAK0qiiV8cUAPZhL/aaMSQckqe4rTYklbzijMziKVz+GgbBLJe5i+pTtv2
Pxp/xPpn9HuHShPnqJPGBoZTbRVMltCaC5cvVrTfa5H81ZnMJAnCzTghUpccwE2M
HGIlqbyRoIwY77M1dOKa39veUIC8fBDpfcktYpUoaHjVyWC0IuJPj7Im5x869Hs4
yuYCVYN7nr7R9r4G91deS30D6mmmPsofBKvysuML07kG5itQs8Vh/du7RIAh4BaM
3cy7LcMxFEeKTQYcq2cqx9orsaLnH+93jBLn6kxG2D8MSfRAqnS94n+BlDYX1nmr
bqqtCig4VS+XZJV2vvXB4EGKPBY/NkHCeGUP+5EmqNdEieExDVi1xrZlb0hbVZqh
AsI0D3UoZPN2JU7PSawMehCS/+E6Kq+RG9x7XlmGG60+R5mdwHrAx/iF68lq91c3
ex6EEp9NGZ8ChkF+r3/XZJl9Otiig+VS8N46Tlk9ov58xrJnDJFh2D6nAez1TFRC
NAA9pCu3DYWloHRBtzzbEQFRGsKVDpc5xMNlydnIt4tyWK/J0IUVwCujPj0iQrkQ
NsBedkt2rNLT6fK6PLvnXfneqd7E4mAUl7yzcG6Dku7wYBA53a60nfzaTmRcTRKI
yzX/Z0lKtm5QjF8NvNGiEN7cYEtaiKcenP04vM5meaYO3BKIJN8Cn/BDILH4tErE
8daOOhBlTuBEPBdFCF+iOqp/obsWNmvzQSd02BKc9TqysqEMmRAikhawyZhUy/cm
RphcCCyTg/Pza4Yab5q3cSYQ5nwfy2jpT8nbK4ibpkR6ShNLB9c0MiaLnnWEXE8R
puQ5QoYuaHlulk7YKOoDr45sv1cnJzoqmLc0Nom1DvqtaH5V0oz9dQqZRqgz0F4Q
LO76gEfGuibnaSro/Hv+RttgFqiSWYuRmXSOXfycw/7B9REael/cQNzvG94YlcLl
7EtRLgXkOwenic0fZQ8yG59SuMtrH1jj6v4Py5kAsmQh9oJuHDN8ML+M+eIMx3r4
RwLgTcM5k5q+7ZYSnfp7igQBdkKtx7DCjpK/yLiiQwqFDqJPKlHrw7bzchi455hy
rI7cFJQ+1ZHkYNp3ZjyMFZHQk/1PV+GOcPPboqNAoTyW//H4NQVAZygFqxe+IbH1
crwDC4msTV1GGAhfLLuFrtXmI/nMNVwIccb1UQf0KyGgAxcqHsJRbGByixclvQLW
DeeZTGB/HZF/oOBH2E2hzSvNaoQS0PIFOoNdwzwz+9/eDkI9pBTs1ZgT2LFEDEMA
DGRU3BYqpVtmhnggwVJAsJf6yelgoCVQ86dodadkFlJsTbK4HoZfwB2aLS7FrXou
JCtidC8pjZWnY12yF4daUODe4e8nNGPQSqlqkDb/sZobfpvXD443DqVYACS00AjB
GjHQLzuEHSq5Z/V7J1j932jrr9/SpoKR3AW8Chaj8ufDX/WlDbjY/FQZxqORpMPY
t685a3AD4p8n73AkirCI4fxJnlbGG6id6gmjNJV3qbaPKOx0mDCD6i7v3tYNlKsj
NWdLdDEgPc7TmKKp7oB5QTNPyKwRSc0kq3JvoKMbTIonZRwCY1SpmlWI0LTEAuPT
+gcXr2tk4+nfCjdoV5Ti19a2ChZZ2k8mykJsHJOSajAAlAnMMFEcUZegR+Y9RGsR
gddIzg7/i7L6otQvOSlFA8sU+cVdal5wEwqbfmnc4t1eNaUqQZMalmcGL0/JBRBm
RSFpw2zKmWJ/n9QIpjcLOpCyp+3RioFz6pWccAApCu/9dGNH0OCTDXgIt4h4pR0g
saFwG4tZenKVsN5eQ5MebhkiYXswBidvcUpLD5M9CITNUFFVLPbxagGLh0NmDzqf
lApcBUFhNPOIlhEDvzD/B9sIJ3COBOBRPa+l0j9gyt/5e3zpgssZWBX73po7dn55
TOYlR0uaS+ValPrXsDOkRTGhsZP4kYiDNwc7YZbedbcYfyxbVHWg8coumI/ZWmDR
DYylnDCEqDD2e2b4Jrr72uV9wdo1qqeD7G/L6GxOH95RbBKsgl9GBE2yOl0Y9FGk
mUgyj2ceqCDZoYB9499igjMd5Eer0dmpd3iByPYNT9sgwLDiVaxOqrLAVj+Dg24U
NtBxTU3HYh24yKl9RJGXKqC8yN9oVwRJ03Gd2OAnyg28lHBfw6y4SZqqNbewuUVV
y5ZgFaGoWe9LXLYQSZQClWyBPKjWS+fYyXdIgM/KwYcaZlgH5r/bpp5MWem7SPY5
blTxSTx2WHyQd2RQHsioxWM/pFlGooO+aqGDxXTg6OdKz7wkPZUSrm0q0+Aq5e1h
bfYbIWDKOhVaQX67jOJEDto+6COrphMmR2DIWIC8ebdktEjxSFa7yuyA96u75QHr
9WXb0pYInTzJwnB9dMFlZNaOf6OwjjsBGRLCwFwx73Sdh6yNaUbtzgcdXWPIu++h
O4NAtOeC+WsbRYgy9syvh04E3sCyz18US4vYxFxEAJ2h+dHUj2KSUBze0zqYxf/R
QTjDf6l9J392g9PC2K0SqbCPMZvQMwl7cCTeP6hJbEakiZzKefFQ0LGpMS/nHfoN
Rynz13J/twtewcknEGfujnahARdlu4DNhBD0oRa4MY4xaNlQcvely9cIQp7Z1aHz
ZMCcBUqHfvhFfWsaBbNycDfSa3U4uxpupw/xrjLmfGasD6SVcpTGNT2wGIgfonqE
VV8tt1ZdweeDiX8Q6AZVepv9pJUi0zSy0YwcBBMiJxL06k59Qw/EvxizlpPLAADd
R6SupeiUCJAk24rwY9I0qX5/MXBo9Wr4QSFzmJ8lRe833/ZbkTBAHlEheJ/UVdHa
svphjmEG5tG9Nii7vzNyeCEMsVz7EmXvTDi682CXLfjBxB+Y3fo5wXoeXS3tMfoB
GK71qwN2X6K1LjlmwVU6R8bnGHwDKjjMNHKnLuuyBxqD6tSCic9DXxq0efu6fAB3
ukn+x9O24ob5D+OTMJm3xnxsXnnlJBJpL2Y4r/8A/XjqQl5ApBaXr+2W/Bj0djNw
cgrxKSCSaE8Ad65eMl11fXaaLmkZm1WTuzxE6LZ6tbQddmBh71ZGD4MaBU8mI75Q
dkiZhFZIWETUavkbZ6Z+TSEUomIT+6wongZ7Rc6ul70WC1lSzMKlTYHaNIBUfqgI
QFVL3G7IJSGIGaiJh/YSbt0T2rsScKc1eS+6JfT9DIykOp3xheS2425EZNaUVCf+
Id7mLH1HGoNtAkavirHSDy8LFO3jQM7d2U97FEI8GXw8zKUe5Ngm345ZJCSs1S3Y
GYMMq4V/rl9FKbD+obVvwMmA2D8dszQmJgBDayFjWBOijMMTtZEAdL/o68GCfC1R
L/G1N5iMk6PD2uxR44+WkRHypJSW04lQPkGYLdHOnqzoqKpvBf/8pTc/q2njbmcF
pzEbN+JFtWoE5pzikxKoZ6PFQX2ZAjxzlP9Vy5WAudOVIlqpThbLwR3Eyz+lj3h0
XivquJJqSsS4wNsao1n4qRtWkqsZJUoa6cqMla/vwfEqETe8YCecMxqqSk3o62rO
9D49Gec1nGA72+vjhGq/l789PslmsVDN3HNBsn3phA7+sCglCrnqG92TdoNZOTFI
B3RbOrrGA6gnbYf6D1e8qPTz1xq2FbqbdmwuW9YmVMe4Yg11YOLjl3ofRUZ/ADtB
GRmXrRDVcC7Ka1dNKQ9rBO8ZEUxQVxHeRQ1ODNjqmYDj7WCdy2ea28sL3n/pOYKZ
/i/MrwBguxc1wvswHQ3VHXMdVWWV+9QVO4VUOtntT3mMcetVRJsuQJ73trK2fs8N
GqOhuV8fJMGNTYrP6WulXu3CYDfBH6K/QCAdLKBwSnAk+Vnp/1C/R2QqHWflcjbC
UoI07r2ghnoPWYbQvkJC9FiIV+FpNxoYVE/pYSnzSU1f91wP8fOiz5O8LLW4mphQ
Wml5bKGkVgyEZx1LGyOOCNEWtzhS45GzxVT46BzwJxQG5TnMYZPuQsQ7wcRyY1mQ
+Xh3QurWW9GwF7zr+c57/BG5oG+5CPsShASaA2Gld9N+uUQfeOyoTwyhtiIRhsXH
jeVADvCF1HvuiYZUZ2WZ+aBRMER5wN/2BAHoA5H63VQudUasa1uHBzfEvdnMUo55
Uee/F+0Jv/GcUMkpEJcTVzQD/88wFy3IdXoA0MtQUy2ExqU0Wvbx8n8i2KNnGPOy
cudURzznM7qIKQGWcXotveWEvrJPUef4VEaoMahuEbszKCes3VKcdKjpOcHe/0Eg
lRAy6UkWWEit1GLMP4FJwg+XHI8BvR97IZQkFEOgxj7gza4vVRV6/tpRr43ByLTE
AvfRprwta163sdN8OHxk5Vu6nmfUTlrTQaG6iaypYQfQAv4t45zoX0ojNEF0nfUW
pixqgARAEMNTtG9bbCsG/WENkcNaV2h8Rx4qcN/S8Q3/XNOjTScVybUo41orCV/i
Qc7zYq/lE2SmK+ujV5160d5F93xEejHDjiw5tWQ8nNlsMyjqoBmiHd8uTw505+8b
OwL4j+2zHWhw9hM1R/o+sFAuB4WgS2XLyv2cNFOV+8jE58F/Z9FsHaQ16WAc/b3G
MZ3UHuo1N4RvhMliKVRMlqlwQhzTIn+PnaO+HOlQ8ZsFwHT0emBrkCZbTiYlultX
PI0xUxhvg2XY32SEAVW5u6ninhLRE/aiRnn3kxpiwXI/Y2ZbuJdJgh9OVQJdredF
j195emxiTh0ccwH18xpCjzxl+PDpE6DouqTPGbphITrRRCYFyPvrbAq7K0sOLw1x
8sYPXAIPu6DqWgaVHJVTqVDh34HfH2DPn/rgTG5XwYev2tYdkQnTOZZR68KWcgZi
x2Ry3XFeHkWhS8p+QGdVJkafKUhvvSF5n2ZAdn0KI6oMPFMDXXFdHM0OUgenGaqs
mIv9zyqA0XQ9pprk+a2ffz0iQF7581FaTBZFf0iXDbzidcheqeF6SJxCGCyvOgiA
jXrvXrN4BW3q/hFWTz53Wjz51h/hBatH0APjLCoTCFF9X4MIMPsyQ4Oly0PK3wX9
WQLTybxN3Bk3+BtfwUV/B02hJjeHF1fHcYJXAV+HchfLfFaFJoq0kDSKYTHpEear
V7gTUBPEWBXQhsMm21st37jJ/BAx6fanYcgRyb9Bt457GuPkg210GEig3CLrc3/i
XuROpIXq90PVlK/6AQSyezhdb5wgH64iSkvGlJ4tWM1ojTF3gHLpCc3r5MtIAJqH
Mrqjkr/RmGr+iHJvUiZDamp5Dc3OuZ9gVl96flQ8l95Enue+U0tfoo5CJhT4Su8b
z14yMmZSai+Z25C8Uo4oLwLShKFvqzjNZQHkdorBxE/U2xw/p532EAjx0+wl6bw0
DOGx/r54+ISoETZYtZDFYF9kxMron9WnliBe7J26h8DU8EobRQ+eKAtpfJF0mZ6N
YU+PBu6MkeSXvdBAj9qfB8Ax1H0M9IjkUvNaVkOgzLHOrpOvya8SURHsiHJntWYr
6GjK6ZiXTLXPHqLhlFShEqoo+6uNYJlemF2cGpGxADA7Oq+dWKXYrJD5V9m+G36p
L7i/xey0AX6/DDhWvTFLjd9BzmwSOpUV2ueSRU8E4zB7NrHOOo5NfA59OyfNLzrl
5xu3ai/zCjb0gcmT5k7AHDhNUsIQkr3ney4HVPLvjhDs88d0mpu5t1zjjpOfYJyC
2/uThnRex+3JDHH7vWGTSj/rcF02rPcMhqy0Vgk5NfIr55MSZRCxVBOPMJ4avcVs
xp5zye9OcaYII3H0TzW2GBBIEQupiilzYw9oq5nrfYt6s5px65iqfy2WHWpoQEEz
yZNCWwIgkq+ntlUKr8cUBO2Ffq/dq6Q42uvlKGzXc7xp4W5uNO/DgpqxRM2zRKVh
GBr4X+42YiBgl0+DQ213qVr9EBWr7jA+4d/ThUSdAj8n9R2/LlNknG3GHejRiVPZ
TYx3bU4dPaOfuCsDkTiAXL/EbmEnMkF2U729145KONT4xYeQ50TYv7wWnemfWg0S
8cwsYl7DkiRtQFe22E+1Oc4H1IwG3Bp/Vb5GePf4y0wh49CMkxfQ2Wz929I3sSVF
mi4YimxwHqChgaYPBfZXbqV0GjI6UEwzszTK30xX3bBCKRcdHMaD1MY9Hu0nJy0d
iHRidGLy5cp0EN/87/9t5GmGn0hnnMglqP61JoyLWblT8WHA9+KbCKAQrjbWEivH
NU8X7WWSTvAMXrC6q8roQzRbVCgnWkTEyNhqEMAJ2Jt4P7nJlCcI9HAAZ0lnrRxE
tcMPMD9PpxlFcg71Lj1VoH7KU1x+1jtywgN6mAatlga2sM0mk8+zs0lvywgJLkXQ
uKvKsqy+ZLWmAN7qnf3lmnQvS3ql2vJBuMM+yr0pJyb6ncCgoUGLmRds02bqtd1S
q4BvT8C4sn4x6ozb1xTylA53zNZxEBAIfqgLNB+oDpKUQjqdAaatOm1Gv+GzXkfN
5cCukxXCCKx1pf0v9RiHqeLQviFfc59ndVunU7NzCjIDCoKsqxGWWSYSbH4NChs6
7hTkxD60XM2C8gv6icfrMZ4lbodVh2lQS0l81tLUfwHBCbo67pijX5/wJA0M2MbD
dMXuuceAR3c5jt9bYgdmG/soiVweonyNXR9DXP1aRAm3cIkRx7oWbHPeYuRJv9Jk
9Uhnpsq5ydtFq7NXB8FWlNW9Gci+FdqdGl8N3dY13+PJq1Gco6egV9ng7zw0X1Nm
VtoeGXwmveLtZkw3ZLrNtBjaapLnoj0HWXyXy//+glQ1X2brF97SpibOMc169glw
pKs4RM3aGqhTfZcO1mwmTV8fcYR+8eU/cxS7gPxAzS+A65xjNBeEezNwEt0dJbdb
bh1UwMT1mkoN7lOmI8TIl8gyJtzsip9WDQ0scLaP1lLCL4MzUFiyex3urNP/2/Yf
Cvm8NLlGsPohSFaQfa5GEmw/8aW5h3S7Q1p11hUg+XEC75W1DMJ0sUTBy2iiTib5
i6HzRcIM3co41C2aBXF4neUVik+Sx1V0QaXFz1AMm4zfVjzEvRWccKXB5aLVqc1v
+QcPFDkGXxTqEOgu5Bwj+qsS0ehF9AvU9Yap8KcWJnSriSReyRoflgZASAgCltah
V5mIAfLJ/9QaHq0XwqQ2xxiOR6lmDsUpYJ9lA9NytSXsEJXDL9UHjrpkkzxtpP+q
tts8W5Wu4GRIyPJZ7i5qjxb6HbQPzGPoDYeUGpiV/NjXc/YzQfmV8+qhjrhyIQQd
MxrdWueHJ+QBSNE0t7xVB9mjM5CKS7y5pLbDljA6qoGmPWw/srykVarw6m5PfnlQ
3DslVllKN5EZtc/LkZgwehG5F+DW28QgboA6EVMvQttYtP6iwfLTEigy9HlNI2Tz
RWvvi5gvziGFxJL0WFiZCGaiW7skeTmyNUFJvBCBCtHj3jPJxI7oQkNqA8xPhGm4
HuT/A0ePonSh1OlnTZpDB2e70PXPuOWc3ddfxsI1XIT1c1dLxe+Kf5EnMYO8fhW9
ZKF7QysPZMDlmkdoPyNNdXZNZJ8kkh9wzraDPSKbbk+D4FpK+ZGvFgrP5pmG2B9j
M8ZndZX6SHmqgQ7T67wbWXakI/PhuymLyH9IrXSqOFqFbGS7+9usnaaQD4Gr9TPz
VrMfKFKwuBtp9qi3FBImrmllHxxJpvJq2zyqw5eXSBN5Y3RZ//3b/TMh8MW1Z3r4
PO7czVp/N6leDEUAUN7xYcOvODgHxPB9/vvtWcaBByaFvJP7oPAoVQH9xLGot/fq
XQ07nM5r3atuYpEv2YMMDYGoR0RDxfKICXgjllIJE6dwxp8pCqZtDBPQ4Rz0xSu+
mTdz6twnFAqOfFM/2T9mI7Njj0Ao9S0PSyGiPHuyZlPXSCNwRjKVNznfCP4Y26t6
YdKddGbArCmezma+RJLwL8pZjuWoL5iUktC+8id73W2PsrsoCDZrQJGDNdrLbMPY
AtsXN/cjXhi1FhBZE45DU5P5A9uOLB2vftfdiSNRZ5wjOIjNhOCVdPjBfego/jUv
gixMGBSUvkkIfQmeFI5whH5jfT6f4g28jRWjvMPA74XecApran5Rrvm0xr7mb70b
RIIAzlL6ALgpdubf9N1RirerWHnOXXJppVyZgJSq2wFE8kj/xFWTWdB8VGlTA/Mm
jFOFt0i2pcmzbiC+iLVIj4r/nE4anGKEW113gpeZ58GK436t8WJ5Y65e8Jptl5Jw
XyzcR605BTqZtwDdVEvuChyaaeUKooi7Kck822AEwYNLEZuT0KJ7zJMqUZouyKwN
Aw1DJ8EPuMNl/ZgyJdXlJSp4fjWA6WdOzOWi4fC85IEOJgvGVbhorL5vIZnuyJCf
H6MuvDyqVGNB2EkvN+UPoiPaEWNgKaHoKpXZzusmwuhZyGNSBA5KNJnqPpZum58J
Bi3EgVM8X/91VyL9wGsHBadA2PaUsYKSmMrbdygHWSlYqNu1J9f6B1TnijS8EhBO
p1XKs0M2kDbC1FlGq4oWsSmmhZ0R3kWrvqGlFT5Hzg/mF2sRF+aLPweTrVHjTfB7
uMyGGjFY2nlsdke62vgyw2t7QwymeM2YzI2SngPyBqkeXS+UVNxNwwCq9Bk9KpEu
bsk6eOCs8WvM9TgxSUy0Tgr7xIi6PS72cMpyC4TKvQJHH2UDlAHc5PrBpSVltvE6
u+BhKhBZFi+UL1BUvypfUA+et2HDJTdaCG1l47gmF4roP5AupfUEGdzB52APaHQH
ytgKA0+FqsVDNX0pt5bKn/2XuyA5RoLDw/+w2RpiVtL6A++JjkEICKktZ7PDZ4Kf
Gs1W21jgyAc18BdzF6f0wvrySmI6NdhVyLJW0uMbRKNSBmhcGibHo/Yye2yO/c1g
7NZfHYfKRQqb6noId9/oO7EXnrm6rgOEQRFqsVAKIaK5PXGfKW9rYxOb7jn062yX
tNpl0ZDyv9ofLNBKnpft3bHTjn7eL+n/b/2H3qEq86S3p3rV+NSHKCkqZlrLXRxb
E5YjlkTH8iJ0F9VPecPKXU0jNnMh7vA6qL7lGSUiut17iG1c2iMWXUnRo9jKkEu9
3nVXJlqKgVPuOG5OVSkC28KW4hGr1KzT/pI6Asgabm1bNtWGifP93nZmmNvKEV/A
/v/TZtjW3qS6AsTk/HErxnKEoG1U52Vku/IpaFdEXaOvr5I8Ead8jkitjmcekwY6
FnkuOr4jAwf4tFbBiBrQ5ArTrKJ4oZw+snqOtla+DYyBJlSCnK9RGb1XCB6kdRO4
upJvrdjrBQhVZ+vNGUCUFut+1bC34WjVe3mK1PTFGLTnilp+rrKvEJO3CT3Q7nEE
F2FE8tkMDR0qi05wWG9gk1v9SUVtgkeepBFa73eHmr+OhwKRH2jdf0OCs97Uz7Mq
n8rHgERNCFuZRwzh0bVv0cyPFTwooQbp44vRVEdt1b8GMGAebmvKzWe7GwLedjZL
zrAUCp/QZ/F8fMaI/4V4S7/Ucheq6FVtf2W3oQrG6QO0Jy7p6DiM5HCpgyZMCrQ6
k+ASEGOI+qDH+xNdg+e3Td80225PoKkIezfpx9zja8ygY3zQ78N1SnH4VFWMZCf9
xEdTg+ykAgfMMPV1TUry6sHiZvvnIwhDp6dcYQXgugpqJTOIl56gnUqq+d7A6xZf
riv7HxeSno0XrMrvlAfPytzu1EPZNp1ZFIvymHOPJQkD5vZUSwE3YVMIIXFRpoyg
ukhA4k6/FYB2wEpx92dMUiyBQBkTUNTI82zSboamIXvteIFz2M2kt1wW7xPcwjSw
294CTSMsrxOHpNP4DKfXSCYVYzY2Vbj7Lp5rN3ikXgxQZ1ejueXCLiEIIqsY++1L
ACRQP2LkpQ4uWcv2V7mzrFIP6mLScWQJeGCWD1QuSqRuVDxGJkja2cdM6jC7e4HR
HhtFZdUAqziYrjMAa6gPIHkwfBTrbEFs7q+Dt8nSIFHYUJW3DVNr1K1xZZuk5p0u
0VgIuBmC9QDJsJW8s/kMuziPxwmg6jvIZL4KZatbLFmnAP21PLKKWQNQFBM/VtTk
mAAr5ba8lTL+QiHSCVmZGw2vmlwOvsJPwRDrufVJYrEVEm1/qlZk7FscQbY+H7J2
8up3LDDDOKFR8QAxqp0L8VzSKhu8Hk8GxrXc17inhXH1MiqB+xYSkzOy1/XqJjOu
w7w0Xcxe2v9fliG/LeDwf2F+R5a0LXGA62z4vE9FeM92FhCHmewg+0m5hQsxaSX0
YRtoY05DDNHBGruSA7Ujn7IxQ+wb7Ar/APhaixR7ZkW1DwpWiP6nZ2cED5MyZ0kK
zVXf4qRNxuuzIw4N/NMCG2Ap864NfvY7EHvQIqv10WQZZhHTyohwe8eNHb6SSwll
loyKnMi5lIER9Rc0IyB1+YaY314H1w5xa4QGkIa4cAoJUw7xgV/IsPfquQLU9Rc+
MV23swtZLDDVunzHzGxSoTa5zdGJN/G4/DktLlkWNz5LHxSiFjBE3Iql/ELOSbEs
j9SxYw/f7F+FJKkQK+nksog8fYDNCKe0Na6HIz5cwgaO5zRmNv1s7pTcn45Y22P1
r2uTjx9erXAxpowCsQh0uRypvLvP41lVd7MTtUroaSlgB7z3+4le8wZu7bd79r70
E/4M9qOEB35jQIxP0Cg07xNcbMhbzrwJ3p5ucUPxtykoRRJt9U4AiEHniAZ5VUtQ
cQrInQYK0GQSCZt8b4NieUooEJF7htq6QzrL7bFzzdQDmBgd45ZdmWe8+hdfOVR+
mIPmKHHoX69FgLT2N+mSjN9h8sGngHXcOp9VdZ8dWcGTiga6Fy9rnLBa+Y9tnV3S
2PouOIQobg+VkMQjEQvz+kDGtIOud7UM2QPLZsBv3Kix/IpF6jGanoZvb9eIGTpq
GHKM+zSUqMWY0u9FXmZ9SHykIQbE2t8IqpGjanQ34xqpiZb+tyDeI8US6DgCcBZj
aNdJjuGPneKgHo2vPsupIOpxyTTdqfK1sq912HfrMtwU2zGAX1E2BK1JAG4gwYT9
Tuh9w55qB4ZVYy1EYFeNemPePxpDXvdJQOsVR06+Jez/XzbpXaUnKh0/DV3HRjre
QIrfVpaTNPIaSXudwmNMX1u0A5K8QDHjJzF4Yfbt2duELOXHF/9PlKA+Xfkhv/5/
K8jTxSSqNdl9okaWNblv/GYG3lFtFDEs6LtlYluODnEK1j3d2VhK+jp5W9Af0sWh
tULscbnBNFBf9YcDi/TOznehFY96OcTCiOtY30l3PXKLaG066HA4cpUBBB1tJ6E6
r8KIGl8yR6RtHCnxjqnDN50oUD2FgbhLfGLurTQoK7np1pst1NXAX3pv9bX/Wrx1
uojN+wFJDhiCO8w7GcNnTWofhHYsyyEbi1uheTUFHVW8Y5Ip3JZgVShPqXx/+oVC
cYEARtnaUBcbceV01zc45utthXaJkda1SOakrLD7/Y2koZdKUcZRVFkZMVR9CmmT
LOHShUFxWTqw+MWb/5Lp3uzRtuEqXdWq/pML7sCNEtdB+8C/yr+ofLw/wg7SA9e+
udOsRMPQkf4wBSpc20BWPcwYwPcgXoyt9Qa3pj79qLPjDCpjjwYjhoredpk5xUT0
N8hASiSS1RVycHih5ZEAolmqk6fzRkEtaG2WJl1rvA51JEkMcOudRHf4qWVSEZbN
ophEupBNjm9Lqq1M/K+X+jMhOVwT3X0t4ib6haDHV2uSnEICxYhJfFmqmmd6jHSE
fyx0iYbub/Q4yEw2DYQZiIeaN7hwAdJQ8R59cjbOjXg3hIg20KRWfRhuV6VtnX52
tf4mDdTdHx38+2YcRfOiotB5bA8knoHa+LjzAlD7WDlEvORrpaVioONHMp4H4Nf4
T4THpW73wgN6X8c/UAJ8Z7Cwd8PBYJGRbpwriagv4/hptLit8PteCyDPPuMyLfQ5
W/YgeYsiwzBnPiLBEPrSNK72gIND77nOL6SaqSyeUy9cT5f9WeOZpw/8/9p+Q3Jq
Zd1C8zgBim8IWLkkeJ1qyuE5zm40My2vWQW9XvAuF5QSG3DF//mLRktSIfFKUv80
fFFXq22SLhp+PhiKfAoMXHKW7BbeSg9vitRAC2yEinu6BZTGDt6v4w0/h6clFBG9
R+FdBnttb2yTqc0/n8fTO4x/C6DJ7KcGA3UgJBQcp0E3GNZeAWbipFvJHyPHFSmD
qc5PiwX0Qsugmsz4LbYMoaAsN28VBYmJyvlg7gJQ+KEp+HYKwT5+YFzVrVnIuu4H
NtnQkW3MdqFgudMrZxCzLX9GdFJcJQDCtOrZYyS/e66GLRjJvEbImX6d5X1hdU+c
EgNKiN91nurZ5cK88o9PMGa0RoYZERIfcABnCiExH+zFi6iKkhFUXE4bCDtleeCb
IrQu3Alpz9hH+SySmakDDG2dPGu2ydF+oI+ZngVeWuaJCul/eJoPn5S3t/etHE+R
pu+xDU6Oeh7SiNLYxunlosMwtAR5QfTYRglspkgzp7bTxYRF7DwtYL+iy22IqUBc
XejZPQNlupxvVa2lgm7YkATta740tKwteQs678b0SOdehGkE6uIwvWp4eGinIbTS
doV2ezdcob8k1J0zEd+7fatuIIT2oxfB0s5JSW6xU3dZtaGWtrBODyAYjrdK5G4/
hLSXFtSLdtIezUPDGrtN8VLYYv22RY401SYPBt6JzgCSJIB2QVtJGvNwiW5v5V9/
D+pu5Ayoi7PVvDs78eciMBT47C0PYgOCIjvE5CGZTrtfnpu4fTcQO27esYfDHuTN
zi7SOg64947eegxhWDHR8YzhpYopo0PtJKrk+vDCLUZnrOgvlI1nKdq506jkX2Tt
iefdw7H8IWM/86IIs2KE9607K6a9m7fp5aFBdER/oxvowEw6UbltVDXsdpzlAj4V
Mco8yiQg/hMiESDVJEUa9RqAS4bQyc9uADnQj9NGFde9Y3xN0eTikfP5BPStAgq0
PQboxqzXcdcVuzr4m0G5/f561DCfer1hWNeBedJ3mJ3wuC0oS7AnH/QIR3U+E6sH
AG1QKWlxXKqzHO971Xq4ceT+ndC9ggbkIWZM2IWgR1GosycsQ2YIUAq+/VWeStR0
mLbCo6p5+8OVfAUEOEUvhu3Zv2yJeQuCJYgpT4nrN7/Oo+CfkmFJZvptsJsZk7rE
6DrJMvFgha7QdNU9/8RSkdEGnQLhzpPPloN35eO4JEHmxAooCgCYGqzT0t3iqbii
3pmnMGn8kVFlHxbO48JwdYQ9jDxencfCxlcTacV66U5FXArw/HA2MBMGxhke32dJ
cXho7Aeh8HyS+ewxpqE0fQea/cc0vr2NX/wla7poO3qhwAIl7n4bB+wnxcauSGNE
Ho6ESHZ6SR9mO1aZCrxTfWw38cUjNIePKHAC52wzv5Sw6w4ql/4oz/UL/MbvQWsK
ZW8iUj2YkMxi7FFKDeVJOu0nSe/FVAJxbNUYpHJMCu4c0ikv8A9pJbe43IXJzeNG
FKpU6GEhkoOebvhE9WpfoN5oxsn23zii96+5n7PmrlrBndUX4b8uFWbODLOSVNZx
5GFHDHk7o8rQ61RtB2DxyjJTdRjzhLYm2ubhw3IKs+Ly80hgm4HtlZzfCBBFOqJ6
3H0d+9Y5JH9+oEWdipKfpeaEtkjRmObwLx9Rxx9BamfsfvbUYgtQB9HglTpnQK8F
nQ1skLO2EjOMbu+ZQMVuAdQwbrOHe2haw96qG8nYLA0X0JjkQcjqyPNkyO6R2g8+
oEeHOTcIBOJRwvAEaflBESJIoqg2azQCxeZOnagZeo6tbwq+D+5++eWBwlQTyA6M
UBzQ9kNEfql9X512F4FsUnQB73fDjsoL4fl0+uYSwJfjw/86l/KD1ofAhWNQjxho
ekMiLFUx0yHJsah0CRNz9IK7vYeSH8f/mc08g/b8cefeXqBjX0ebw+txY+EMbYfj
UURmWoeiyCJ6E0Ej3tNmwij/gNmazLbny8DkldwM7PBa+vEHC7yhO3Wn7pWHMS1g
gUjIuKSN9bl/v+JKBXcCzeWk2QkSZkwmYy7Tz7f3baKnIA8rBjQoxzEmvVyhJZwq
ZjbhRtZUu82T9Udsb1qFqXuyCa6jsDc8XSXTaDIQjo1OWk4Kbbb9MR/QgBOwdZ0u
W/QM/py3Q4ynZaZaqS/GLD/32pC3UWjqrCXAm7YHvw0dsYzDcyrxx91IJ7vNh0H7
lfFOqfyJa+sFLUWBqElOUwn1tbcOX4Ohug9QYcpBz1BwZXvJ3V8UJr+0ektO2Wqx
1MBxumyMzlt0KTtA2jnH+nM8Ao9TAY51xOPMhNn6zxfQFIWHs7SoJJLv++vjr01w
ZswNXvI/BN1ahq3b1CXEd8SW4BkRs57YFRWF958Jg2vkXc69ZxzJSMLzCtYgBO8w
wsa3q2QoAiOolnHu89ns2T2P7qSFMlwvZT2d1mD3aopXdgKXDitPVNGr/uor1av0
wqH13SZtIjm5AnenkauC5EbvNFlfWaq9+xUS9M67maL4MlPwqhUjC9KqexUTIssq
mSNLJcdyKBniHERw5SksRy77FtHmJAubtuc+tp5gVAp/h6cUhahLJO17sMYdejpn
wPKrqB+yvsvE4b1Z/5ttvksuUZKIp0/Hro4bP89msr/yI7sEKQJXSpcWn2ajTPs0
GfXo85VXmJ869mIkcWySRvaRcxUwTaAhO8n7KOW3DBFBz7ydwfvQf1dEKly8xEtS
TMzNGnYS9ftLoarZFgz1rYE2bXrrp94wgVW0IvKcPGtUBe8Rf5ldBOHAyYzoF3kL
BeVQ9G5xjXFetMzEQMJ9cA75k5OCX3RGFMhw4wEuxF5aaYKtzB3qyvTejhK66UxN
WD6SR+UsU8Efh0i41SH0Ab4Zd5TSzNxUBeWgittxS0wF8YTxBLrZV1OaXKz02fpH
NqhPDAo/wOTI5e5Te59p+mWYfNciB4hsMhlnJtL3J9wJ4PAxRrTpGo/aKY2Hz0Jx
iyrPwbDnuTyThpo6WM/h+maUhUUsob/XipAVJi2jNjf+H9ERd90ag0lDNc9EtZFL
vDHtByWAoNfEs7IowXBXdB95neoINRhRMOHBSNrsmarSEkDOHLKt+ScevANKGW2j
INpH4qqvGOb78RE7HMXggMMKDgf6I8/Foy8gRD7A1P6383/d5Z0T83fLgcp9urMT
X70QCdUdw3Tsh0DhxVjkEYLc7Vb4jbf/1IO9nBOgFFvh+xJIJ6uKS6Tkfrvx2NPn
z6MuSvRnNBNg9Gc9xyrC1AhQkXJTrGYaIcjXYKz7tGCDTgsNkhQc5wZYY1Rqg4yP
ovqj0ZocaAJhMcHU4McfXyeAXm/kVXwSN9PPKZU1Su7I2WfVcjgxacBL8iiGiKE/
oBve6ulkdqOvIEQbciIjSdO3mJFpTH3QCT4ElwFKFlw1hb7eIn4yZAsYngDRNfhi
KLki/2vzVfs6S8pwMYZVphA0f9P64DvRzqtnA3z7ZP4f7d/rzQb8cykElJgcEih6
jQuq4mXa091ZMBbc9gUdQJpB4dZrej1ldT7cDmAxXKlbO+RS1QORLfvHE2lF0Vlr
1YbhGZhZnSjPipxFU2MombAj1Zz9P9R9OmiINlgvEgc6+gKix+P+WJSequexibQG
/fYZ+9pqUeCzsizKgK2UaOxtuW2Qoa0couio0oNYV5bTco+8Qa1fFh6RAohRDC22
MsQNVwjO+yvDqbzqO8hHSQ5NdAk3OrmBw4yPOSiN9L7CjsuNHnQv5Pj2Xawm+yxN
dioYOU8uzmAEkvVeExG9NwgXomOCehyjiSeIRQYDpt2nbr1P76Y2ZrMh2XmIikxg
aAjLS3JTGWwGEYNMhTWAOUevxF/hYfDsE7t+r0HbUKKQLNBrHzQ5BqLj3O7zxwqf
Xf63xjZku5AN5MToHj2t11RDml6CZSYG6aJbwzlNX+fElZwOrF+Xdl8Xlr7KRaiJ
PmVg4PG35Tg/8t8WVzayPr1QGSHp3rtAmZZPnSj9rkuj41ucncZuReEi0uJHK2D0
sHWG3EFGijs3qFUCSCXZWB0o2Yg9CYSzVBR3eAghZuA8pwDmv08EWiF11Tkft0rD
X0KN8E7G15TUw7WYJbu/WjhnVsCKEu3fj/p/IqWxxlIcbFwTZm8NKJh0Hq9YYizO
W0ATsIobygy3Sst4xO+GWPffw3ibOV1ldkPbeQtBgWHN+AC1n2x9BQYKIuzQCg1g
qTRwh5ePvaQVrDbpwT1lFYFTym6MRl/66zoqzVgRTAhN+FVq8qMTkC1X6imRFLWB
XdbWqtxI4Gfu4NTHACehhWkarl68q9ICmCxDpdrERt5wUtnVOcX2n14A7dJshbmK
Lx8gtPOn8CdTeeNL9xu66E2iOa6qnmusSiMTSv972Th36nfirgC3IOcx8M4e4K0S
oGkDGj35bUk8NGcQLjllfTpPq3lnIFcr9tPWCii8oZR0/5C+0Vdzdhl1nnaI5so3
RMwngNajOvXyhSxDk6BbYW23Dy9wJbPVuE5mNVdEi5si1m4LxyfvwR/WHx+5Lhgn
m+WOqp0X/6kJBSdJymULzj2t3tC/+6Edr/tCOeZHn9OC2phGXcl0eFJLYWqz3vv/
OYkgh27rJmJpn+h2hs4d//JMKjH52PxBXnRgN6STqO0nx9nD+FIS8mfGUSjA79HB
xXHPRaEt4S42MLvG0KjgUScid3VVxWNPg7Xly+idBI0tfm7ZDOudY/ocjv7Ssj/C
vHxYg33w7xVEYtU9tjDLqWT9LbxhnafBTdvxiNHfl0HUccI5A1kOqNgOByIKhp3l
cPTjWc5ClOccwcW9tsNaSBDdHA8Ws9VY9UpwJ4CVYs2r0uM9o+0noV8/uspy8FHC
TZsWwAYY/Le1DbDNjcOXBUbvW/5xZUbmNCmxyxNTrJ5ZPXUwcvuaKS4v/DBazZZ2
pnIyDQNuICVDNjbPJ+8iWIrNd/Zz+kUqy3wHxlW6MhlDI8CJV44ssykaEKHucnhA
5g3S2lW9eJfqdT0QmjzCIlSShbRJqDWJ7JhRAU527y005aolGYbTLqu9XDb5QKLz
mbE3V5VmDrf6v6pAyBmrjh/fTQrEOoPY/WicVOdt6yWp1VeasP+p7ikq+gaqLrrC
ucIISaP2uaasgNEqvEVGPSAbZo5WU0XqidDbUkM4j7X00Br+N+1/TWUPQT+HVgx+
BduZeyYMv3u5H1C+ofW4mmol8CRb6SCyIJKOTGwLjWfDGH+wtDxTQaMoaiA74Tb+
WHIB2OS73eWAzQZdR2zsMcJ8j/365AmtxLTuMzlVQvdBUkZLmW88cUo5LUalWicx
12iB0LdXLVVxCYQRvCxn51U7LxanDSaI+JN1OnfM2pbsUV7kUucgQz4B7uQMdOSL
UAN2PVbDAYRapWsb/+woopvDfJjtCgkniZMo9T0yQ+bPi5MaCxpl80fMAkZej1Oy
6/7O7KeAK19mN/HoSaJp07O5w1a1W1clU1KNZFw3sLoPZsaqnSxP1wdrZ6XxLCYj
IhArk01T2k/1lmEnCfjYmrQmbrWQY/PxOIWAsm6q+sA5w0uKmcFfTn/YND/H2q80
N76USgSC9aOogJcJfxtz+U6ANBHgWcU7p5Zxt6lMuSvKO6ATB8bQnENmY9eV0xd1
mCXrgctgl8WWPpykW/eByTNEGSe29vZYuhqH63IF0hq4s+/JYYQooWCTfVcd/wCz
k++TUlpkCRKEdtmgUq+2ivSW9ycSovbSrbNG/UcLY2HKvevZKALbVhnVzLqKrDPa
Tx7ls2k3e7oRoz2WDPJ8Ycb1IZ/kbhgMByAi1an1aHiI40s5qDZv+23KuqYLqqKa
bO63OzJXyeDLIsACIb9Oo3wRN5yljNrgizOnciwvzuciXxJV3NSrGnZ5sgApGKhs
2VpBtEr38FmNYhtTCXM41Qc8WPSWWk+RYgIyke3gMnX0nyTblfT/JwmyILzj0o8M
TISBPMlbHMy4eXLwfVm7lRt/HONI2U+8wsINweyBvG6cswuXoPTABSqzssm+bgRo
XuPkm/PiG3UPrBCRKyC7bboZHz6RVyJbo04Tby5x/jbla6BefvMkDd+0wPzSpZMM
IQNMA89EQUNlMZYfaA/Np75jHE0M6y/RA9WtIekz6VfTsKtaTzCqahqwOzrBBrA+
3FOB407CdpnCfkQR9p+7thYjvNrhkeLS7HeY5x4sekK/A/nNeE+FdY6szAJyx/Aq
pP7dXbXoHR6Z5OVXSma13v1WyM+JNidFdGcPdZ+MpDc63iwlfOgD45Q/DsUCHa4G
W0RtSX5fQHaNZ7/1jbNTFM0DQspFlCGCcxnarUp8ZY9xA5J6oYqGKMz06g/qfaZR
4OFYtOKn4nOQqVHHLRzt0mm3yCL/cHeF8TJGygfvDZgBiZsKPg0UyxH0K54bNqHn
x8rd74j3ikPz0vCcYWW68fALPmEVBEtTuRhE71Ks47i13WHzUU2tBxEUtU2TlzSn
2EMjV7MQ/cMEXl0uwUIDMin4F8TfcOpvFnuT+RctXa1MVRP/3u9XHmZn7QBT4e0X
40XCjPb2OdSmPR5zZaGp72XvOMeQr7tJNJNc53IP1p3Tr2BW/uRhwOUasKS7oJ5q
mEuezN8j3pY3YaTV6TFTZpK1EPe+cSs3v9bHmx77Hqtqj6xmH4dOBnAg/z5IdSSh
h+KLp/vTrToVM4ykYrGPXF55BOP465bBaz4gxp5T0qhS+lOimR0tyA9O77kZCMD2
r3htmyqABDXexBrdheUvejLWmWWbA8vgUsfTqaqmFAmmZDSpjyPLOlGAXVtJrIyf
ej5l1UpUg0qP+PGIgsDvxwewjouK+A5urVNjEJWGxZSujOEfQak4pSOXzotP4bvq
5EXUnHTr5e1nAF/Y8+fMSLT1fW3VNU5cPrxZXYHqnGO0DBJdjhV3wkGRIWYVvdS0
zQFXDEi+ydNsl69V62WQ1H9rgOK7OiqPaw2kBbio5j/JcX6jHo9e+LsTD0S5xc+l
zyOwQiWhFrAq1OwPht3VYICaqvvfM4Ie7InD49W6LXRDFA41VLnn33gjlbzJ5y1H
xzeLgsVBAXos+CaM/g2XKr//rEtOvsinNRwdvJfKPG9tEQ9yx3iSjDaiUFV0V8KO
CR4MOT/tBMRCCP15jb9ieTfvjoEUcc3nqT7YwiyulDanjtsKWaKWmG0O8EhPN/wQ
KIX9P1QLqj1d18X1CoqLqjnBGi7oc9i05PeMVyMdh9t6nSRMf93bAuL71KIXumaZ
QebZ8ah8B6shsYXep/u5BN5E2y+27gY3ChNahxwWWOxJEpUOgY24N/Ec0DtjOJZn
cZFRWnfvHTYu/mgtIMpt6tgHpqe707DNkse0gE9m8ZUyj79WyDDALTrluJRb/Lkt
fIERG1hA6UeDljcIHmfGbuG6aq9sd3s8fYDfbNlgY8yBs5A5NJMSHfInvmpYUJ4a
9UggSLnn2zQFGYzYf+eVpVgwK00K11lkkwV4m7yEKDHcLP9vRYcoK3NVychwotoR
/4d+ZA0WLPPLW6OFXMyqc5unDFyzZ4Qt2d0uz8kagNlLGsrOym3sHslYqQXoItlU
3qivrFH9Y6IRUyeavN1tZnRCfjjB7Mb5qoNOZl2bYwmqvKeO4OSOP0hEFIam7WnZ
/J+Q4x8+fLoJjaiWjyzTNmohC5z3p0R3iKZyv9QICWUcD9Y863Mc/pALk0qvuq1X
KLg26Bw68S8iZLKl1Z308JEBuNAGiZXpa9Zi2eOR9dF7AmeYk/69lzvaw8szjnDR
sp0J4I0XtXlS8iDAMmvkfml3q7DZ+JcYI/OxtJIAbhgVygC4ypwV4g8pydffU7oA
PBVmaNfzXX5J6uBlK+EARhPp5vhlxo/xUB4eGvnkrvNSC98+z7NamrumnlGlKpd6
j/iYj/4OazXLKy5YlCF2E4//WV2Osq/Byi0uSeQH7uMBqy/8FCK3Rb384S61rqBm
GZG6tgP3jQaC8L45cvhCXzrbtQegQf/E7YM9yOa36VEd5mHoEq2Qif2Lf+FLvmB7
iH6HHewAQtWKXex8+pFgDolK6nx4WcsalwbL+jEtIaMxpwYaJCA9TO8lceN91NsH
2oH5ToNeYM0mwIKM2E0fWb/aUCfOA9VaeO/rkK8HhMrUn4JpnC+8cRbA7nTGHXjd
mu2OTRGTot9bsmBoUuunje6svSmdKD6Je9THzXEUOQVe6OY6WfeAcfZwYeqJHGjm
Atn7X4MkLKQ8CtnrJv5d4qNfx7HFld519A7iIOP/q9x4UyBbMSMVq+AyVOVb72xk
jDKMff8AZm+LJ0gShFDhBV7d89pWLu/0WKFUqBbh4FS/oiXDuPdpIPuQzTazaj2l
0d3NbMVUSzR8ZV+ZiEgNxw7buy28Sf5b8kslFXOzZyhhWmsJVj/lUGjyZ3C4Ayl8
gJHSjuF7jFgdi8RnhUCh2dsAiXWoGGgo1Iw6V0HVe+Gka4UPa7S1MlPyn7EOyYuV
Z9eUPBTnZTtzF2/0T2WVxLRPgyGWlps8mwuSnppEhF80ssXWXLlWVe/5ZjwJt+rl
z+SZwrVkHgTEXry+GSqcuCkyBCPAklRX3MXzCNq6+lhzyka+LLgoL+KZOMFHaKW1
3avZ7fEpu5ZuqbH+oacY9/R/Oo+ocBaCVfP8ujZE0dv052TU8w3hEPz2v5wiVgQm
wL7EQjITgBDE5Z+qNeQacOeFEmBXYN7erNf0NM3BYyeLU0JgUzIBEvSw6igYkrSL
3SD+QX4gsXfKHQEB9q8CBsrZQ9LQfaz53BXfiuMhRMWH6n8UC+yxBQI/0J1Bq+rN
ILXAqal5hr2Y2aCORUXNz1qq3IfWszub+PFdFQ2FI5ql4/rYZy/FwVTsxCZmyBXw
Cmwq/66z6AiMyJiSfetSK0rVIX5OgL7UfAYX9eNUHbQUWk5iKTU65SVkzXMQY4t0
kGhBovO3VPsDv7eBIoioIxFGySbDHrSXmBngsmvxbaGjBoHr3pQzG1u86yMoFT54
2dSR4HOuN9JG+ldZLfFGQNowBfx8LafojMkad+Vu88wJVtH0g1sDTgVpuFtttfgv
XNaNr4FjqoXaUke8Oy3SnjbR5UuKov/nS/2LQ7uYLxosRir5s10/oL+Yq4ZnbmyP
S+qoOo2d77Z6bgXAmKmngNIGwWfN7JqClqCnJw2VsZVcs+pv5tgjxMtojZO8PHc4
lxnA9MMpSMRc9uDLIsO1Aae8Goh4INkWmw8+fgWO396el2aM8VPAMxNiFByJXvFK
311uQvnAZ7YOfCA90U63Q37bYKVazrn6virctyxuUyp6Lv06SqBgakIMCDU64yhN
XIGD3E4E2lXqkhjq4KgWFZOUtkPJ6On7VL1inSzqiFVXaczAlXOAl1QL7cmlmX31
ZVILt2Rw0aYPkq4u4i1Ho8tZDNLe0fLuC8pfOZqRplZ7KTHqHQoZNKBz+XCI04eJ
0ebkl2excxc2qpyeWXEXYHEleY+GWf/0RrBtPekpoOkBapm+eSeUd0IwM8gStJPS
vkBA7T73YLcy8HsYL41QALNIzY5IktollHnreurWg2hUU7+njIfd5cV9BqBK5x09
xEFQz9FIPF42sK9LoBaDoNSdzpIZJtaHwNf9jzsTcc6/FAHDra4QPRyW/ptTWCOx
qG5xQ/RPCL/xvjO9WCdWTyTxTqFE71KhyuOBT3qyhjbbtfl9fdE2w1ChN1GGXE1f
lieYQza3mjoyoqUG6H88mzpMKs6+RoqPTqxXvAWarcvzrPyJ2S4fKmlRh+sE44X3
4/HsK9Z1OaGMgZ8MmJSYmD9VUhP6TQ3qZTTtBG9rpTeYa0qF/FRizCTkVDEwUGoB
csCTk59VnHnDzcxzGbY+XNS8Vh9Om+cXCYTx4nGWpTT8bnl0AXVrV8VwC60J8S3y
RKigInGE4hmyoWejpKQOY2l44AhYEzPC7iTHWLWu9EGdQ23B9EHvh0iT8gMJhGTx
9dU4AxYxblcQkOUJjrmXsGDm7avn0GE+w7IYzCj0trlaUj5dNmBChe+JrU+wHhp3
hOK/UPeeEGms8qCpBgg8uosXyLWTYQQ8BPQxmS9tNoe6Ivl6Fqs62Llx+hGKfvH4
9rOukOLijT70LIlEBq+CqSYD5Weqtl6fOSAGgwExKCL7JhGL4nJFy11cVHxQBngH
YQvun9Fc3eq8cNMt2I7kKrZUzn0mHHRZkrxY7orMKNdd3uCJgiwhHSIzJBQmhdcX
W/bQph0JSKGcyjnymP1eIptbSvIo3hO6tpn+XPfSFh/Ss7wA+YzNzPB3UswUr1rK
CwdSRGaq76NYZrHCAVH/cWIN5o+c4Kj4AN9ov9fhqSWUNET3ydU9YEIJB+ZpeO/p
ZYBAahtL18dghl0u7wZ+RFgEXW4pbbOSM9coqlbXNJZjj/kp6Mrqs/0vU72U8rqy
5Odx1ZFeI3ZMU/FHzUMTSwkOChuq+wSDPxYObeNwuoWbRiPxzBoUnNrqgWW/0Eyc
2VE6fEC7SwaAF1BeUfWpx/X4F3lm3N7aNJIseckfqEG04C1wMkWVD52wuViQVymz
+J8kT/JDxzaMywoofyk9UO3wq7n/lESUtkuMjJ0y902Jne947kpn5BxJMuqcUDhi
194jkuZGol0uGAYDayL4mTZtaVqVFWB8xguSUDTTbpTeHV1KletKKMDmuEomNLWd
CoSbAF1v2vTjBp81V8WqMzDAyHY9+0FTz3D/z0dyeUUVu1ULn2BfhkSHxiPSKzG+
4Kk0tcycxpbTXw8mSEt4qOAgRwyTBroct8jx6yNJP76/F7HXr2eNMF1hNOv6/ofK
eeXQj7av85GGGABLu7a8SrBIc6sHr04feXAq6dSOVzrPBv8q+WPWCL6j0LUs80kp
NZuY5LdfIphguxbuNvmUqqMkEQfOyeWpq4qnlpJtXInjzQs3JzfU3lkkXjHbGGuD
7gne+Y99SCNVV2TPhmIJAYqI6VRLLwJeKeWm3wHsvGgUrDZ+AgXTXDehPDnsJnM1
bIsNoLEtLDGSuLJt4TgqJ0IkW6lWUX2iG/MjxDnDEKVm1c3AmOjUbGjsuDo3/R2Z
yBro/Q9OjR05Bbad4Ya0BxtRI4q0Gu2/ARKUkAXo0RKCEj7GNFP284KqxNY6o0EH
e2q9ZyY+U6O6zdPjoQqxYtOxZQwpv8oRkgw4s6pD7YHyviKFRGNfS+5Rw/fqrOyY
aYqVfsGOTWI9CA5wsyoJrPjW7p6IPHwwQqOVT6NFoVOs/HAld1wGKYTm1OdieDSB
GuRfhb7n1Gt04yYKSoKN9SDKyePOy5xjtcm1b7ollXH0PXWME+QCfj44yKrBjWaJ
RGbnsOGa+ABgBjtfPPhf7tyUd4U1jGNaqpoXxFB68BCN5Dks93qbcknlWdiF9NhL
ZE7btYxkisM6mEOu6HtvD9HiWvsrMKAoefb8s4IQ9Jd+KxaQaN6k7iXcomBP2Ste
di9/wfj271xMShSbdTd2aThW2hw+2BWhu3WrcCkxEsa/nxENNAGQbHm0/O7/0RIJ
/wB22MF4oIPPHLh2LrpHssNF3RkYC+HGT5l0wKkyppyakaAyT7/54g+5c4l96Z/9
SiF0ukaTDYnNGsTF19KPBEGlCr2skb7F9zB26AY+r2zk6PKSlhzBx9z1xLWNKXd3
Q8Re05x6vChmmlzvDxtnX/jvbE1dkENcO/cN7khPYeNziTRK3iHvlBYorqAziqa4
FRuL39bpqpyI9JPi/qRIGTMH/tlffccIfXaEdWUSM19O/wi0om3br7/Lqs5wOZyO
qOcsEqKWqOJ/60C6+riWP6ekzOFvahMsCMtoeJ6j+ddJgLulYBSIBtPpFbYZ/19x
94EkqoXSYVXP31j6z5wa63KAchWwTWURgS13PNoAjuVQmTavpc17CZiB04SxBWxH
kL+Y9P8ysUB75Yo6Obts/zg7EJydGUx3rlGkJ0PfTH6Az6MB0irZ6tap7FTGr6Wt
UqC57X4ub82gNwxzM61QMlgVR7WCt5dk293doxij0febxONJIRpPo3U/3pCSth/Q
z8p2vPvkenB8JzI9NNJrnYNzTK6QIc87hZWTSotTGDpg9XclVShIcN+6QPEgsKRM
v/LbTRVlEQp7GPO8Zm9Z+vUXAgw+m6NmjGvGkSQhlA6EsaaPqbt90lyqXHi27MCo
Z9BwN+iAV5JcglGEbPO4WiOk1N59oTZwLJdY5o+pov96x4fawyIcwKyAzGhEbLXJ
XD54xDKemTFfjlzzTZNpBIUY1lHNaogiuXV/rYFt8v1Fb4M/27hTHQQD9gG7/grz
TlchWz7Qb9s55pDvE7izGS7GyhxBz8/YG9KcZxVFEaj+cchYlttuXXgn16YqDvZT
mVyLwxjWUPSmW8lVSJxZ4x5JrEqTMexDgZmy1ny9lvsSQMCFNutGonDC8oDGYkw8
KxHhSxoOFpXlk5+N48dGV0PCqxrGTIySRXarEtfPgiI1YfTWCe8xIGsvNYbUSmub
JYukyLAZy2cHoC4Bpk8R/tlpeKSnIrtG9Y3Qp9eqvziZuJP9KXyJcCddrPueJfWl
sdOSbIiGVcfRTYU01Xs7kWm/aGfJ9CFYZ7SCmLjufHmuqQN+khdPwGA1XcMaupBz
j8aVIloOh2Tt/SvPAGhuU0wMxOeP/Kd1JjBpr9hMXaL4ahvHkxG+EyHF6FCmqR2a
zDqyNfrmtGbv3IDRGv7vAdnGsSDOD4UPLRex9ZvUIaotYKTBp2tBp+qMD3NoVeNO
HRH8tJrhuPzXI93l1ohG1+7CFySAJ0TgnEXaTns49MPboSIfQF+f/MqfvM1bGHJs
BkitFEPalPZ0f+IAg0BZ23ka+bFToiWZg4VepmYxhjWnj8JrfJK7mWY5W58HziRC
L6UTPpKGT+VXNzZvcZlY9+OSYi17/4P6s5s5GiGKXH1S1QgCR7elWnEcSEX1bEvx
I72eBmV/O2/X8HdBNuvTlJt+Xe9HHn9Cjmz6ktCn3X7GPTu2e/MgPYrl4w1gU3oc
IJGFotb92oeRqh4FC6KzDLXjkyRyDJcfNyNxbXO+3hk6XNFL3GbB8Hm5Ir3fepyg
9uQ/Gon3NB929cDx2INcFr+F/w+N7nFZjnHRgQgYM8TSR9ZyPOBvl9yKB1lfKQ6s
Tq02kzHxHvSoBU5jHFY8vlFwK+0ul1ifaOMugWOuaxDlJoUL3RTzJgyKE2Xjv8Jl
nbDZ9sPS2vBSzv0zBzUe5YlfJ8ZGY9iMQGoJmMyGvjigv0btIL0isVkoXGP880ac
PBf0oWQQ5RcD7uCayqWb89MYZVdrtMkbPVWSTLHrx7YHbsqUyPdLFqn8j9JWyG8z
yvYEogCX/GuWawdzcaNvdhyRhxohUoO35CXPog08/eUVCSmtnfC26wYhbrFgS0pN
jAIJ58Q2BLrcg7U9lFBDSN5UJHQ+IRrOxvwxkrGIEp/0zSV+aceEgMqBaK6iz/dh
SbugTTfRxhVdlHnz2qIQTc/SHZ0/6SNr/SPdMa+QKq/2NyPtjBclCqiut6PuNODf
Z0oeYHLFf5Hrw+zup66J6V3IgxjlfoW+oEFf8VkTnqaAp2SVrwX70sGPPg09aLFi
CjYGshtY4t3KYJ5thnrOg1g7xymQ+Oq2W5oTcdcoo5+WZ0Ve71tlk5zONmTrOAXO
UHPuxF3NtHoSc/rljZ3HgpLh7zy7Y7SAZCPb+UCh3bOSq67qrVyP647BGi1clMp1
Hi6+lYZI04b+VjH0HhU+VM/6xoJRxOg9rbww3jDFUmPG38LJyw6nX9IBk5nDfEEx
q2WQqJcYM0ZjZDw3oMPISHZ9kP3zCDKH/K0NYDVkhVcc91RBlVCb6ptJIVTwoxpB
aIKuq/SkostnmZSnov2xAKdbBRJ0jYtsFvraJO7yxOtNet4kVasxRdomzFh1N5B0
xF+nbOd/CDLd7lJITicxfra8iGtfA4ItNl8aRa0lz/yls7qK7QGeyWQQpdzaK1ml
VqmL50ASZooq6MgtgST0fbgjMp7OXiwrzs/B1/VROmaArItrJtAQbAmj2n7nQR4+
HnpYr6uWR+y444zLPIy7u0Me6H6BI4ZhS24n6pKYkyu88IN120HL+98TsCn0zRYZ
YkbyeIEX/Vkx7HLOP97EmyRB6KDtKiAVDcvr8ydLXRfJFVw1/upJgTy6Lo76EMdw
tRaddSa2i9m735sQZDcrzeVf+F+YgJs2cy1WZP3FMn++mJi+mHZwCp04F8AakxKe
/7shRMIy0YVsrdJMR9+6y9xeuhJwyoPCv3Y4tITrN3ifl1SKnM5bLQNeG0nkMYjT
s1TIj1UAJn+fGgBSWwoXDWMi/y3JzaR7yMG6UPh91tM3k8Kmjso6FFeuvndSlSXD
h4OrfgrZcg/1e/lblNgCbDAN9lCpL+RlyZSwTKmUn32OM4Qyq/PsUTRCP5ccQ0P8
IjQLBnwS+pucds2QXZnbqohgzqQx5tMRYSGfVdhLvwde+bc3xfcngayUZC1fNMfZ
sTkRNeOOdq2A+WW/617r0cFVPh+5JEIpNCbJweJd1bIs1BJVTuYsw0CEMgZwRa4M
voOSErJrnyU2HZW1y0m8dLMg0ggYykhNmyMKY/1329Im05a6XziEI/iqVX+sl8NT
kYtfnn7JAKq2p3AXjnk/o3NTNdpy3gjVjQNJgZkkH+J3vveXqxS6rGyoK1hKtlHC
EGMruuARAayGpJtsrfH79YgixgfPp4FDx3MIErQql7CfOYWy90/wE3q/JerPTVLb
JGpeEPSbdVCVa/kx2wj2qrelcWkq/fytsZ1WMnNnh5hQ1NGEqUyNq7sRo4LmWA5u
lfVFZUeUn/bEcfjIqXfYr1I6Kvi69weTbrNra9+dIyfJ2iSf15NrteVLKVs+X55k
HRo2OVYLJkg63fhk6GGagvMlveE5TqM+/EBcNXxzIMUaWHXouRqS01N8ZOnT7IF7
TD8pkEiIwIlVnKCzk16wiJqyIEWtBHemc/0aZAKkIGHKATOFLPaKyGc3OtVWMRqV
8ZaC40fsmEbZK/97HgtXqShAOhJM7B1hI+lzXTGsyjWluwuyCPgTpGBfOt4EbjaP
3Dhd6QfcApvwq4TkiD9lWn5nSSW2jrrMVaeggc3ZEi7Eu7aJdLO9d4Qtalq41ljc
BB0v0sEFVAnQ98Z733N5fsws7gl5u9VIv+uAxp+y2bbrzWjvfVSbTaDuL+iNlvIj
0lVZaF1srjh4fp4ZqyZZxOAWGXN4M5OJi+UKTr2ZGJU9J5OHd4W/EXup77BVIGwx
yYOvkFYGTDCm2DYUsMaMTUwocZ17XKMfJTR/n3h/Y8xEw0nI/+fJn6ntMtFoi50z
gs28jYd9QdeOfwpco5j1uQqcWT8rK1YYC5lCTJU2hx4dNqZEIHrlGg73Jtk/Cam1
X1K+IOgEuVg0YxGJqySRj1doi6djv79XyM5LGYAREPak3NxzjTQ6yfVSY2oNk4z8
zRczssnITRSH5B8FZMLSvckslJpsfSRUm5/fu/XM7mE622p9/t0FyB4lA7SJuFt9
icU46Ei1OBSd1N25i0ebqc3WspYOZCQb2h3r67LuY6qo7Auf/UgYomflz+NDhaxH
EqcjQ/74fiiKE+eQhsBSOYN0UwbDNVgw7VwfT9eb7v1yWvbR7l67JRz+2UzY3GaR
pCXv/9CbeC9Cdxw61XdXVX2t5rknyu5+/6Dd1IydT0GAWpX7Q6IR/ZK7yki4kU5y
Qeacy9rkwvBI4nnOk3h2lnLH+P8xhJB2Jsg36MkdtWgEMJCtPrkk8sq61Mj09NnB
GZMYPQzPFz5ISrE3nICy8UHexhg0S9Ab4MiWwBMsTOIDc4RXcNGvsTpyBj2/En0A
VsrDB1rCFfRX08jq9ZDUKSx64ZSY/SkZ9B0v6swtOR1kNKUgKdWeuGu1gnItW9Ev
BZ9NUv3KojautYlv4tTgWMbTInEnlqT7R3ut6WIFFN996v4BCAN+Ib5IURyr9C/d
fktxCOpnafnC2AmHLY3nR6s4EWZRCKG+CeqjcYwUcUcWtuDQW2e2myrft2htR5hq
XJ2hgTg1ZM4PEZO6M85M4OxYQcNAIRxSp9f6G/MdVR7VGNGCDePVCfFgBzHqSki+
rjxaQVn59TlCoXtvd4fEAFrPcjQBdUfWdysi5s19HuPIjgV6qr8YDYA+NN0lAM7X
f+c6urwkHSs1J9c/au5TmnylBizdx/vHcxbJ2FKNizJj4CZvl/2OpOCJw5YyqSMF
b4zgwDCl6yzRp0eUei0Xf4F61Lt5iSLpUIrqqiMPAbxFNnqoCm7s+0zUi5FEIuD4
EkTa3GJOWOq3cdsTxFfZuTQVChXS9KH+PPA/N7aQLU6zmYwwkogcauL0CvYS5tQo
1jpnN4EqsI+JcwsRS6x6aitFEk4Bpo/TkpIg1aorxfCaCvHUsaOQDUX/eVh1sZv+
VM9Qqk41KLyX1n8+OuQ2NXuRURG7UDuWhzuwnztmgKYBVFnoruT+gPCCPCPGNz9X
V+GnVjhE4cFONpezc6aH2hnop5TSUb4nEs8F5D5Hh3PekSn2/5QKdqY5ujImRbPP
gUvv2Xp5NZ5uACdZFN+XQ6m+K1KY02988vkAshwPChDA06XMmA8zU5X4i8eoEgpY
EdAgTbSmsx5X5Lp+QR6LqxsMiAw13lXEV+gnrs2mXUsSP3RqAhFhJgx9qRET3/tx
W0WfiwMWYFmO+C/aWYZPXyxGAlsku7ZwPYPDl+MV/VWjjZMfm78Rgp8+OsYo5D53
zll9DcYKvnAEs4vXzeKPVDhDqQhmPjO2Pn7Ovdn0fxeTq9dWvTm495Peanhemt92
zO2WPkX0QLDOH2J1yhmyX/cAzHfE25Vui4s29BnXND/d1uQKFFhQtMomH5CnCslo
t1z1ehHZV+Z2b+7oKBByPWzbnkJw20bd+gmE+eSQ6mzlwSQGAtnvUR84rtPBo9FL
S9AthXHiQ+/DJHqLeWQQN9nnOiSSxfm5zN6aPRgX4lk/NlofgRVQpswu+ypjg4Yu
Ji4sjcDLTaM6NiJEl0hHT4zYVCDAsYf/lWvBllfdRiSbjcUqAu6UWqvffW7+den0
8mCpWWa8cjb1ZoHnMndzplvXL0NCfCp0FM+wdpmcDXzuG2KxF6NxP7nfrc+kAuJq
mpwqvp2Lm5P1bUHW2msK7TtawZmwit+bdkkY4L+ahB/iH2EtGBBLAPEDAwdeJhMb
gxjoXq1CgIDjTWR9oO+m2tTr84DXfHJybjr+FdIKY8QTG/UA8FbzU6YmxoDQyqfl
j1kpT2RADBXUb/Rmh0NYG9pb1McSqTPi8kfV+aah6BgP59J1j0pPucww+YmS+fuH
pA0TFqFVewQFRHZYO2/lEc5PLGRVNchI/fu4Czd48tHqLnoxtjMg+fQax6ClBHH2
GF3cD2H4VyoGwrULApCi/FNLw666rzja6i7tkle/e/noJjbICjkB3ATTUm5kUGrW
HJ+/IkHnrGPRdq7cPidGtSlFNYfsHSRlyMXNddyprxItmTxy7XSPzfYfCAVN9A8D
Z28wNJV42/hCfBfhFkLl7onfyNEUwmW9E79KwY0wmwCSnGM5EV9p1EZOdFyutbPa
jsn7JqkE7UqoHAFoddQ1DGBv6Kf67Dq2Ciz9zL2oOYZg6xNDwp4QUyuxBbHllSQd
Cy4c017grjzQq+Uav40p1F2m7UZDTA1LzDKtJw3Rs2my0MgoDysb60eG5Vrwd7A+
WJVQU05bE7IYGPXIlXNUgMqbcy3T8u09hMw5nBQIIYv8d/fLEVc8OXTbaxa42C8R
IzEfVux3XC3KaXthI+dxkLZFpTNuq5wmoXy7FSVS5Wzbck6sgMelZws6oMQ6IxOp
S5NDux1SGRd8+Ao+3WDjgdjerN0XHbWdGdRVLig82hQUI+XYEZkMCDtLBW9OK7yV
xyjKY9B0gqXrcxLVAWPkgQu5IyKNaJbPAMgkL3cNLwzJ4+5deAOpk5ozxY6T63xi
Z9BSg/aRa38nO0SFNib7hH7AoSdicgqWBy5oy5hL3wLsOS1yqRa4zCvVw/T7fMDM
MlBLbfT/pX0pbg2Z3VqYl1HlG0qrRMKgvkkC/Sk9XRq/DUpuYtyp/HwNHoqUSpy4
E7KnOH4cphZGr2fwURrf3AcLo+Bsylk7NfVzX8dTuc4jT0SRYqZGJpLPjllUN2yY
lX9IrwHoeb4s5sz/GuWWaVXJadbG55BkFkiwD2vMZfvIsZnrHHVCASGWV4Nm/eRI
lzAup+vuoD81jTO2qrbVwgFXSbv3RCdJVLw5vfnJViebNL70eLGhvXskoK1I7oA0
vYNWVqupvPh6je3chxvoQZm4RCDY1itbQQZ6chGF3Xh9tb1K7uIIxMdsGzXmHesX
Sx/ggkkQSZcf44ZCqtsvBrxyM8ylDQuMmWrvuanxTKHNyGKeqscFjHUdd8Re1CoA
LsWNC02z+m5LWQMeVUUU9fMTu07rXXreBhfbt25zGkvAalBHVj7hm8l5usFH1s9z
IUlJ0OPs7TdKQAsIsUFfkSzF/CYRTsR1+F7kkzE+1D7U2lssJ2ZZu/a1kiRQbzBg
M6C4EPigY1IdbEHZDKM3riwAbxGazLa4rtd0F3gjxzAwIhQ3xJ9NhibZkU2W9SVh
zPK0dQ8dcYS5WIKjqjFCrzMiKv/inrupcSpIac+drMKIcjUbhIZV5ke66PrwF6pw
uePKubcW9XvKJeohLeooLIs+Uoqrell41OlFdkDhU1oRMFBU18kGH0lz0kP/28VG
2Jv5tc3IsgWCkobTa+8yYjAuXiLRT7JzuKZ8lnYtPBfKhYYZsjuGDqU0vOC9skIR
PQZhCJmkGjclBwVDIKiHMGBtw2YO9l0oVm/vkogHOQC3UCmrDRM9i+tebtvciJpb
yAXemV2TA9doLpMFLNVrLtgnyMwH42CGaFBQ8izU74M6SE32Ya8wGSDVXN5b4pSe
f/W9BubPwktJGNE2sy5PP07q5c+MeG3VOyzV0nE65lIRPzOeET/vcjtUgb63WhCv
87Z6QSqFzyjh/dAlcJOAm1/+LFLbdHmuaNCBX4vVBb823+qA5MbWfMwXZOLh37Xj
PWaDdfRDCNEVlL31aINjWuucZiopQxtH7TT/uWmU1fdMzM7Se9eFaKxuyTnOJ8L5
ex9sJ2Olk0QWC0Kb2SMZsS74id8GmQAwuEtW9CR4dEo9cm9+EPD1uzYWPWDUfWxl
tIJacUyNPOmpP7cKoLejdgAcHkcNXQyMYBvC25sg4tBh+22ujIy4AHCi48RM3SXE
ecdlxafR1iHmt6dzWhMVUh7GGDCyse8vky/ch+iia0nqd8ngxW3cIMKgzOLS7nel
Nlgth//CXEu0l9jDk+HMiTTjuKhOiG2tZQ6Fonn86usTWNoLdPTdxPa8SySeu2f9
zTryaK0hV69wDYcARJ+PatHC7DD03pjcx7hVGVDomI3ZlN24xQwJPWeOSuQhLhgf
CznZKwCzcS5Iok2Nn3PGun8Kt8l/FdXA5fiDgNiS5GyrkFXF11xBYo7lwFSU+xIY
DA01BM3wvsBVFDI8z07XRciVuzEWzfCDHnNS9zDbgCC4y/O/g9dXiASk6aXawZFo
3UJ3dCXollpYBeyU0kaC2/67z8i4ON08QO1TsOgVo7+7OeyKUayLYuM2765reAtT
h0tWePdqp9+W+L4l6XLdYcIoUMcb4YS0LzIlxP2mG8QpA+Nxyij9IpAyPaHdYx6d
DhvIrgPoTWL592h+QLiP4im5Ax/HWKsIerMNw67g/u5j6NuMWv1GrMHbJYWp8G2V
zpH6jEU+nsAgokBMulFnWVLxnysP8sC0OZu40iA5yyx4uCIxQDB83O+XeUQMwWlF
2PJ4A5z33g1RukYj8HHtUnUs7vZXiPHHUwon7HnrocalhliwcaJ5GNEtqj1Pbfh6
B23QJoXiyn3zMv0rj31SgdacWg4lZHhBdBXXCN/WqAimOzqp2IpFAVIMgPOwp4ai
C4IyW3YqYy7viqCm3kTcjOfhxiQxtYvXCjfnbpftnBQmSLMJMsqt+sUGV8feWHIO
e/AeDVCA//PfPJPgV8IjZZP/ujwkm5vb6VLH4Bq04Tb3jiDHitmQK+IsU0C0he7s
MEjmo5CvYglCnLqM4XgjdzK5ULTUnqgNsXGzpNh7ihRYc4BZdhaFgAdy56I4CJyv
tjGNzueHV4qEGGBlFyxDnaNTwaPxWqiRYsiZ9FBViOOowovos2ykY3RA0Kr3JFUE
XcWli5SxVIvksDpZeATyPFHLnQC9TubULSKgxyVuiGCIKCXa1xMbqsXpphwpQUs8
ak7ztdCuS9VPiBCT4lNYkf0A6dB/cZm7cWT07tr49hIS5mGjXDezK1oin4b9ql0j
VjR/1F8N9kv1ZkDf3khuMll9fzWQI2csIY6nv5Q3rOkrsMnsgMyOris3Ywr9o2vG
WDJYjc0hhexVvatoTgr8fdnYofrqJqQfa9wJuXFQxsKq+VdHrov3VGYP2Vz5KAVp
F3dIN4iX1okRg161hpxTFF0GI9j1visp5yoR0ZB6v8DNzDwP39EP6yFRu566nIKU
qgfzVH7N/YEN3WKptAgpak5L7dzI7f7QvC5Je6KNoK2TK3aEYmClJEmgC7F9sHjU
4WsblA/Mx2ACWX0EatXzhFi+aGCkmJTO6qEFNMD6vVxxGEXSqd00YFl8yjH4TyNL
Ji4MCrWnLj1lFD8/nNl1yoy5fjMUHUIc5R2TO5AMwboyX0upqVJLF8Axhv7JdxGv
Mmtudr2HM2ug15VhlPGwo5/lZCPC2Ai0s0Um3qmZYzIfg6A0OvofzSgoFDMXxFwA
bv66WPImzzeT8Z5hMFT/rkbXiysIzV9vICAvYZSbC9HwpKQguL55tayjtIFZ161Q
yQFdTYWMysd8st2p3VlVZWsljCIHilmLyuhiYlXHJItLlLUQQNG3pa6jk9R8w5Xy
ZOTsgOaluFyviApYN7moB4kXgZrcZ8pTUJxyWYSku6GXaBPdI/AdvJ7BVpBchxic
aih4qtg6obxgNyvidAGCsHZ0IUPCIYivCiV/qC3cN1jelFgZdUtU19g6tS1/dmRc
Q61fPLTcK00ExJOrMyRubq2MscvvrKQpGIqBl2BgydPzmXvAyyFAsd1sGdQV3TnJ
F7kAot4AMvprLlYwLtaVC1UCZwLYEAiB0pOrTETh4PByhER2H6CZrwQTBX1exr9V
XtDUHKSWHCin01c1NpFBvBfxzDKzedGglkhZQn/LlegDeSNlDo9KBhhihaO8PPeQ
3RaREKFRTE0aDFkOMzT3Xmx4UNKIMxxJSCd/VTxjd5Wc4lKFBjyNb+gKYBROJ2Yj
uy48u/s33aJEUOpmpIGwqmG/Uv6DH+YWyFYJyUsFPeWAq+aXOrlEN5C6a20MaH8F
mcDzr2NVAIkmnHaay4rVb7dvXyZr5Nn8YU+ndiXMe4A4Pa5WiR3v2a/cx/7clq8k
yghC9qzxEH6Uws90SIoM/sySRiG2v+a9rZDAMtr7PuGPIvEZcvsh0ZMx1W3xd9Pq
32QIwwIqkLResvIUAltruOdFKnaVK+8zozmRnjAkqQQuCxET5BnG/b3s4nfHDp+H
z30BMHX6VhrsRzls3S21E8ip21l0xusQMZKZe8X0NgVk3ByeOuoSrzrCItX5vYRo
GLrL8v6gCLQKbg/PmlAg+mS6W0/Bwm/wFg/1Rd9G0zz9S3XCVkLIJ5GMXLHpqF3x
toltJL3YlggCOFbFuRkVJHiUd9r5SEGMfVnjqSp/1jFdJlYjwXQkwbMb5tjHsXka
TVtAYSyyZ/puDYTbuRAFEDqTeNiSWcLsbjBR2WW/5oSY/m9oNVYHqQBO8P8IdOIf
yfQEPt+2cCUX94bYWBRZOWkK2Y11L2w/txFmdxCr/iCMSHgICgrIIWtRl0kaiE6Q
Q1ZUtV+EXgKWB9N91y1NhWlZavzTKVy+MrD8wGNgNmcMUP2CEB1DIdxEstvRozGQ
Nkf9gvQOtJVj1sM9jpDJXdcvRT9DkdyAKSAaBsXPV3cytO50b8IEh+6gdoTiBWiO
8S/lyAkMDLEwo/Dr5N+KNRN7DfmfqIylIjemlU4s6w5pnP0OBOOF7d7UQ4kAA2n3
8bx3W2S6h1D6jJTJWYOK7Rqqb2GEsC2fqMZ1g3uvyvPmMvksvwL98KS7VcHOIyK8
ak4/P+r9S0OnCIXclpdBfDDhFTalustOwhJTc2mKBDo5zE5qOjYt365Sq+GdRGhs
q/ULAfwuumFOv24rDwwI5heLNl9fThLF9jD3DPrYa0/L1cWXU+ntqffuF6RXWv94
ZPZ+y2JQRE1ytP5cB+3QJRS7anHNyJU1gPzik4fSUOOGmsVUGuN+PEugB49iiywW
qOsIAJzFJr3ea76q2sVe00G7vTCbhSAH0ARW/t8AlhwECs0gVJvkKmiH94EFi53p
qYJnBIP4cX3TVLPpnj3BmNv2BRIkM+qdxzfWtWQlGDjhPojeGh9NfrvjS8vDHxGS
zKb15aikIMLC6xu/dPxbd3SyU9oS9jmaZupe0XOLyd02KhfnRHMunFEHKcSiXepX
xibLrnx/sCuQu+5RElXZOJfP2Td35fGWdhzXMuEsCuCLZK++0d/Vr6t4jMVZ5uc8
W/FdDdr6Dz4o9In4d+ZuzP1MThmCFzWoP6clehMgT2tazMVam0k7osXP1zt617gh
62PPG0ENoYUNs61x3lFr1vw4/c2+05I01pzGp1sqxAibBaAefChrmzan63wXpb0S
G3E4b79zRE4V302WLMYX9CIdVV2OGyWeWZngv30xL71HZcwH3sYwU3/aRVH7x2Va
et5erHIWTurQ2KX09KT1BJSGsrrrAEHk4SpehVRb5L0cC5oAx6kDRlWzDev6UaPr
AbAmOIbETzdfG32gZ7XWcMoXKmsJvsPRcWweiEiJiLaolmtb+CG9Pbnq1SsqUt5y
3sOPhzU8yTOg3rWgj1cL72r0Y1qQxMeAzhtRFSCymeCIJjdRdmDbqlofXX4BXYUQ
ljGS2cGo1byGHoeqA8wDSgPS1wVMqB48e7yxvlKEhYtqXhTJ/+1u9+NRbjHnNkE2
wz1xyiTYx2S3+N2gPq8WPWZ9CZG1p6z+sXN6qdq7FNw0e/7PSdvKbjFdfLTWycJk
F7w7DMjop3z4APs45K5MaP55uj40Crw4EoTbGvTOTYJ6EKTFxl9J8bDf1izBjqdv
i4Ja81RwHVAckKhYzXnHN0d+zNvkppFKJ/CBO9moP+J1COJmhve/stCXWPNoNpgQ
s5AE2zUC2Npwtz17D9T9E6aucIB5Llp2vy+vLpR0ISFqqRlSp3P5TPJ2HQ5jHqp/
1mOfLZCde3pWDc/ig8X/kjt1GXz0xjBf2X9NaXbEovuGTDMRErF+gPfn11kq+cR2
AkIHunaQpvIq6llnLYEizjHzkX9cipUedHqCzceujAlpFtOwRFVSeLdPaEypTboX
UawvPbc9M4pzmUicphM3SJYoPTcweuYjUh8fHQ3PYz1TLdh92+PAZYZ/D5q9MZHB
sbvgGPzymwLx/H7XK6QBmpwobzv70DduV1TlE0epEW50j74Hv6MjE1hlfzxSjVmy
9ddysfZ+0l9rxFp4ho6ETIE/U51P5F9TauqWXL3nehjiwwb9lDmJprbM316Ijm6u
hg8oKYhhwU3iBO1iAJWhQ64KWg0vd7iShBm2229mbt8XCE9wkohJdiS6JopiKE9/
szNRpop9JhJLmDCnWstbn4ctVS8VWaEkIbBpYVGabiTU/z38aqZ5dwAedLPaaJWe
vsJj7Xc+ZpJbqU11rGnHENgEeHvjajth/OcFTlHpt6bCxTLiD2O2fbbDi6QpN+nQ
STEOuHFKPBInMYsats1LnVe0oU3/FuwEGD449FTloRTfNRjU0tGlF1+iLroJ0ECI
6RH0TACMoh+0uL4Ykng+ZGM+mEqO2caaBYJ5jbMUQVzHI4yHGN78qtknC3+uhMVw
QrwZliW6qVU0kK14Wy/u5eEBnrmZ+cn4TzElXM0c867BJdlTNjG2zxecaKmSbu6d
dVIhXvtRDJ7FB1xa9NyAZC5/h6+gfsPhiB0Far7yAVO1uj4WLSfqdbZZmIpG2R0I
aC8BCAlnlbtfJU3GFyd1JRMPJPzOJTuHPkuFI5Zp5dSjmLJ/9R8+eyvV6vFdZIRe
RLJ9f/eQBVFmzg++9fubQlfn9SIiZp6vq6U58kLPzw0LCu0hBBX7T6bTW5qUmT1R
cM0VeyXgN8JpjSVg5zOJEe+1QVbG+QUXD2a170AsWSzWL0HBwYe0tNayMpj6UP3U
zuKksqdvQK4UEPYx+iwYPHRWyAxzvrUl3Gmnmgrr5AcNIJwxyVTFi6JJ1ocqdEh/
h8uafIas8KFYV5dfQGu4UE5lyiS7WxGeyxoCY+UJv+1Bm5Cw8cC9DYtZt251zGdk
oWLXQXWNcW/Ui7+kpX+KVrw2Lb72sEwoTlgEfR7y3qtaq+8c/uJObJkfy4Tryobw
sOGSPrLQ2V7wFuHqq/ILoROx3lhVVnRD5pcWbWXFvkfPGZte4Qp69jqiXlkjOrS9
b7iRXXJYe2avrwBaZNuo1V+oKVRLvIBya7hR1RWsf92QrzZUQqbRvFdZm4EqzIhR
CW+aGI9AaDlejm8R4IT9Y3eeML85fRHr3+vhV28xiMa4YKhG2pjBwP4jg2F8jEQE
SqETbeW9UP68l+2LDd2umdgZ26Z822Jf/tlamQpKD/B+3iQg3olHbjhsgvN5ou1u
giZiFu0Kjh14lm4JjfPCUmtsb+hvJVX9lb44rrJxT2G3zlqWZkhfXMPvINYFtrYe
1N9hcTSbSb5CmMorQdTdyp7460vgtXdM2arLDYUBY1QmoejlI6IbX+HsguKwoKsc
Ih1jFBgG+4YxErMjHZPoGY4G9B1Jzy25csPoSI1qqVkFudDvmxrMYvTYOaJ+VDHZ
t9EZ29w7gAatA9CFqsyO12SSDt/s/9YTVMJ7En0QhdgwvJZimfqbJTrGT4O6L9E5
9XfhJ/QARskXn5LqkGHkfDIJVZuu8DMJ7i7i9fQJdL95BH9mK28TR6vzXAodkE+z
D9cKfC1ZwAE+ZPN5RqOdE4CB5F+EAklml1xQOD5vBJ//AlEBLMi0KD97QhYcS3Ds
jpLclW8zlkhoZ8tPICz7tLm8ekYYlTuostDa+B+m3jcoCkKltB7kiC68kSu2MWly
lWaxKXFBHVj93IFhZz14e2NE+6c5dNC678XTRCJN1u/kF2HEn8Nt/rVOTPl/Tm51
v1LFCQpF2a04qRqu67ew+zMNEVQy9vxaRQzMCqqVGCykHTp+AL2uYU4HjeEx8Mtw
V/6/YXmncjQHicZTLRkNG6Cfo0XT9xizo7IgnoIhzrMEfSqDVcwzMjO08j+AWlWw
jA3s2ucTlAtP89Ms+yaBPkR1IK0B6s7Dl0sZpkdY/+snN35V9blW9oiskepvXUc5
cAuC2ImZTpxCVoT9bmEF9XGogQ3vuxNt5fN6GilKLuGy7cPmukI+Z9A4UXDXu3w8
2nbYu07DyG+Px/F3s5ut9RctnXV6lVF0tpllgTw5+n8Vq9ssNfrxJSv6OgxKTcQF
QP+GnTwccrX4CsP7PNawzpo6ciAeQvg6NQz1/qaZT+tOQ+PUx53Bv7iUpn0ws1Eh
1V2UXgnNMUaj1mUej+2ttE3WJF52OEb/zhLgTlHlVvu4Bzwgoz6pKd7NJQSoyYXA
uTYtQHim1Dxwbi9l1/SFEiZZ77CbiwLOxMuMeb+bHTCqUqAi8UgI4a5TBPlWJoUT
TtPQ0PbA+mokM6eOBhRBvBG5n+IXe6e+7kc3cTX06ZHbAqQGXALHDecwpoIWUWlD
7YJl22dmXRi+LoIvzFz8CJfBy//o8442akbWYWLzc+ITgU42KGdu2oM1CiRNiTKx
sysNuJwPAWIShIeySOSdrpCW11rUCBsIb1zr7J6Ae4eRA+N7287hrUdZ/GkYqdHB
NPidKsaxv3IRJxREtLaN0S/+O++oqjb5y7HUgH9nxYaPOJ5rWarsePQ4Sh0g9Nc5
Vj+sh2HD2uJG+ADNTnbEUECpMxD/sECp5Q5xvupIjwrOzSDqMgknEFgcGMboLT9u
exTHfAt1ZbPV0eJWkuoZiLGnjRMbvJ8SuTogXZBXdjDMxw5vFo5N20+5GJ5UtLfE
xsmcCdgmIffNNb2PQR0nwN0ODrtvzjCM7tNYcCck5knTrK/qrxj8iiFgXKEBCspi
iIGjl5c0ryTAWY8cQoPukUkX1qt4RpWM4fmIsq1SNGyeutWHOd0CUEPlncTgjAwY
xUokpQ/q6R3+NzHaFJFDOcUuQbgoymEUPxpADPYZ3KapBBqXjq9qqNgd6YJDzUI7
q6k/JBnVRt/wvgYH2jr7Wp38IR/EXwbPC2D4wIvAd+smMFZwAGLtA4Rn3pR8nxOI
ZAYz1CaiNaMUzI4AXwSVv8RYn+5uzGn5b27C5RVFiRGddC1/I23DpOEWKPvg2aoc
IGssXakF99+5ojDJ00hGTH3FcRROpR0S1Wn0V6RZyxRuQh0PiiYoBmgcnqYAe4fL
TOWZ7s2qyoxlnQ944yd9rvCIYYfHQkR4vLUGwKCKIrW3Zey8o28eaqNnNelkGjJE
Q/FFBDvxkSBkFipt2C6/4ed5OdyXgbh43dX+p/7Viks4WPO7eIqfB0uw44rpdNXR
MiQm5OUwrNyeSaIQ0z1gq3FVC/BSAxPhn7URwIrFY0NAEyPCLl107fR86fxT3o08
QGOWLL7L0ZRjXzfV1ABIlmOOdhqEdbYx5f39exSOSicRyL4DuytzJ+CNTYOXSN4S
Gyh8Th22vUWN0VOewTWHFNkNZtx3szQkCbvYnC8ETzvn50WJa+CPVPk+/HvWCONS
aL46QmvDSn2/QNfXVPZ57nUAMum0W1QqFswt5DDcdgxSGmmn8vOEGeyFJ/1ped3m
FgXW+1uSKqF6OlE0hoNVjXByJIWvLo+pwRDD6reubB0WirHaEaZkzd/WWEHEWaiO
1sB8Jd0fKkagepmB0ORlUmApvNR7vYcQxijgb42J02MrNVg5LvoMs3vyynlS0psX
6V5kEHJ+t1mn7ZxvIGBvodfRX3Mvsbntju263lnXfPYCxBGQaVlvBzMP0ksZQecu
SrxiwNx2Kg2z4AUF6mfLZXooimzjps6Jy+eqH78dzOq7W5jDRZU8tZgNlqgmmzvw
YCQIQAWNp4IL1VOXOfcIKePwpgHY+7TKvW060JN+x0VbECpxZcYm0M5Fg3+EL7v2
swGdGc4Oo6CWQP+X7Ts4U6PO3F7RuaHfVTtj3gG/qkwCgLCqzUpYPQwUn0u0A6Do
uwAxMLpzBOINvVOqp4Co3t5+JK6C/1oSgJzZW8oBWmvRBSJMpX6dQb84N0aO2/PG
kiUuzZbddJvjbxiwKmVAkgZcfJyPnQqbTC1LfHiDFDgn2A4Qzu3Hd0NUvAFeZEhn
4hvszrmQdGVFrSpq7WzzLoeYz2X83FiZifWTtGGoqS/Tv+9OyDe/3DwpAMYhrkbm
iTo8sppi4bS5KIsJWTdDcx4dhh6bGuL/B4mxReR4NWH9OYCuF2Nv7mE/BieqdvHB
whrqJRna3v+5PLoYZcyA8pj0L5mHphVjFa/D9t2Km8V2CxmcVIRHb7S60mV2XZFi
AG+NcSaGsBbq9LFJcRCCbTwVEnvPymLGIHzAjET3qjUy+KsBRlZN41PKGmysZGtb
Bg1xlCl9Hkq7+ZXK11voZnSqngHzfpZw5k9dIxpVGssARW2ZL0+j4Pvbq0XOaB+9
vG1TopUlxPQCSJusg4K1n9ap9vm4OHOx7JMMrJMH8uyBS2dz69TYrHwVOC81mMvh
0htddKW5Yn64Kj3QlRGk9XKKaJIJ3JF6UUfbqtl/94S5uomrgEV3uZdAjMJMOLyq
p1LRM/+HabvZ3iKif2EZUZHJx0yU4sqs25ttCUH1HiZBz3KvryppIjCa4drfZQyo
F4uZ+kXbwEA1jVm8QGqQujOxLZzOhArz12WOSi54vo8QCu/0wwjQkpF2d/N++wbP
ke9WlWLZHMr0z+tSsVVoql3BKaTrbMuVcTNsQc6euCAjUxA901Ukg4Sa5fg+1ElZ
aEl2e5dPpcKhkNhDT5iDj5tzv9bTnOJlLPTB/d/NnOWdaQIszEga+qBWGAfgbh2a
WL/gKmHfI7zjIwUzBweii7M1mLBo9DMq6HOY+IBg8HaEhBlpcWZgtla+X5aBPsbU
/MYRu730bLP+4e7iPq4fKKFU0K0X1IEsFlj80vRqQi0e39jZKnd4YEpsoGOAZBRF
l5dsfSEojvWczZ4KlAFirlpt4ouPUjABVhEduqazkcyc9GpS2x7KByB8fbwqDDQm
FNmk0/v/MJwryRiM1nkRt5YDofh6uL/kGcuNK8xEA4Ga465Z9g2Xws7ulrVn3ySY
urujDAm79Af9iy4yBCA2mHdIgLPDEI49oOkRBWInzC3UNKRrb/0mGNrGrMTZT/AG
cMff/QNPMJZ4j9DkHzZnZJ2W+spBcQTWmYUkNBBz75PuI9lt3johkDzWEjPZ5jj7
HRzI2gWBgy+8z5N3AaAShUrl7h9Nsc3BKICRTuWteRdTooIRJaHsL6aMXPYKwD5j
0xw9kx9dcFfe0BwJliPblnwReUF5SbgoTMAlpBTiuMGcWlzWH8T1dapwrlnDrzT8
CyXamu+TLLOXqnEpKXDJ8Cx0u78wLQVJ2/PRx+iCk7RIx7zstZXV6BWtcrHVO36s
4Wn2dGwhFsOQ2any/oxUjVmU6rhpLpcNvYGCz5BcZxLmrpi0PcGO5BvvSmx4pNrT
PvB4wWMjjmqdhCxWookG3Ta3GOIFbum0nGoyiYddMWIC8GiCBPbbFo6xvZj8q8FP
4swv1hPhSxuSl5Uu82xBT+FcSBJmumLBXDgtYif5OQUGwvuIvjQvRhbAzdE/F1sz
cp4EfwgkgR9mkVhLn3cBWieJSl+ZkWhJwfGcEiV/RzCRvnVjC6+VzMVbodq6SKYO
qgg9APjQVc4wZfxpYVBZ2QtaDJ3L6JvWiKfUhM6PAnfn03cZ8qinGqTNN4Ornb0+
EckmbHMcK1d8USek8QhmgiLnxwBW2lISJ04Ju0GDikB48t3ybPugZoY0U/j2po5D
uxGFDxUhsFNqABIEurRuCDDNQSxsbdoBoRFU4dtDgpy6oInzFOmkyCyDgIonzO4+
2K58G2zVZuDT9LrAQHzxryO8vhDPk1Ad9EeN+RabBnPhB+OlJP0+t+sot3pqGaS6
DjKGFdEnScvuaG9B1IeVakPPoy91hIng7pf8I/yTZuLdVHjBVLPBvFJSwXT0fu0C
fmeRwHgGrGaiQcl3m6wKX45VfjIgzyfgaKVZ1MIbUnuoA1vqv8JUTjPBTLJWppqK
PO3i0wGSt4X3RmOOKKWDIu3GHCcbjOlGI0FXxW8u/LiImU+0LdCPyDKzvY3VounA
eyiWdz/2Qr38gtXaQ/aeGvLONCNbUL95BavqB06B7okrZslftCvzW9Xm7GOfK8pH
6c2h7LPFRcOlyDmfDi5IB6kbAIuSFoTxzVPs+SoMnwBZ88w6x80LRCGuUE9fGGlZ
Gw1NG5qfsKMDtrcWO1Ta6Wz2Qa/BjY0ucn7+HgZtOIhBsFwzneCpaH+Ul0//hXuf
qVSuzQYF7ET/9l387UpEuthoRM4mYre07epN0ZE9xW8lyjV7Gw0CeAQxKBqgfdqe
kanu967/tyDOYrdNT+RPiZChdBJCUla4CVJHd+yvKGUMc2U55zfrFywpm9zvM3+o
1Y4slPc8CszsTL4TasUS7B3ikiVSh/+4dGOVoQ2v+66ZlfnDgtmSLeYX6bMBEYNN
pNMWo6lPhQOyhx0WQrOq9/wZtPq6xaAcr9VLq0IcOQxuyMbcvT/h0wY7UAy5MICi
1/fXKSMyThVTWDEdWk0KUyCNHp2zCwHdwzAEpSdGrxdLY3Sq9VzE+MyRpSjcO9y4
GgJfc0RzOjVo2mlC6bqpOX1Jt25fdwsGF3fEcxK4NZUe3djKFlZdbEmsk4sQnRGG
n9o0oOj/PTdFI38mKIVeTDqy6Hpl2RSbifhSH80TOHEE+l1KGzfAtmP3NAf98kn2
XvJaU7ExdrQd/mQLGgHmsYR38Tl6egc9kWT8Z1SpQNzOiVic/g2k6dpiyP9EqoQK
kXAfRnEXgSZ2tJrJ6MxTAqdMcxhqCGVj8pQDWVjMCkp7S7c1y6b2OIqHRWh8nXQc
E56UqT0orZ8CyTgEWpzoTWwdtNn09ZVZkuSPzWnqvrbuwiP7CKrCmVketm2JAr83
Ocs4fbIY4WDH18q298At4zOgVELIgrboOkLIFPYhqWY2KU6OlYjx8OfzA9R93HvE
mz0sKZmI0RCDaT6MUPf2GIgM91U2GVSz8EJjZhwEPyErYpSrbvSpiUTjZTJcnSD/
KlPyZk28/9Sou2BisVUrAfMfg/0jtR+71XWy6V8lkD6sB0sZtWbWPPnLevH7X1Ax
FHgVXHMMjdam5wV9oBHDEuShKkChKt87L4zTeym/TekyXZP4CEMuokwgvaFP8YAS
TtumdEjQXCboJXWFHJKV/Nw9ozUF1bWHPCv4rKSJXGpmcapmmYZNjkHMRIeIi8bc
prcaoCvNqSDd6LXmx1Hu0rHeJ1NwTdBJXx/UtxWH3jzwo7elGveQ/gMEXpw0BU35
8kugYbUVjMtawTB0TZuajIjfawhiTu4OdKhrRGtfnfaKYUFKw+oZFcI6EmFGfOsR
mMRkpDO2oKb70ZrkTinkNwITTQ08SYZEo/fsCX7wHDeN6Wfe12tW9KMDB2M9Tjvi
UAMcc0eec+HSJogmrZ2owQORZQ0aEN+R0sNTy+po+Kuw3+ZwwtxmnUEs7viKG4aN
m5w0oWsAJt5BJr4+XGcfCFSc4MesNOBzRpHWcjcNc0ymcTPvutnOdCEgdsmSRR9J
cVrRZda1JbS+Ic+DtuvGZ14+DWJJG5BAMzUs6BgLBnXhmf2wqFSojKC00QhANmQi
BUatljMqxq2dUpkr6yvc9JXCJ72WkqgJr/H5ko27tv5LTdetsN3Wy/+7BCpcpDnd
iPwbsb5WYt6PWdfBtRv0iNk5Z8GuTnfSQAnGhneTCdgqsqO0iXvIf504RJb4MP4z
CPWo+3Iw/N04qSd9QX1E93cx9FemtKB4VdeLpjpZPznSsq+v+xJ7vpMcTTP8uIIQ
8sM10SHqsQ6ocnxFHSdM0GHvr7oxsrAzdv3HyHLPeA4azc4QStcNKsS4lBtO+aVT
4BxATlnRAonVFggnhIcz40fQgnq9WuX/cspIxcaA/5Zke0Jq/v1noDQzudeRuVwb
ejKiL3qOBq8OkUPIJM4r/KQYqvx7jbeBdPGiwGbfjNa01Xs+YszRE4XrjKrky4cC
PHqYtIuBJmCAqM0Tw/UojSGEUFK1gi5yvux/zxo9blD8mLQOjMIabZOy1M/OPG6R
cbb8UxkrzDbXnbfgsXmMeK5J2SgXBhPoZYwuUnPwdaEhvmPpQOC1PO3wpmUD1xBk
IJROHAi6uOVIeVXzriDoSEHPSHHA454CFD3wnbaO7b+jaozFm4HaCtuyVnkcEF6t
eqlCKh2ShVUUepot8vjaWPQS2Xyvbowx/Iw68OQa48UVScxHJ6rT5pq237ht6GSX
3BImstImkXJr5Gcoz7ajdd8tWX6zAruMJVpC7Re1fLWi0Y2SRXVpfXO/RlvXdywj
/aI8yzj5Rg0iqHeJUogWzjbIpql1m8k1oYUG7+yKFkqFrVNUjjDJxgqwdfXXfClA
Kp8iX2F4kgbKJDmmiXubYArSc8aPsJ+NgDbco+CURGogvW9ilNceNGIW8BrylZuS
OwQ8MCsPMVeD5TQDXgQGqZEFWf6E856Hysf0l8p+2HdV7Yd3y8gsqqBEFCFPRNQL
FfDgg2e+MEuRDBKQZMgfxcbsrzUVOPFRouU5dmP18iK3XZsPP2VeAuXqRuh2/muz
f2yjDeEOUTpvb3d+y9+aJa2VTWz/Ykjy/JLC4TSeU8Us+dpISZH72TYp+XlMTUNu
zq5F0RHGkLxOB8i7IMFA7vRUZphmS/VwlCz1HIURNPfzKZC6GhCcZrW/1BYK6rra
obJnoIVfNmzoowHUqvlSgMD9UqZPY/+ffLvm5oUvGI6fsnl2Ggtq/x4U5NpacN+c
xysJQLpQuu/hKO15s5L87k4iu/ky0wyBfVOeof8zI+HHKo55Jn7J51ap3MNjH90u
OkvgMWPsxJdIwpY4/9U/ve5/jdBrPbp5r75V9286klekHI6XwKy9V3g2DWCKD1/c
nxv5rkIqLsP/8yvUzqAK+4i7lraXggKHtRbLz1W++7rOIBI4yBAgTLmXRw/CoYrE
Z76NJS9gS0wtxKjH8cCJ5sfFFGgwxU+4SASwk52FsF73FbcC8lSiERI19lY9/Oyk
YHuVoHVb1Jvz7EGoTSSfdHv2TzsRr2w8qr9TcSl5fRoE1qUk+SfK8xJC3JQvmGR6
DyAGgEGT0wO8tlkdB4/Yiwoe8Y08vciBHtI7+Yofn48Ezcu5VgV2WVZBQ8Z6bKSN
ZlYcsguCMyU77l+IDKKYcHpHc5QggpdbPcJJTfFjhlR02JiHmVp/A4KGy1xyXybQ
OBh9hKKi79gho9grg6auz9JA973bPq0eWymPtSB86Cgjv7PB1LnkGutpW8jlJw6k
n1CZMyW8CS4LCpOBKMTYXlKTt3tfGaS2aD/bOjp0wz4O5799FtYJWhHm7Lqt1nFk
B/ESgAPjXSm2E9CH6oz1AjIURVRqVaszIt9l0/lcw6bRmWV1RLdl/xNWiEo+yCtl
BiSasJAxwDIOSnSmihVMEcJGxizj8NVuRKRZyxhtBAk2mhTViH26erMIR71YyDoB
QLAXiSAy8qWpNH2AfQxCzCzcQ0NpQ8AGfs8sOVym+Bgp2HXFrC11ITkvk8IYzYkl
HpB0r/+djO/kGDDxlC9/X7/rUSSKExeoud4VhdMV/52o6ReEn94ZZSEJ7O5wCj2T
aNQahulnFE7UI1byaLjuG1n1ZqBSB67qn2agSj3GBHAGyw1az9w7in/W1um6Au17
UmfKJuBhbR/ss/J816w/RODRkJx0oPAuhpvKcZviDNNrTUmbIf/x6Sk6cwpBrNJ6
dGGD0J44amCcvBLn1t2eXOy1yuQaho4IFjZaFcA4ijr3WSrPCRB5Jtr5XJ7d2vSc
LLiZJHlyXZmZsmg1R7Ufd2Md/gpuBALftC/A2HKp4fkJxUmng0eWcQ6nUL+AWzDC
AwgiAtEdN22uOD/Qi62Li9KzA8BU3HGHG5FA6is3JjEIrbD9zerFCII9tauHMHx2
u6c/LIuJPRcD4jd+On0xoz09p99IBedtL1980o+Mz3IRFadvxmkCTaXPyaRo8Q1i
hRG7O/PrpoNqOMbqvMFA+4+jGyUgnRJup0SHevLmB5O49iTTnYJWa7K8uhjsmxfb
acpxeMGhv8SSnSXj97ryaPb74EHwXgSpxkossa+4yXOf5D+tSWxNoBZglVIl2/9G
tmA4i8M8n+VVT0kAiLWUe4k9S5Thu0aAnTJosGpY32V8gLTRueiWSstickLtqeax
/VuhjJlIIPpDrjTx9bnzj1mgx1e0jKSfjzrs9Dtd77Bg6nsdL/xd+QRVWdEAoVXi
6/YKIBlFm8baaWUZeztYjdtkueFqikmhhM2TsZQf2a4AC0x/SkEUSYgwbcYa7ED0
VfG024bDKwm4k6tjm4DFl2MkVa+QUDFRUpok79lXVNukA3B7wpBdy7Lnau4zxnJp
ULuOmoLrCEEkBOTtJFLnvmHoq/IUKyP6obWxExCFjM0CjMzQ/KfK2yG+P69/rZeG
lqI6EXrXqN89al0Z8qmMXrpT6FxXxF322cjuhVnsYJcAeai89zEH2W563nT2Q0Hk
1vNbWhaKXkpFWwtNDV4SouwYmqMGTBR2s/HDq0VDdqQQJtjLvhqmMikEU8o5z8za
wCWB1b8Ch2IVdXLVEb529Qt5Iu1PDQAWH8654+GS5FN+vnE+RYGgONbdA1t9A9aU
niq45uhc+6wTH/pkw/DdvaVoaYCvcRXGnjP3D5wKQdI14gY1TMFWVFCwkkl9bHSO
xemRWqxOiP9NHkwmGPEb/bG7YHUwtlCXcJFTf/xQ8Js11awhZYkl+LilV632qNX6
WaZi9w7khM/ytBJqP+p+o/zDnXAHAWU0vBv2IX7vwrbiNo7ET/0NX+0Gk2VWagdz
F9hNmBBeOcGogn2ArlQ8Nhvsuk90m7nvazXm1qKHqiE5piQ+17qbIGmf3XYw3NiK
HQQX7bwRqkzMqjzOXmCr8EDqG7H8CXT0w77yGaosFjuem/VWmRZnfdTzPmhwsjUt
8pU6ai+XIPQCvxE8pS+g1pkzHADlgvSnf8FYckISFMQe5cthFEOQ+G9/8PVF1pjk
4XpDmcWVsGbEWiZj5tb3Ke9YRAo4U3VLbNvdPUSVtAddqMPaEgrek8p33tdMOITG
1A6URineaWQ9HagRTADsaB4d5wylDbFUZGEZ/BuCAw6LdDZ4Yw32VDyq2P39eBCP
zBvqPJ9KzVqnWvAT7u7OAA3/qulibwn25aZCbfgEsczIWcTjqt04uOGIiJae5HMh
ZUSksP9B1fjmRV483PK9sOQdOWtqobS0UJOQtnAHX8Gt8lxdpeKqKQ4DKQ+34OX9
t93IOByg0+9umFXc/hmPMB9jIjZjVS4Zg4vNvCCzNUlAYcCM5jFK16+4pkYeHQqa
sghEWcsfhqyoOl2PONKDEEbSqz6eky4G0NR7Qd88ONdT9aS0ZVd0ypUjqXIE4Rrt
oTUPWJ7bTIMWiIiJ3WAtYqjjFjDgY4T+sGp5SksDk1ABSt+ce9XYqKYodf2GKa1l
EkIpViLWQXc6QKGRsGjMkZTxcM2/oyahJwrm7iEeUjrutXbdxTUumZCwEwfM6aTY
xZZqtlb8Iwrfd/o1Yt/cnPi8xF+UoPVdd99tN58T9unCyTi7EMs0qvd6AxsFnhNd
QMQjDqG3Tvo0+cVZTgP3txJnS+VaVxxeZqIocgUjJK0JOxs7U8ETh0OM8+zmfVzX
/Fw3Xb140adxoLP1W7DCdYFSSwjdCw2e4PSJWZiD2FIS/T+X0UrazFPrFw/uPjuU
ho4dHgOs0QNnW+QHqpzapLbu6qQ27YNjhr9z4Y2TqyANm5t6CPyt+zkodGTtHLSk
ibqKidiNKfM/3eqRZiqCbneJdGD2rBN+fZdcmTLystiljxBJ7LwAfstUeCkjnFX9
88t+aG//TJ2U6LCsEV4XKsTpHMxb04yMqTC6KyXSweTw0SuLZm8m1X3S67YRYi0d
MXsX6A/iC6JfUjBoZT/UMcZQZY9q3lzkb0bNAD3MPVfvZD6J3e+ClUWiq8EIppHP
BbQNforwqASDLsewbUTx9rAtPQGifMGS3rET6wBypAl9r3jNQ/th/hmKjUO9re9F
jrkfyE0Ef61MEUIlvagpqh6F5aCi5BHDtaRX4h9PaVUYzNJmncvrs96TGBODWful
dVQaPddoCnhysk+GAUqa+yQ00Zmy+cmq8bE7zeRjzQT1aC+iTc1n52VF6SPdIV+Y
cD56oQm5gSNkU4BbB+bVXWCWgxPmpNQ46H94h252lqR0MAKCp6gST3RYHt5PoDxN
tpUfoxfhAF+9s4FWQEO0eIIP8UNTDBp/tft6JSZxK0qdKGG+eNrvVazHbqXwnM+/
NmxTq7j9ivHQ7hDO765nml9W13SNx1ghgwlr0P9ulSVnNRKGu48PIMA0l7c0HCnU
95V06MwLNP1jOTaOP32DO6BvtKyY4rzdFEurkeJYsBVn2VwfevLQPeK6QnUxPyWw
dsJdkVfIq+bGOGOXJXPTwNWdH8VbeTjJDXU+hF5cULK4xTGulLX7OeVGvsmb70jA
gfgrlnnXHXJ0Y8KyMRQWP3HTPJV3yZvBRpo8ftpl78I/hDKuW1a5loS41HlkqK4w
gI9wtqKgaKJvbiD3IzZhX1qLuycAry7vPcy5KFe8EoLtB2YosKXoz6sEh1IeC158
MsrD72VQvHwqpua1A3/xhXSCcGuFkrO14x3qhHJrPEEz7Rzsl+3Lxh4BgutO8+FY
5pgcmTeYQ8lh3tzuPtBYqe/5nKZvPbOEJ5lyd1xeTFZTA6SQaenWp7dZZhDNbqz0
DzhOr0P/2rQGyndzdTGeD3lkUnLR7Uph78rHuKMDrIqxwKSA7LX7m+e+7m3t6Nrq
LldAblOfyiMwGxgZh37Ee4z1dRH33nrnlZqWprXzLYhom2JZzywDYDYc3kAVbG8V
lekw+N6Le1QdjJ7gvFKyfHz75pMERePw398LdOBIan4UDXujGEqm9xqibS5ltEp9
rXE4Y+GPrAxHiGf6WuyiRE7QIlVojHPcSJDmv31aidJL7UeyiQhnofy2eibsrpho
L9UGSZaji6NTrRPQrbJGx1SNHSifrP2rQeHKw52fw8OGaLVxmpqH4HslYJivSwgX
em3p7QyiJ6Du+OWDYF4MmDiGwKqHP5KvEBVfYQZUe1U7XJHfnLGAtGIa0HJkAe9f
SNpeFB2lnqIilps34YUqLJHUwLLOhutlI620sg1lY25QMTkp+NATFHlnHcWXa5oU
znra/VjtyoeilbYbaF8VyuACW/VKXtuMJs6tNhu3Zeo62H1vmxLTzDAoQN9xCTLW
4rVBqUqEHz8w9hoRTF2uM+UB/DCZ3Vn0K75k8nG/4KLZ3+dTDq3kTElNi3hENO2t
Sb/tLvwf3slzCLyZw9hR1aV8sWgnoo+czQw4NDIx/MUf0koEM9aNiV8uQJ7lQMJg
OXtJlsKisRa4hU1DrwWmpzhVaDCCkDDwXfArO2dc3U/SfM7CHE2I99f4ufvcu5v6
u22ZAch6AmKkmeDwpLQSEo4ESvbZvt0iedWyNmFuJlWI8N+utODv3wRlACjZqD+X
glRc6CBuhnZrCQLqoDDb2gKp/L6jNHaEnWeDi/bFmo1YDHSYIXNdcsNci46MwTss
A4HxUZrRydfkzXMzxEEmYEkUHTmN7RZTM7u0iT6hxjrf4Ki7FuLpuIBQ9PsAueOV
h8s0R7GSY/REsP5q33pXf3N26wI6hjkLK8glmN4uZyIRjrkoJiCF6Dp2pweKZ0qn
q4o0E1Gx9ZrEYAIJhyHJBXOfme/YkNolQGVBxK1KfMMSUVG0tz055kjij3nao+eF
DIR37h5AA5pm4fxXEQCV/3oudP9cJD5srCGFKj5A913FInuKM4ep7F8ZNySaMPii
RzpzsCjAFTf4D2ciDu6kNeb3KMUfgX8p2YlpVe7K22UWozx0oQKcHhMSG4bt6z4x
TIjAbA5cMVcMvi/A7jmXEd1jf1Axlu5E8E/1MSvr2JXCKYK5RJ4rR2ufR/fo5M3f
WF81PqIkyVJO3pCVZ51NY1qmFhie/GCzwLOKmj7JtZ1EAzKRUS+B9eYuk1rVXSui
umGnaGTeS2VVbXdAsy7gqgmfXllJoLPRwYOKubx/ggB10AXBV6H7Gq5nQFZrJaEO
ZH2sgnweTnTAv7KpnZSCZLuSLJStPsK5cf7ldQT7OQPMc9O7o0d6vh9gRqkRRlMq
QQHf/xGXi4swCc4oy1gDHi9EpPXw1ppEy/3SIdQWkTNWDRnetj6wLg81WaoFnjDt
kAGmBv4wYIOzc5MWn+PI3G1LUw4Y2+l3ftM14Rb8EuDOSIV9i3/3JY5n23zZG/W8
adGmxyXvRckzdoub10Tn4cprPcPd991LKTRN09x7f+UwnoXs0KDttmW27CZ+C6fq
9xGxoQnBGRDDr4sV/tAlGo1UzvswR8G6oyyq4hLn9c4Ia86jUDpxcA48O+3dpRHh
fKny9Hgx96vxVGze8TEUPatO7wXNhj8aDyefHFWgco6owkTW+4pqvzU7/cYIYiQC
Gkv23IkuAIVoRUjwLVVnXXHyxNrPC4LFHqpZLrkGxB7P4TLc8Y6LHhKRLxSi1Wfv
zza+Rjcbgg3l2rtu0j5N1TT3iSIBuL+cnp/cCtFUpYGE6ZN/F9Uanc8MFamWTKts
8npyXqhHqh+nUbvtIYxIzyeHr66YcpgxqYvtsXWX/EWaze/SHtqnxOVxMkmmEc5p
jIlfHpXZ7NLADoRipC8chB/tUKjy/q0pHNA4MZ3i1pTdlt0h+gWVPBQhhLLdEwE9
TtfAkE/TzjFD8zcdwpElCczUMbbVtnPA907ZYLcAoPipG5kmuhGQxyT1jhb78Ynm
OLlmVAgZjxmm9PqUJ4HF2Ed3vK9AXibwRPdGCxGbZGU3o+UvAWUeQ1ko4r7u5ukM
SAFfR/ZfHNY+1RJnk+tarGpnAzOLuMEOQfyWYGY/viGNh1VCWgh/LuwjMV0+iA4y
/8dz70IRdPC313TeIn/hhkbZNx6ZXybIFFvD7wB1p4l91yrZJhoSiGqFcEdtKqQS
Sgw0nEzzKsx+bJuHBVV/4RFRDcpLRyAw9Buy6h0IESpW9X5gMj2uq99Zb2D/GuBz
WoW+vIuRrNGudCx6K7U+g5jp5JJph3cd9uZ5kGqnhsjTkNNZFK6IZIG/IncE8VQz
Ea8pNB17hcQjuefRFg+/2RTbYE9pAVFplDDXSEezF2IKyPc6+BYRadCmQuVgvZX9
4+C+s5iKktnOARQPPfz+gYPlxCjkw73n0tcWLh5eYFRGKjrfilCRNZgDkAtbC8Lk
ktA/gmQyGa816eJ2d5BBT+KLVCppVunKAnWSXaxRUBxNWjExWGKvC028f2eYKnBc
zetR3wjNCiyyeaMYECOZHIdxwZ1kvmSAIEuwZAEjh2bNxsFfvFkgfOt08hMXLIKJ
ltgdMikbG2UqFdtkolIexZI0oCldMmCLOsvsGkPbOlQNkYGURpJymKIi4Z+3Ls23
jNst0UwqT8btapX6jwqTe9v5JmFp5sMIUDVChl6ZiDRlakdqwwFKmcqF6F2tvKe4
sMepU8y8zxBi8tHhI8Kztnt64TSvINc5DPoa43FbFjlFxlQdo3MOCJvyYQpQWkDd
7tG7zJZtEGCukiJ9GtJ9oOEPhlvy2NkoABPg1Qz8vEMZoEknFewoWwmfwH7F3s+Y
E9dwnS/soB1ae47crsqobjD65RaEwbSQWNyjln3Fg/sboHr3X4Bi8pAFXM/m66+A
JdSXvqvuiKgzbfCc2NcFgaiIxUnyFpMn76G52+UPIx0B9ZRb7n/zUwWLLrqhDKTj
uUb/gZcsacYsjnTaWM3dpyj7MG1wfoUl8cuMJHp7/+nCTNsK+Li8/o2Bqvycg8de
DFIDqyQDDnzMsTcFVf8s0LBMvwBGBj3wK7diYdYppqvMc3ObpeD3xK93oJL/6HD+
eluMLD/ueu7yQGIK3Vew9rSF65pplordRF7B13eyq618NnjgrXgrl02iPinRV6m1
wL/gPru6PlU+QxBHOduAAW1Lapu8975FkHSCzGscB+N/1UAsuEV1Fpbq+V6rIE5w
pRmA+GxIju0+OfTFoKu+JxIYD8h5wlNHJMKyAbec9P16XoUzZ2QyUbUhITl4I5zE
P9makKg4eqN5FibuBSQR0TM67jU7jXYBTyOqSGvL2Dvgrnabhu6IFNh2qOxsT4Hx
LRVF47CuZwka9hA5gPen+jzZD7nl1KPQZSd47lZqIGsXSnW+2r3jUUgQpqwHR55b
fQP2rzkd4sRGf4sZL9NF14FKDJ5mg5xq8TjYoStI/usiwFhwAmcyZgZfPSBSf69S
HIuZ+5EGiJciOlI56m7EG/MTJSssyiBPu5k2YWVFG8FXRdoVN5TAQAx0Y3zM+BVg
WlrfryIZp9J+HPVTnYzvzoag/emgRqVzTNc4MTExxQ+6D04J6Y8hHI2mLKxQkaH3
+VldJ5Oju4eF0qPvG2+9s4C0RvbThllKvJV+arVwenIC4agCIbimefA3usFQap2g
OXCgL1xCvo9w41yL9rU/iBrAGsVI+2eA1xhZr+5YqAq5qC+oXZUpK/i5yQyz0IEM
5O8SzfQipukFR+gTZ7/6Wr+QuFOeHv7ixuG8yOfi3NZ6HwckXoMij7nvvfXQSEQF
3S0hJfe7QkfXoQv+JWkQB/LWT51xzdvwc6zPGZE2w1Ykdl11oVXfLerTNiu35m8y
AaOaWrPCKiQ1zy5q6RSCMtnCST7SV+0NM3AWFu+Z40PSWfCVEpfvQJUw69KvBnQE
YsOa9DgrEZG8B5xuHtiecs4aDD5r8pgD4208Re+fcloBUAmpLmqKy4JqjrEwrUgU
1s81TGjbklNX6SxwinNgE3oLbvLALsZOjKqrtucbLSBjYZThWAjD8+8fHhoeF208
aADnOgz4eH2Q8gn/FY6TDvhmD4KEkGlrPMFVqegulWFlzULfrJorQ2vgFip27e5/
6HPPMx7JPBjJ/eNZH7/16CuKB1yGIflxn3i3+/olbW9b4evgI3LZJIShChAk8+zY
5G1HRn8hnPrA5c8CmdlTy+Ct7GPGbWFQgv/cxv8l8/gONeOM4XLKHLFVotCJfwgp
QmGXhgNHRLpg2qxcVxwtm/pQyk6iA7GFoTQ6fNmuZr3OIU635aAxkvvQgDAwGMQ+
4edNWPWhTTkL1kJCav9cl9ZnJffR5cTXECEInlsEHSUH02GoTKk8bgU7781FZpxZ
04ldnBO6cAhMNsT9GjBzHnHjFoBk6jJsiZ1aoRjam9DqqPkTJOTBaFpw7h3QKmH+
qyQPX2YnW+yNoRxkuPG6t3IswlaM7Lce8glLWxt78uHMju4i7mFq4KEqvKedln51
i5FAJr3BU8AKhMaihE4uPfLJxwMN1YPllpiN8IU/rW9ka4Wi7KYfZoV8L8YI81jA
MiQiSoVvG0YDrZqoFFbCp7NHi7K7aezCn2OO6JrjmqTxzAAay4k8+h3HrkX8+7W6
8uB/FCPI0vza5azwVGJGvtKLN6El8Ycu1naRB2VGxfAy8Xs6u/EGdcv+4c7JGmmc
CLaz5HCDOO2xa+1jj67PT6wYWzWHPYPdFQ54KeMqVpM6LdUoyMqDcLF5dwqPwrrG
AN5vmoez9NXVWKSu5Zn3ZY3DEfwP1Cmfjb/lUqbo+p7MPQ2XX7L0VcIasB0JNTOs
NOOodA5JN2S52khwfxKq8C4TIdc68bzlhhkTZepsQ6OxVvVLRlUJW2WHXU5rAtGp
SKE8eRzSKHOGhTMhLMorVAPjkwRn8uNecy1ZoxttXfU1v8AY4Bun6FN2GoJT+MyG
dIedO7WTfn6jFVITplaFvpxgo/Zga8HqyiD835AMaqHS6PcGVE1TD/S1K0eoarxh
cAV48MxPcWGOoxK7RePNbgFLhvhHll17T8sm8FTEgLIKX/VdglQhWiLPsm7wGx6i
nXYF9lT0ClgGHWrjXzZ/B14NCD9fihjW5waaVWULOybFhocl03rs5nLdG3PdZY2m
+BAj2Im6U7dX9uBPopk6XQF/0MokthgnTTHBC3WRzgvZBciH+uW7vPBZbf+leVFH
Y2EeK+C7VfCIwMwZ+/pb872mI9f85Qld8IleZl0UKtfGomE6j3rCk4X0ECmDBwgL
5iChSUL4GKvJRmbE18aHLs+WJy1zUiFqor6FsDpHtOdM/a0Bc7pH9Qq2ebEJU238
xJ++D+kZC++DKpayO0RmfOgTzoBmLe3LkSijJGLa8qBWZW2idH3lYFIcwv1whxFX
/5UasNLrSd1TCbMIV+/JVA/S0RROtCPEaR7SjVMErICUaLF213gK9jTZ5Z8yWuGx
WEy+LBSG0Hd0VEgo8I6aFnIyibARAhS6Yl8emlnSYXxuQU8fiC44jcOEseq/QBWS
LBZx0ihC9VXkmN4GhEDBIC4IK6aORvdJqc54V9fWpfWOuO3luj2vPbn1D+LYUplw
pAqvLfHyfy8kDOraMQwB9dxNchF/GX6nY1lXjlXVpnUp6O0pZuvgjIPEZxkuy+ZB
WBgk2277aEnOeI+0ZovqYr80VyieB9BGRz8f6pVuovXduYoBgmWaJkd45JbgKs3o
R1Eoro5w/sLf6xAvY3bWCSevpT3qXzKy9RhrHrvgyHgGEwmZM7/g67Vtxy/0M2dn
CoDChleWVVTdMwj8Z8i7ukQMKFcV/hAtSXpi1g8hNc3IdAlPRk7QoCbH5w/CK5AE
RzDA3BeRUSOOPm1Lfl4eYUAG2Y60BP4T3pDmp1Fx771eBnj1qs2HnoPft1IUu5vR
4e1rXBGJG16M6UBjYFD4JDS+/InxZOOqiCVzBn2knrHkwnmQahAvlZeEZ2fBAgwE
UBQcBfZmFWcDATz0NaTX+5W0KhiD6rN7a1uqw/yi3a25I5SCERcw04zQnvh9fSga
lFWiBcMRh0QSYuNNmNhQOoVpNU+lBd+9VrHUsw69KIWZf7amaw2gZDEAwF9JyeiY
KKKkytiBRY2ebrouIai40yJv8HtE+LLZ6khv++VdENA7SM2o+7zw+EwTuyKNA9LS
XsBq3rugdtqDeEXQm/4VAVnknCPAYaLgVEDK38y+OBrNaRbKl0lp4NXrjx+kIa2f
1F7sGA7nwR3NkU4+MwW2AnOcE1OjKcCW0hJS6q4H1h19AZIwuViob47vk7J+DISC
jR+l3UgzV2BUqGY737zf1x1VggNSCjRz+/WUD6Qzcpb5nYWNaH4+IicB3hUVp3PD
f8JnIv9hqmAEdzCSRTugxlCZLUEjZv7CS0F7d9rNJGrcdfScNxeQZ01+bBKGDkKN
3RoV/v4umNod1i5WUsVho1CqGCwEwe5BWRCtrKbnS5E0KliqtikctTqxTMIutoOK
LapbFT8r54pf9HQIz9juwbP/j8NuGiAH8sKZ5l9EhIw7RPpqOQtVN46Jf/MIqNuo
PXMYHiitpq/QlZNJCL5v5wyPP+ykCAW8fAYc6CHP3iwhs88SUlZ533Wuj0JyT9xy
dBng/XS9e2h7uuJpJaElhWwLKKREd2S7karWtILsQkZmEZDQTlqqduP6iFBCQxpp
l6qHJi7h1oK8ei+v8LDSDEuSxYBwGWv0Jifcdj23dBX5iRsuyGLouvCF7IDQxm6/
j5wVXtQINytqV+2ROTcFlJfvDZXq4r+T+z4/w0zW5JfXRLuGWq08rFXka0fjBCgZ
Ng3/Q1SzpywWV0zJjcKPvbEyFJQVlrGbNOh6M1/Juoj6GkE4/COWSRkBTSyWHRpx
exmjjn0nd8o7KmLfxeKx5P7lOu9rhtfQvnf24kR01gNDkTKXLQ/3m5hsFgIEhVuk
L274ZZ3PpX/gl1FqoH4cfTl9DmCRskCeG8ybpszTqj++MDHKBLGy5CAkxeIkfriR
zyajNMX+ccEU+p686XqV2U0MOvExNoFJudRKnovdOJBoGwcZRkG6AlC25GC3pG4t
kV7vK7AJlKzi6Z0lfPpTHxaWMhK2TfqdNRFZhOelLOj0c99A8UET1lITnzdQZcxb
PglashNIIPlO/VD8eOaeb6/FZOOAYHOUk7/zNGMUXLLr2h9aaDAvr8HtIQECRTMa
5U2YDNjZPzj4GO8/rrneCDYtUun5E5ciYEJujihrlcGFWcU8mBvL+47GrEONYFT4
o1WaEUrXzcYQa1mtUQbc/0+CKwV4UWMzhKuHbN/fl4TZPQPphzt2fNziYBgDGgtt
3t2Sp7R3L7X/1R5FG2oSCJBcVKgG5gbc4TOWuIrdA8kPWd2tM1KgNlRo8UrU9bOx
E+1wMPatAk9F1e+uP6oejQ3XCFpiK24QZNYyV13JkAn4kY9z7P/xS2hXDtnY8q6o
j/hxZZVyMN4JXMu5Ldlm7c7xTXzWVeAmEJN2a5KfgpkmMja0L3BZnPZr+N4po1Rt
Rpid/q4bvOqSMl3JETy21EfIUyxpniJ/aZoN5DvelBEkWfASM0PtJsfuSlkPnQkN
u8naLbn8tPba0pEhuULcf51PzbZ5RYTySW3cyZpzTIL354YD0OfAvSuJjkNXQOG2
IO1n677fM7m+KfGNHETyanbJCkaupweOjl7AB4W8YGEzivaQSygM0/5kpmlEG0HK
u1dgxefI6uzDnk6+l/ASAJp+700wtPWcDhs1taF92NgCqi+s3S0DeX2iiLeTSLPT
CSncnkqj56X0RuDy/bKkuUOde2Ym0fXFsR1Brjx/lqHFOI1iutnuUu/t3JNaCbLB
5zFciXWKfIS9/PyQxM4eqIa3KI9sPCbbJ0xVtg2uDZOMqHBYUx06sycoZMMhDJB/
7kf495ZY44iNNx7sNVRUnR8X2js5CDgaddjathe7tUIVkZZdZvxNqz2kx925pOjc
BXL83gwZGoe6N8zuJ2y7xx8zWYbGzFFI19eQ83ESRwski7EX3bNMYEieYosOU5l9
qxk5um95jcAAl0YP4+IIMzzVetKi4/QH2BooET49/F6i+xhXa5mivFXBV7gnK9uK
xEJQgSms4rmeUEX6a8hpospnHWi5YZ/EWiyYeL06xndiiD/20dl1PsueC+LsNiDb
DI16zACtpOTQXLWZMHhVgJJL/FYNhR8Ano6QohZctOOOYtnr1Tnu5E/y8DYGikcK
6nkZK21+l4O8uwNZGC5U5cMln2sgSv7o8q/BJsZrE3jrzM3L2hJOcLBK4+n9DhFh
zZC1TndK95PthuZgQhbBj0z4j3r6//+j4+ckQK9S/71hcas5+nWBjU4+SUB/G8Ng
qly62zDDiyYi5G+jm5MXxyBiEDqBWYrPGX5cqBo8A0mZoJtWsvezXlzTS7gsDMvh
w1hFMGHcnxLrHvngKDzQ5jR/U/dwiQ7vBPaigdjmMPyMmgZP53i/5KQtbmOu8Yy6
mOve1dSElEEL+zgxE1/OYA9F2dJkmqRqA3KH40qdxPY+tWwrg1lgyxep9z565Or6
OULtb7bwWSl2BgFLFDG473sNY/wLPiSwfsyDyn8Rxjl209KWJQoMFNxWwOe+zn7G
CIOtNzC3BXXsGXWt3XQKyY0JGk/aekXzpaG34QAzN21R0xSxonLNbbBMz1+9JQBj
OrUNdf2gH+zurJ/GrGwYgeCxBGhknlXE5UR76MFtbtXQUBtVR2xdS6qtcFWzFkIR
hlhieXVn+nZKIrumW+YHTvNzwK5zhVtYNG0OyRcln56T163nJb+79CEMUIMUJzdz
uUAmSubMIxjw3R1vN1vgZMpCvCrIKapjY26A3d7FhLT/AZFEUiM5PAeB0v0GcWPW
Yz0J/IHZnM7UnJHGUrGfvmTGnT1E0E02X6JKd5t+IkxVIWpyhpv9z0XnwU7Ao98G
MoNclskjjRq1hvH50srjDTqq8uUmox1+o2MiZbIKiTnxQUGocn+ar6WVoxv66AH9
WpYD5z2yKE9SwzLEVym0+N8juPgD+MhuabTgp2exQGEEkIJ7ioW33N0fQjwX1qMX
eahLlBv2Qu0rAIhBJD1I1nP3YkXVPGWa38VPqsPzbX3RS2tKKxnwJ2lh1/hNhSP5
METsPJQsCQTOlC87LFnqNbG16hJS2KASSJaINAbsf7wa3t4L2JNZNv77ziSQZy7s
aBgE4lEF4Yjr+7CsaAKKQiZ+uBXfccLThVcI1nvDitFrYbmgppbbKVSQUFxx72cs
QPV6YhE/PW3FSu3ZYvSnf1zo0R3VXzkDySvxt6c+eHe4wFy99/8E9P6qh8uKJWKM
oZRrURijEPz3q7uCAGoEiEYUMfqbnlBDFy4vl3F+1lavp3WcyOJeb7ZYIuswiAQ3
P55cBJaJzW7S7HKVcb6W7EWliGYCsSZR1hlhvp9+6WV3sjDxYm2MH9fKgkmyWXGo
obzFx0rMsXf03nxUDImopfvrzSBh5eTDta3B02QVZA3OgpHz804wc32/HO5Di26p
SdFJ6oWyWfkVa2xXqDa9WQ+8oe40v3NqiMEzOA3wy9ZF1FsaxgwwUGN2mkjpZW+W
dnNDxSxJrzsHz0STpajpOuwc/z9nMdsnS/SCm/o0ErO+/4SCvP1A+ayq/UkcndCJ
2ahnZ8zD2APRj7VKek1kyzUmpIbtxptqx3lH3n53NgVBsu9CcJ0OXMNSvF73p6Gk
mtjube1R0AqjqrF1irgZN0zpSaZkCRPHG+ptNDJJ3fNCvX3nWl/pFnRhcjJgDcLA
CI457Xginq8f3P123AHdxxla/snfLgtr+AYjDdHswtgiBBpTu68foSWYqt/Rc+TR
A9XxCKBYhs1QspfoJ8cNzgK0y5+P8Gj6hX7wYiBM+6dwc8I8shfGOhzldV/POZBF
f33RkxdiyUnH6j8ydLAiZqRhw4ZnbUgh2qr2dtetkpv5E+AssbyNJNn7H2gAYTTJ
GjhJtYxYs3rdoHh2oM8TZzv00ecrxL3djweeKchY9V+orAlsRZWIf1pY734Axhmp
0gcw1Em7Idm2ygT5TKPh35Hu65fs9CLG7o+aDyeM5luNUsnUxSM+FFz1bkJGOzYV
nckRVxv9fRfOSQpB/hjNUlTS79S/m3dRKa5d0bA4FaJRjTAN1gTLAdb3gCsoa/hD
AnJATPUMeZgf4xktusnebos9rBFroDabuJNXcf4ciurLwXU7Mrw8PGkDzEaMgFft
fekT97dMv8jHn//CxAmaLLcKHaw/M/WeEBogdDE+UCdjW3BKagPyhBxdGzSWTfbl
96A/LaJb3BjqPD/dRtI8Wle+q0lFy1n3/1VDduFc4O0gt6u5VtYWMpgC9iGk+xw4
GPYDUZVUx+7SpIx893+RKeG2zdFCX/ML7C7A7c8kfXj+9iMBim7TRuQgMxV09T57
eTzSTwGTbgMnIN5fWgyL2iclyWs9y/PpiI1Lta3Hg6J8OonQIjfpqXMFxS7r+Ren
VFmFC2YhLXWHuRvxAR4EBYj6l6oR5P3BMStQ5yT0oTJjMN00PSTYm+cjMMWvI8d9
63ElTNTXLqCSdTpT/l0CyuhxMjtfnM5zYLKs1Tk+80NhYldrWXNC9ZA7maeLJAtc
rF8TWBQB2RO3HoAi59cQOtoucygEtcMdcBk9j01ZMNpFUazeQqGftxURP9P/Rj8S
nBeaFgL7izFAS3IiQm4V/hXSi6rv4QOufIRsZl80p/VpcBAcsPZ3cD5+zLvQBOth
zPXuumcyVFcVj6GUieT0BrcoA8MXbOwe23reChzAYYBbkF18Noa8tVxJmSJfSJzN
4SLL7nkjDHPhWVQvriBk8iAWXsCeFL89knSySVOL5tDFhx3gM0DfhFYRJ6fcs0AM
tFuC7n6pSr7Vxn70pKhVnHlNG4RITD4N77Zq8c5x0fAiB8NetZqyPdkksFplX8Ce
GF0klR0J9kDbcWWgHMzmjYlYvHu1CCFuKYyfRMM4V6tYxCthOaJltZS/cGyzaUWx
W2sZbnlhduLOmO7rxzjVoEk2XAogiSB4AQsyDJiprTPRP1IO9kBoSEOSop7oeT5E
y9k6GK5qxiR6bEJfpRGt8rpQAARLZx0BmVJTXguSo9sDcFTdnaWeDKPoLKfMGDP+
+qdiPD9n19yeZbT6aIAgGDHEIlEIclZHNrEowEJX1owcZqCeBDE83ZFx504jvoBO
/Phsjpwpv3lSx72AldssOcq6D0dCNPvSz5mWJHoH96b3Oy81F5Yf+t9f7oKIbF97
AvVwHuAk3TSEwgGs0sonO1Ww+/xHIwOm+aDUTr3D+DJblkXIlw4I/WQ/+laUKlpN
0kzE53T6H0s+rN2lRxrQk7ySR2XjpigDlNlW7KXmfL3YurBWC29pBt9TdEyAdn9M
jCC0/S56POzE3UJBuuR8CoJy3Py+31U013Yo1g9w4SZD0raDNy5DX/+QNwAp5Jlw
Eqc2uKAnRKZSbo45A8O0h3dsSoB+xeK4JIx9YybuOXGrElSDN00M27/v9RivPMS4
noeOC7QRgRrsaQoB/y6ayReAUgrvqHHvDtY/d2IoxvvTdG/gJ56hubyth4Y1IgT3
lvDPt+gUihLxf6L2FXLX6a9fOYnRZILwxv+3xlqLV9m/dq1WvzVvYX+BTkT3gCkk
eVzPrg0Euuwxyug7STlx8jqT243/8qQz4n+O9k5/4mmV40Hw9ZFhzEHGD3u45SNy
KPrxluDxBDnXPfcX/ThFIdSiLtpywMo4tCPw0ammAMbqs1IKqxMO8b2kLXAiS6qC
NQUvsVzhC25jjdJsGGTHtXyDkM615ZBig3tIHeyw5L+z6ZTqxQidy3+U5qLKmPdT
i6Xsu9t3uCE4z3N6sU73w6YAIGT6/2M+3QNDcqe3z14IahG+7pmcq1Kq47R/ih+9
2r/jzsO1W1U2vjh/7DNnJXOvW3FolCDJ9AWxw24tkDVLIJOeuZUtfIrKbfbyqUR8
u+yNqpLMkQOH1jydayMYOuiJSkFyotbH2LOlAaPZbC6JX4rAESD9jVZA8uPOIiwS
CaHQjgJloGydHUp6fxItWPiD6K4AGiM2Hef9G2hkzdbznhcgyQnSyRt3Jvkcu7SR
da/MESd+pXCmbURc1UvkzkmqixTfZ4KO/YWw9rhb+j5lVJPSWjMPKS9MIv/ZtHpt
GwFeO8T86I+Bg3rjoGvdSo4Vt6sW0VBzEglIyO8+jij6LmvGgOYOp4m0gIkAgE7C
ZwmRHt292JL4u/ka/k9/TzYmoxJuaxbJKNPLhUhF+buNW2Bh9NTccKIXZmtW1RGo
kH6n8ljjDd8Q0FXzcoacwN/PhXIAP5J1KqLz7s4fJtbncJjoWo04torxFtjgh4PC
XXcsKQBH/vZIyJm3T/n50j7eZTc3wW3rjgDRxlbiqJUbnvt+OWphswYvDFnFCdWE
P9FxaVm6FzQ7YhL+u494+GHFWCr0qD7hh+iUB6Sr7oIXyTcowkV6i9FHHeycxeRZ
bNMOG0YI+v9iB0MQJbBwVx+p+BB0Jb9kBJP+UkIHNCi/2TS/v099vU8eQy59GQTs
x8X3BNUZ2m6lnAlC094K8V5nv6CaR4/4RUlXSzJ9pfWTvffKdJs/1JMphnzgCsQm
gHZhXfwBHlUuOhDMmzU9eSOCoZqiY76WZhOni/1n4uXPgMjm5Kt2SPTiJi8KOayd
q2bl5CvSg87EIiY3QOUwqFQBvJo7dYsU8AuOli2DPCZh1n7E/gZC/RmnDJwM4Zfz
3W9Lyg5GBMHzI1stSq+91+k5ml6C1e7UKLw6uInBBnI0Dx6ZRLYzh1odlOiQBwEC
rQodLHNhjgpFximizUok1GBQSWLnfILYt4zVgZFi7D9FBEQ917c+h8H9Rf/D2O/I
7AqLqxAOw0q7hMZ/1ZBmVebJ/NGzasx3CtIblK7HerwUG8ZsB7HUCP60uTjuLuxH
uRcL2aQMrwrRrfktoAJFSLDgHVmZ4v/5c0f86QXUGulnoC+MAKrvYjPaMIRDoFN5
Zh2pvzJ2gHms4RfiGvyS5BjpCU0GkRwyPNSIm/3p/M9bx0pkKa5KZgKGpvTka/oi
nQX9MiOeG41MY1hPNFFhge49cPSKUK4VpGeAx35TlIoxyXt/FlyiMLvvYUf52oVm
Ue9WR4QlIGz4pHyHIzdhzi5IpvLzba1d0y2YA3K/piDhzQV8YJZ/BJTgU3nSRhD2
UMqOpgD6COMzNst+AMrIbIJ7l4W2/iQ2kPRsesG6DiyXBiHKIb6hUCAoRG0aN7OI
LJPTmnJx9LVAiloJrnEa2UWwDqTSjT+qxIv6E1/0+V4CTvbjcxWuT5b4UDK/RPWT
xOtq/tAujgRa+l8Onqo1pbMPvmKITHVgS8EpHFJnYD7VK49wVG4s4d2GoP/jp8KA
Wt8/hD0BZGNhEBUXcbjHVhWVp+qEeLVJzUrwCdzQNZERmkCyC90HeeqeRH4Oaebq
s+bPDNLtAAAlxUphgxJ04e0wSCZbnw4io3cY6uogCepQREBBT2RHkL9e4LCrsSy/
q/RP3D0XxAw+v0s2MWyAgsQE5hy/JvEmQyvrQcBxnJfTomPIpcTwT6UG/Rt1oYun
hPbwZuHujhbLDSdbZIcblvmhf2CItPW7t2zGoHzqDlW+e0UVypzT1pIpnf7GdbI/
Spj+yhG1CTEstZdsUjQhTIq3dOHgjs8/0klyzUnuAexUD6a08cW7NTEXB9/4riNW
nT05B1ILwE4sGBQEPX6T9cEC/7/FS454f+1kIKLFjED1yvUMx2AeWnWhflXez0VP
YPcNjp08ct//hl05jE1NIyg9cVGm99PcPQFTN/sYZ1DIa0nvFgfqdVbBB62b7CG3
+iAlCUKp0KbZ+KT5jpW56kv5wVEKKEHRcIY2b1l4bS7vQ/csabmDvABI4cbbUZ8v
HHObpVKkSO20zGnvTddsDBSP0z7Ai1IY1127QSKQi0Bjkg5FybQ2zXNT1czo6D4i
W6wG2eoswNpRqimcUE4mlVzJDJcITM/e/metPZI8oUJPLqOriFetuXxBa0fxba4U
qfjtAgSl3V+EFlVG2RQBz/NsyfR+h/vp35HCF4Z0TnGfIbSN2HfJ2wrEpO4pHBG0
GxDmQtj2eYf11YjLvQzi/tGfNbKlQGdHK+eihVL2AUiAfe0cLfT9TzJMpkafad16
muEYlL/sjVf8BwUMWA0M3GhQ+k7nT5itFby4OP9gP3GMOehW5eySO2/MmUEBnwHs
D0M20JJbfMa944nrw0VhJUApdkGnjUYednmVrNdj5sp2j602E5Gyb8QmVvi7ogMR
DDBr8GtIMLc/lXQr3/GPVhNma7MKP4J/HC+75AtkQFbZ4jNkBEugYCq2xeuvdTjX
lLS5xIEYrKEsOaslU5qoIt2VD065oyR4mJ8WeOmvoVBVHavhV7e1Yl/x0Oe2ehF1
k7Q5l0mSl9AwZeiyhBbpbrdDNxDAwTW2UNnJKRHLlwgF3vqZhirLDUTo1PzElaIl
34bAu+cr2qs7j803cs+MfuUf7/c62QsuuLYrT7DP48AxuSTCdW6oHsBcCUI2TZJK
Qm6V9xk+OTQrGdzh9dkEJFmNbQ6k3Oyu8CsA8Lqzma3UUfrXyREw+Oqmk+Xw12eH
by0jpAXScVdfal5qSkuY2cIYNvbbdoD1wWu3TZrV0MB4aogCbVPHa10dGQ/lvBhr
IGjeDxqwl3sSpMWi/H/PFhQavOaCjv6gj4hglB5S4eb2rqkfCgOwru0Kck7YpqeV
SQMQW8rl/almH97eHqkCDi/2rcUJRVEDBo0xldAMVsaThE+SHeOfimLltMto6ZAr
5qRDi+AlO2VRobVVxk//P9aTpaOzj09Z7PgCjkL47tdgWpwOjM2Y7i1uiDmxyCjO
kQiuDVlitdjNFhF1OEGSLAsoBTRqaNDJq8eeayS61SJBiqeSPNyd40mXaq7xIqY6
jXe3BgNdPx5/MYjDidBgPpaqypsZ8s4TSQZCn3O3ki6oXQJ+kn0lsfhgqXC3u0LG
ptod5xzFHFOrvSEeojU/DQ7X3784/pWeU28m8GNIRIohHg5TcApvRDDgcduBroBv
9THyat2QY+LWRXUF9d3WvThCHf3jMRtcCM/NevM0fYUOrhNrYrCecteVBGLELcj0
eEZta32ACLLcSSRqbqzMtR4krcMi+YL+TQHImZ6Y+Sj8znIO66JcH/kPzhqHtgu2
lvS/bURTkiFy6Y5PCUHHPiUAg+qv/TWdobaPsWTGeg8J08q8d4Td5X0enqHd5glK
BS2sywknFDNWls2qEYfpIYaxBDeQXJVgRSwn53IV9RYCHFfzoxf8vyStp1MmVwcn
H3Cs6acEYuL28k9RvfrFo5vuC8cu55yeOBxjyHg2Y8ECYhHzf9m3vqJVR2teYwzp
BFA66hG6hhzZ2EJJI0kuziBObuG3CbS8/86NDnQ516xgwiyQvgrQg0LdM++VJJ0c
JRHTZ9LRnYXhlswk+9yt0FkjMS7CkhVy+0vmibESUit6o7XYLnJybLqBU2M5XJQq
Cheqlx+RoCd+aa6jvMDldRcr/AhoI4uFtnZcfFb0dcC8jdujLeod8/Dh7qLDR1qV
6Z7cK8FjTm0naxD8WVR6AVyn1+cUFXUdlf9lN7A4D7lh1v9QauSpkhwp3v5Sp/TJ
TRry7n0iaf6J9OAc2mMcXEQR3hRpBYOpv3qAbmS+ji2sB+v13XMfu6GNDy5ZNn9H
mUUzBqY1Ua1qowNlxAK6Vsftr8TPy3bQ+vOYgvAZWPxiA8IystlzZs+U7OTn18iR
5SnjIUNPz0Q9DnOZVgqW4zyBMUdwBA3nRbimV8axmm+6Rur5IGNaYXusC8PC6pNn
JCl6EnYc7fWlLZqTuwCfSx/mlK8de8cmlXKDKbyervCmev2wShiWIaay/7qpwdNj
qZMgIt7u3BRKwHBKbqnxQeeKeAO0lQHiZCnfADrE3AmAVvyYLWeqi9TAla75Zoqw
SXrpeiWEaPahPXHEjkndeArJU1r0p7EAQKh5eCczy3eC8QQ6WIltGo4dc/o7s0HR
ugdVeEKnj5C7c/se0y88NKSXZJjFWoUfoPP2ygHuh6aoi8YHLrW7nTbwEAHamw1c
QXDgPdv5GkcpTAfdncYTxThrBv5dHyeDXq+8eaCE7dUWWH3fenBNP7gsLjGgXwmR
rFI0XNZLRx5V13sAR0SNEyl2qSaiwNX/v06loOAOvOKle9NKekIRlYiRagPgvu3i
j6JgCvlWWcs7p3qmcLOylooOkzjBFB8RFYQgP+iC708UFkWezoRiSzYNkAKI82lj
8LWV98X1Ylx9UQFlqTrJkyktkR7dSM89Z/TvzIA2HU80n1ebmIqfKuEyaj6BMIh9
dKipwZrJ9x/qMz22ExE6lp1C/VC4t4SIqpdheWccZXIjyPpIjCBxVQitPn+IajjI
ODB0l4P9Xbaf+hSZH3s5Fwtd0CS4x2NhJRI8SlrDF3k13yhQdYuNqfxPit5EQrPB
ovNRN/IKMjphp/WCRFmE3SoHpWYngSIIxNVFJPoyqljsOTQy89f1ztuvM/hYIrCU
z+n5b5LIFUvignsAtFYw+oKwHIsbqSuvsuhIF8jbkJCPSqxQdQmAzAkbocrSt/XS
B9BATl3GAdq5I1qvNcz04XZnbzQrZhQAUFEMzaoGVtEqCTs9OM2NWvHSVE3/S+QA
C8CmqKv7ttvs1BfOnxfQmHqhUzbWQGaW91C0+WNJKSvi3CSwM/w56ZkfN7qlbtUR
YuzxYTvbrFnfPQjz7tUErDkauGw1/2hO6yFLfnCVrAjx9EDZqN3GxTipmUdCPVJU
nOvM/R3FQpZ3jV2n1gJIGOf4TW4OgHpk4ijQ7MtYguVCM4E1JJLeuvKxruMvaNxA
XSuwhfE5qrZin3lW+fzk+egqrVOzDdhkpqIHE4Wt6adiF7koQDhsWHtcCNVBTIcv
EvRGXC9GqURPX7DoV19F/DViPfeOdL+cOda8D0a2OT6UzkGdM+R01o+ltH+lDjjD
8fLghmcUojB7uwDdf/6tOidyZa5+EDGDb+6k8nulsrqjayTY8ssp97Acra6pYBUW
1vl9VbMDDxL2+LavTdT4zM7UMcsEhmT9da3+QC4y53q81WdJeHo5uDZOxCL60vER
H7JdN0uC3Jr2wteyFePLenSC3wL4LcanBjxBKMtXD7htxy4W8SdVsXvaqCV9Zw9I
Ov9LaibNwYg4OhMhBJPSuQa6FGgil6pu8I/TBKX33fOegLxJMcdtmx/gZewusnVG
Dx7BgBJOakpbGSI/Af7qQDft2WREiUW0jeD/NaleAC5hz2hcFltHfGxgNzyG62yI
ZbvHAqyqsce9/FMipOJ9okNXo9w8aSWxoczC0DLB8tB838zOFc69tH5gEYp1nwVI
G3uiyaYlUS9n5hsWXZjd5DbRl4n8jqa4BoQ/W+sowIJhu5Kdx9tRBxgulgnlSHiS
xn2GNyc9+2r6yu2tXKUJBzs8Y/Z9wM4mZfU/CltHD4+uirW/vPG8UWhRJxsghANr
SJla20deH+kQtEJdtc0djFUDO4kkiJef6hopkAVzGGGurDGtjGaPGCAYs9/51C0A
4C63vGPGsZ9L9d+te+EkNvnA/qQxqnAluwDrFnS2b2qjYoqyubnlgAKy3RNySRJD
lHbOCXwMd6QAa82SEmBdoQwtVoytNIYxu9xKWUwyhQO01PyFpRl6aHlTD3tjlebV
Cg8m38Q1tCaiMUIFccH8XbyVWZ4NAqq71b2uOeNdQMaNiQ8Aaw84UVMVN4LQZQO8
mH3VDbE/gMquFOK/IdzDyXG/sXLlzXCMAZVlBfDvW3kAeJSNnNvRSacmJFxJF+nS
/CreIOKEKbc0NQEo4oqt+UVsewDMdG2kSG3pmJeLtch8/APq3Stb6uTIAmioCvrR
P2ORUg5eDa/e3TEkRT0XXbKUL0/NPRsbAqFjnepTzcLN6W6YUyeKCITxjqyow+U6
7qdK5sf8yr0VzQA/B+C8Jme38Y4euT/dmiOpsCRX4NqGxwdDd2/azqSa9eFVmk8k
l+PCjtefzZBYPz7oAqhXo86u0yKdERpcpbfWPFbMsjFVH6GBxj712xuCoutvVJG0
YgVH8GVZDYUyGn+krCKJYw96PQnZ0vRwtk43eXLtdgaDx2XpJwrZV4bhpQpjXIqi
RvalD/SBXcUWeDFsLan52lajZyqhsP99y25BpY8Rzn1OV6Ch/BYuvwTvJFipZIgH
QkDysQriDGw1smb2v10wSmArexicvTp0NwzwdoFQnvO5DFoq5TCLLBg3FAFOY/0X
33+O/+xwj5oMDYxzoluvmPnoHe3QSTjgfI94VrB7J1kDRm3SuXQYul8J5C2B1NqH
yxAWLYKXIJM6TizmXbm1AoDOmXcSAMOmeIDdgVY/XJU+HR+83NJCR3/Sx424V4kf
d2bRYIrhfrXG38OveYt6Cosy6VhLcH2UfX/CpGz/dJyfhp+KmXYhvdn2wxHhk9C1
RZgTMooyeX+5tThsDXMPeaz1yw5KqYmv6g9E8jrRrusheKj/8OkzFZPvZi9djSf1
QmXLX+HdAF5qxW/mQSXiPJIqgg/yWGH75x4K0ja4wAhVUZELyEX+W9FYyfGCNfSK
oyoArsNPPlonwmWJCtjhfiswCUr7SPWJLHcBWmab6ztj20urV6RJL/gJ2Pfjw7Pg
MEpZ0fO8woYQcM6m6S0ejLhCPg8/88E0si7c4ctEiEgJK1rD0aW1WmVJ2oDotzGH
oINBo3Eoyrl67e5LxqEu5Kj3igXk11hkZ0wHuEBMLvXG19chuwMZs7bWC5h5FanN
0PX7mBexGx6wNg9MtW8gJruFoTwnmJfEaBUfn0EoJpvCBTLVZl12vi/sYDliIE+D
4jxBDLqjC5GdpJO+/zYO0TDbkzugdHlRM7ekpyqXra8F0hXP+vcaXffvwuc6qfm0
WpM6UGusKOguXTAPLGy1LyOqh+mWwVGRqqXGp+CO8Reo/95K/tyCbq3fi/VZEtPW
qDrPEoUBYCYa51VsyOfPUoxtj6sA99mOuDztlQHUIkD3ctqfxoC9R0et1vOC1jS5
vZP5JOLTc6bkcfhEd3hIhsat69lxj0J7wNgo7XWdL3d+bCxWTjF77m+IMwyOsh2V
2IfHZpS7o6+QwUNwavWr6IDFnSkNpSjDJXq4+eMm5H7F39nTVA6sM0iZA5vv/dPH
Saexb59tGNsUX9D/EsY4JUfz7ApOJbyJrHROvGfqvDqQlMOHvha2rj5v4ujCLF88
esI5fmOuXPIFAg0pWd16gvatZCgpdfHMLEhdsJkXNvTQmmtm256YkxUu9Q4wOZfT
UORmYCBtI3Wy9wkGdqMY1X6+QzWR7aX6rFFYzceK390EeekNOViYYWVc8dWAw0Nj
fKcL2QBjj0P1OJHBSMBxxJhMmKRgw0zm0EB3QBL12GpzfUMEDRcbWcmvapheYhnc
Q80nXiGaqx8an9wECbVHneySQoBHfLBF3BOPoOnTAGkFEPIB2n/V3aKJgij/3Y7P
Sn1CMxyUHXCGiYF6LYtnVVHqFVg+jksALFDMLg8lqHSz1nviYAO62iZiuf4x9JKg
nee9+DZMdiz/pxW6nshZoFHRca0Ejit/JzEKws+g2j1EBd3XxXaayd1YcC8FDk+X
YpKrFjrDCQwz0gQjMexao3zgFLHw3KrHbw49tNMMmYBpS+p6yveyPGoeykcXoRPf
ozP9qgum9bIeEg5IVH/ICAe5tTnXKhy80COZghx6M9mRTLpaVpXU6szz6nyhdwRI
Nf6L0V+Ko+pYH5viavwun4nu5e5afGDocuVhhrwNoyqCPw/jdFMs7BVWtiXijvk9
2xm3mHiN4lZQ+jGzOhOIH+T2uWdB7TubTU3VW5Hi3rYG/q2K1192P1zlrOPEcOfV
O9an55DVpPemtf8vzC+Bb8nhO5tC+1QA3jtnso2IIGLSs2qADOBHhkJuIM24OtKu
q6Kb2J1rIaDvlJFeoOx8rK5ORhvku6bUU7Equj/c74OAemZySWMsQJoHjRordd5A
eFZCGF/T91NnoVDpiAUp+yPal2TLAQ+AGMpwpBp5I0PrQ1psNtw7MyxyPq7jFRpc
57NjYPi9pOxrCz3lAbpJi5X5neSb9X9+JgdpVbw8G5yqg+U6F6gqptY93DoQ6vqV
+AtWSSYmLGq2HhnLiuniMGJ6BSZWYz692wRepspbzqjUxEdeHXNbs7jT7RAOfM88
GjGro6X02vOnvgi+2fG4PhmvsMlBcd/rQ5XzEE0C2kHMoC2ZIh90fx7suSV1sNhr
x3cIeF74+qmYimxanJsaJa8bT99aJ6QAlxKRLuIdewyQ2dn5z1ccaYf3GgrrGuK/
hzJIbT2slnq0/kvB4ew5YpCMycfmC4Re7ZzyRUuDcgJ9ZKNIPdJXs7EQZef+4sZa
Czggi8eYkKm7FA2c/OYxAjFehaK8WR2qxxilk7nKg71Q9ll1YDa3s369IIlPZvuY
XcQeYoK/RW475VN3mUVxV7coa3guC0zzWhlS1CFuWMk49OQxqdD7LycSaHgmodIE
dCLGw7fQqoL6sSJmDFO+9nkxx3XB0dwlkwkdNrql2sbU0yb6V9znALxzT9gSOrDq
jN74RPvAqDTaRT1VXiVWFaY/uzfpfl0lG+qNWC83bp8CKFXh55s1fHlj+YTHYMgP
/E2CfAniamAfx2OMFJqDBS4TIUB+DedhCS2UQvagllc3sVfdRbp5SuhGt2b2ZGfo
KbIYoFBDtrnyQfaXv2vfn09T+lfkpJEoqL9jU6+4cxNybOix9THLSHsgs7pjhw27
FPNQMpeWr5In7I7j3xZVVABPpHuegFJQMqn/uruwcNOjoWeIC3dvlzlab7kbkTWa
mQKolXD8nK+CyaqyBzviP12r54gsdZH19OkS9DoV8qLW4bGb4ADQilLouoZC+g6L
joxuFhv91/zy+s2+bKI6fgwnxBe4AbwaNgRr2xRdkqbLD13gbgYGg9wIQbOdwwhi
Z3G3figIildmbnqWhp5Kn0hXZDDhhNj+wmwcf0YXEpTmqQTNAIBzyRibT1AT5bm6
//dda5PnsTVC1oAvQZwXPh057jroY7isY2kVHJyuRO/lNwX7Ex11wGaksKhFog9K
uSvq2PMAnq+dy42wAa6BXvKP3qG+wR9cyoMApdQ8dCwdX1p8GGwl8APkCdaTw+vV
XR6YoUqho7uLqPPju/jjnOxX2yBSpuUIPm31HISA7BkOET6c8wf6ZNqhWPyt47OX
g+/CCb8JzppbPb1eMaQhCSmNnWb+wAf85nmWJ6Ai8aBJ1uJQY7vSzugBHH8s3h13
SXNmzc6upirwXUqvhl/0VKkwFF4zHsw50Gq9jVDwhts3K+UUpFKy9LmEtKW5pZMJ
7dLVW6aE3WjDyIBEXQzNEXO67cUlzVngB7MLUDlBgf8y2nl7TUadfTp9du1Mi3Ky
7sTVMxNEDygGESnvzlAaa78IZIEXoRFBtVzQXXavgNekRwrehuUlxqb8geBqPVxQ
RnTxb/Wp8agniDgNLprETodKy1d2qDeDber74Ft0vaLhd9Uev3qbvtjm5rNAtdzV
rMlS57aot2KMMSat7CSqFnnkZiDG1S4F7AvXrxjmi+0sDYS56NMnNDsgQ548W1BU
xUc59d097OlPia1pG4ptGjBPhmR/Az8ZJBhQ4KC+9jPTLL+kE7gUVJ94NWUfiuNv
T6HM59jVl/5W4dAr5qYoT8HMjPhQtURWG8n3arswu0mlzmu3SjszXwIJHDvZyHKN
WRF3wmO587vEUlHkoLgRi1PF7wqwtYpJRYpdguifUtWOTFplaDHmDxsC2SnYtnnv
pW4IlD5LK4thF6nAX6xJVmyjtFDz9giOMNcMlsV1s4C/KVxgeo9QXCzhbE2CuxpG
O95Djw5Osv1cRy+c7zw5Rw0r4op+ls94mDXAmEhtZAIgV23+6y2u4t5YX0ZZhQ0c
3/KwXHbclRyU69KUVwm3JH1xttRfac2GrK3nryW2ZpBh92QoqH+HW1O4ibFj9sjJ
+tLW2kbSCln6TOoMuyf+Flj0Wlf/Dc0vGUmPs6o2FAAguXavgRoju2gmz7Ub5otk
y4yzz37qLmInPj7OSYCeq/PDm58GTGJdN+O5zhd1U51sBvt0wSsejiXQ4Xw0ERHt
ZxblbBFU9epgIY15dKDRQtzA2J5fZsnBKDmAZRJmtLsw6WUCIpH8YuJN9+wRRTj8
8xkqZ7eLn0J/zmFy4W61jeAg0DPDu3R4hBH7q7rtW9jk5DPVSDXTCzVB48B7b1pb
yHfUpzpTldd2T0tcGKZ34l1P/7cO2qVv9BrHVRyBAJHj07zn+fStZArdLeScTn1j
x+g0GvkHUGLAD7tuNOr7BCY5UGYK3ew42Vi6HLZh8F7VW6h/XhHxIDtjaKd3tjhW
mBd7W8FmNRFSBbfxln280hf7PABY5MoUdnky+GJZ5eTlxPkbnluHmqJs5IUf4HV4
61jip7aU/XG2rQ5wnyXBD5Gyy95RJfJQsiVrH6JL0SDY2JxrLdkJDAoPPIWNupme
X23GsLMZFhY1RySzljZtBOHvXrCPR24LDe6vac+72QwzJsB8FQ/oIzS3JgJKtPC/
Vwgqd473QU8+eg5AQ7Ba+o+i99VOuZPlheLXbHrrXy+gSeRM0xhUscXauU/56ufn
EmvZuP5anlp7VhnINhUB6nGopHOF88vaepIHVtL5P472JSoIt75M+Clnc5NVUWKM
SAFLDEjXced0Q0/uFf05UWCcmzliB6hr3wfM5ZIoiX9fYPwEB0MNYKAfBgjWBxAk
QRgisJ3U9MQ8TZyVjy9UsKtau6pNd8Wodc3y5l7P4UTOY3i9i/MQ3fkpnsjPryu3
cqlLI8SaorNzzwvVSLhEvMo4oMfnSbhCA1Ru2lsejmCna6Gs3cN1W+ih07b1KNZB
PLzqxGHZt5Ok1AYCBAaRQ3fVnTDCnqy3/fQ+3S8Drde5SJEkUiPrdUAMu/kcTn43
ShxOif4GroCkj0mYoSai4fbo7KSNtt2cFXwolu/QyoT9MekR4VqmU8/S/gXcYod7
tKKktYZhsZvqmHQVvFOAu7Krwtz8fet2fPhO3HkitKhu6nMSx4drJEC37VL4u0HA
P+yn0wsQbY8RHwg1bGljaOU9LLep3uwD9STqpLAXMf06VJXMOHYwMH6OCX3ZZCij
W3h0akZdJPfhS4kV/CWgM9AB28qq7GvH8EGjniBaGrmyFeMaGMFtQHZpoRoE/s93
LjkvUJnfEVpHVRDwPL35FEdV8TO26KuTyjchJM4qBtv+E4LdLkOVypZeRuTDE5kh
Fz3S22Q+LvpXDcYXo+w9+N9l7H9cll5AKrZ0rVMuPnQVa89LawuaArNQCOW/j+zZ
rIMO9YlWOv8GUSqRZsDAHSXR67Kt0Awc01tEk1/yD8GXfV96ojoThBF0JH5IAIrn
PLhlzjCIMvX943ybaYHDkzHmQxVV5+Qsvu3zR8JbbDilzx1iP4jKPmr5Zs7T1WsC
HeCzJQb/9H/1QdivGFHpbBjoESr5/tLDI5YuP5aonymotOlchNRt4McLuJtgah4d
Ct6uTVWwxuI0ZBHaUBA0oUjui6i+TyyMNTyqeymIDvrEnvy60reA+v/7H8GMqbGY
WBgcj3rArHXpj28c/d3tQDRn0DVknVtmpZdl/+QMz37JUuCBdKuZ2MfZhFf/BrKY
asL61Y8S7BK3f74nskLERN1Wti64YGBl+PVorFPE0JwGf5m2XFVF+vqREkEfEgmR
nLOU4D9nAr1FHMQjgKjxLQhou1r3jxaoZ47nCpODV68Lrcm8s6P8c0/YTmKkx/iJ
H3IOnyWALgGMAdqbwf+k5HT/8Q+X7OuToKWNbOsMhDWRghYOmOwop+92qv1bMEQS
aXJBAMNchFQgqcsdw7jU4Nuol0Zxv/rqhnd36RW3c6ksPR8B5REH/xqlro0c0GLc
HFHhYl/M0gePXKQLMNxFcvGh7G0aHv+C24QLGJ8cAvmVyDxDGV7aai8dcMrVMPt8
UfHnOwvBGlWZ7gy/V+sNxuAQjXWjqaZ1R/qKxR/iwMfWJvy66J4eAwE34EbQqzrI
7FQzX+mM35/0C0kRR8oyooPv+nHr/NzppIJiLP5WUR19XU7XpBxtYfq31mJZJjdq
8my9l8CtHYvLzwYi0/uQggu77mKiOan28rHEk+lQDR6/E/wRc35JfJDKEynDuNKz
xmQaRS27CNPo1/peryLBaeJwVEPpVBAt/qjB5Yk6qJVkjEEKEDa7GPVg7JZoS78i
FRq+jiZyr5gXYvQ0YFGyke8Xd4ZrqC/IIZaWXeIV9Q1da0GkzERYV3iBc+JW3P4t
K1vBjprPoFMqLthr/MTT3e42u/Be0/bmre0SIlFwFSj/Df/rBBOlgQ5ExrwJSmK0
VJd6wZbvkXjXH3VSlh4d/Jpzr4XoYtm0pd2ZpCUUCAwmgicaO5+HDncMIW2w+01p
8Ike7AwRw8G488dmy7Jy10neJp/D6BTy40RMwS4sZSlNXndlfRH5krG/pZW3Fwjb
X40TWHsEnivhO5B4zbHLqnT+1j++MhAWqUSPjxYGmf5Y4SdG6pxAk4/8YccUNZG7
traacoI6gC9XRo6yIK1RyFPCge1pooaA+RZntTAMUEyXMIPZ4/K9DqCcRN1cacqI
wXiZuGhZsQ4I/XF4BB49DOv9OlxZGfXqdSATzjRtEtBy5Mx7uYgGdc5Eihks/j2i
tz1Fnlu+xlJyHD9U+lHj6Twt9/xtWm8ayVOVVkCpOCHujnznfOJHBaiMuBQXLdcM
W2h4C8/MdOVszzLe3pM61282LBisR7pgvFAD4lywVEF7erwK1clyQ1Pi29gtVx3V
YR+61Y+gAqM3poMx7Axay0Qa7ITk4mumR2ad0P5bn1mjqJzxBSSPpzcrvwUaDkI5
9hYE1Jn00y8z5HmLsZHIne4LfUOQoO+oUZyQBBOS9f8hNEG5CClyp5VMtqQ8ycSC
1md2vlh5tLB04mWl16xuTWUu0ieBuURgvGWvO5C0KPVMwxoFCAMKuDxrKfYt6OI2
v28h5LOqHZ+ovVkIqpy2daO9CHU1q+dyB4Oj1AsAIWL6KlwX1t3VNYn1XlcWgFbv
lXdNzKEdGFS6kXrWXCnSVlAczUp7ZcO2xQ+9AqBio+loo//mt0Gmb07Pz7S8ZkDH
BktCz5C2H3qx0KFip9CC0oSG1kvVhOmdOYri2MmcICUviym29urEOW4IbFOMELQg
a7R2m34faX8Tz8u+T/U2RZ1YFfrLSeA5LH+8h4WR150NCQq8cYx2V3uJVm+AYbry
onNhNoZ6H/Klbvt8bXDlZoSWFIhf2T1jP3NRSwr+H5u+1VASnbvUZnUAO4lC7Lgp
Je50X2dZNSv07XkFOQa6zmP/+00l6Cevn5ulOoYd4cAzBbmtANCmoAl9dfV4wq80
ApSFj0LZhWb3Dmf0bvgpnLeke/kRvOlfb7v0nsCngY+PMsH27fFZjvB8kQtDNARo
TC5KwbKI63AD+4chd+9aAjoYc1u9Z4ahUcaWmrP3Usubdva5mUQqSNm4g/zfX8I4
a4t8ZS6YNAUP7wihZyvF6VeUfg9DqvNruufGIuL2RKhCF4nbAqw753lPdM4ml6o9
5K78+FaXEb/vudwsm2IntDz0+P/k87nJ0MMRYDy7O8HTmygfB5X0u5yM0q2RbNF+
kFP/Y1fqhALWTfHbs5XJC8BlT8QPwsvdKA09sXqzaaRW5wWgCl/LVsOUfmv80eRZ
sYAAiGmCvIiwQ4rr9gJ1oGFSIYni0/rYo9cDOT2AsDpROis2ZlWlXPJ2hd8i2OnG
XyiEmqOh4dZMi8nz5UKL8k/j7ZUNL9U+zCc6hdeOX3jxExNdRzTEEK/0wdujJRbL
RTIfhYmgCsoZOdV+/uOOxeceZFVDZpd3oV5PkTeBy3jPgB8kGY+MwKObzmeaOXIX
kweGcvrxUz9Av9Q6WmUB0lnlEMu8XRxhvCJmbhvveJi3roMCinTH5Gi+u8OJehO2
Du1OCLBt7iu97J1MvewdbdRYs+6LiPZmeyLxhCLoEaikhOWMBoLPWl+Z7AAj3fCO
FGemkkM9sAGyCWCrp7fnUDORxsSqjEcGHlykcGlqAIweS6XN5vAsHOQO+biHxIXH
A8Ow8+GOZKZaENEirgVo0+RExUcm/KLeAdJLhtru3cTaLCRtVrdGdelPDGMMecow
0RwNjv/WltaymDvHS50r1uUYg+TQwQw8Cke8YVeAJasVUrRnrwLUWjxh6fWikXJb
sWENDoF3TBlOze9gbAkLe64GKJWKOCDfCfynoWwlD7AnRYu9XzvkhoLo3yAEVaON
CKod1SBgrMyv+EBI3X1YzDgpKFum9wUQzWHv7JWurzGJnG4kCMLfCpKyHjMx6va8
FtAB/EV+f2nuj8FvSYOpyO0kqw9s70+Hhah6w1lTZlx17JT5TD7KrXUZNwgAXHiY
CBIsLtaq6e93vDPZkDwf3Zuvq3nfXQsgpoyxpYy4zzXk5jK5XJxIQzHkGuKzviaY
ZdttLsiRumg7pA1DeSJL8nSMWFxngibVLnkiBZPyCyTipefatUGORQ/OBXSy+XFR
ccSoA2lnS8+BkhxfLcQmkMfi6fTgqsC5qit6E4LhgBWm6SIZnntpiX1E8g0E5ryf
aiWxhwIZ/qzmJoJ2/8v9KwZze1RVe8FUQAXML3EtsMrZzGuTXEyz/CjxY7oypdD1
wnNS6CgOFIZ4z1s+MOz/xYVDrcqg3x4VXyTzcOfOsJbkTG7Igq7BrLMPxnqvedKf
VwnnjGXAWkYetpocJ61GLYclZM4uVYAaNe0Ax/0VvYOqQCTM6yYUyYKeJRUKDTwM
0Nys3VSzfdsMWsaYSIW+vilokVRrErhUuQFnIafUBBWdE69CIdMgDpBpWoJm0szB
v8NyvSc9ToyIA/QPlNPFZej0VUS+9wRiW0u4FcwQxd7VDCoheBIdn4CoSo8x4VoV
4RJwuRjBM8ZH33iJ6dYFKsZrkGhH/mFs5L8PDICWeM80fWQoyfaF1yLH59e6Cu7J
6T23aQwTnA0man8gD3H6o4uYjzV0A6Bolc2BJMOjCFbJVZaWQi2/Z6jHRsWTxZv7
9JfYxYLSY9/fr1VacK9HOgb9RIzPL5CPv9bCpMwAMs8jTLmJXXg2jL6H/hYwbONo
vEVlxo2QgIu84ZuKFpIs6tJIqUqAvY9rGuxmXoDgj6FVF5oC4/Nmi+XLB+tSAfGp
yO4rHdjH1pJi5yCl8yL2OfY83V2Ss6ttBqMSrEcdhFysvcF50VgWSNxA2687jQI+
BJsbtGf9BYS7DQIwBW0/GBnU3n3WRtnJn4NUbWIXmx9JzD2i3AHy8blhK7F1LWfW
380ML3mh8PXYWf5YnBHx7RSuAPn6D+tDn3G+aTcbKW0wV3zGawmykq1Bc7PKBPWL
Lqh9Gxp52NQ6eGCvVHef5cS6Y8xqq+xPMqr0uBUXDFpi/GHI7mnYRybc9Kii/sro
8zGRJxOnZWsoy8GBuTEE8DStc41Hr5tkT/opqqoojtO528aM3pKl072Kh9zjNtMV
bJfx8KVwGl8NY9q3uWxRVOX297d4EmGXY5P9beqBRzE55s3BP9OJgX9nUfqxsj2M
q/5H01FIvEbhZQJt8Rhz0LRvq84bkygOAXHk4qjjc+MdnzF/EpaWMdl3yqasG5oU
MzV0LDyu1+269eDDG+hKuielYFjoZFZzahPmid9CeKeZhFMCg+am0Q3a59PNokQN
U3EoFAcQsTOuf/Ve6s0FEeHsT4t3gVaJRbh/S4g61bIxlbHAg6xaSddnd9sWCm9O
gut3s58AIyMrZjEdRTtwy0YaBTCmkl3ti7vbqdj7/I2GWEIn4x+YuSmDghOtmENZ
UuVJ7VMKLf4FM9Sf+t8WSQTS3Bo/ieFU/h+OfKTEE/3onAHpG3jEuTo9/hJvGVze
oFAAo0ZTX4ffTuit0GS0Fp7BWsFlUJfKweh5tJeKKUjn/Of53dQoNieCFPSkmR2N
0er4UNECxNVNhN4AYD7vB0f9iiDVNJClKNzLJPC3CfVOYxOGht5J0KIixLXNJApn
z41KNPWhltcmvEQ9xBMQBkoF/DVOgen4bj4yhY8n9H0IxlP6s64AvZcoeVFnre5M
fjSDvbtmfSAwaq/LQyiSc3C6Egrk3UPX2fznYdnaXkQfg2CNsdfpAIlOUnxTim98
rVBfQ4LsP5mKmru6KO4WBx0HSIQDGkNUPbvbLdFfQkYkGbn9BezO5znnIQ7MjiYN
quwWU66mPAueJnv8DMeVzfZqDmwtZ2ULnjoRjpchflwsW7TEAJ0pIbHbR5e1109f
CPKX+6c3c8lrpJ/GNig2c1m79HNRwyJ4Xt2L7qZGIa6Unh5E/HRdAu18iXqw513/
Z1Gv4qp+JsTa1SmzDN2RwlDnvhG67KmckK9qMwO75CxiC8UFcjH0FLULFAiFBwQt
8Tc6EOt3RstHh3PSl+mLz8etAuZfJXLui/OplH8T3buc5FcaHu9sh6D3uB6B9zO1
4dqhW43aeW2vybRgyH50NpbDRp13SO/qBsvvbSrqzYxgsipd1SVS7ZaYsQoJ5IOC
PXAwXrXUE63quXO8LAxjEXaeseeb2eyy4sMSDE7DAUbipCDpJt2o5vJyHOho62dN
Fcvy2mo8yRD/Tww40dl/HYvyLaGMglwL+Zwv0M1oQh6TzuqkajUEv5lIHQ79F8Ex
dFiREblhHOO8fS0tREKi1Tp2nk2YrzW4kxOpqzhvxMgHdpRot6FtNQ637VuCkC5R
I0/7afChnMPHWoIZxrWyl1VAEsnDQcawX9b6x3ZAiHYzwXOQq07CEazXwU7yomMv
7VyrPM8mo+rwesfFNwVeDmu0sjiDSWw+knGAO1pStZQjHcgHpJoNE4nCRUzlEEcb
MSzQ+toKxIu6RGjwMVMv1knwV9WmzntbZ/BrOsm6VhNGJsSe4LN2OHr9jleMXrUD
LrJaG41gPmRQFeZCcOW89tM7D4NvHg3Hhf6O2+c43SDFJMUdJuAYlWa+Cb8+F+OR
QIRNmS9g/hflov+kIfawtsQv3PPll1K/5tASadTp8D3guLP1OKeMQwMcQm1dBLQZ
JjAyUZtmdJqXsdIEyMpHDpQL4l0FjWCYuKDwJQVwCjnu1aY2fD5tuGOYtTGBhrTz
lE+pop64qcElFU7NFPC6fU73CZ/vAkDCWAyQ2vWGMnboZzTx2PSldwynkJnvOdBx
OH4eBewVC8RsMWZc77fv5nUOw3IuP4WL/cF5pEizh6n8nir0rtAxC1AeF5plSRMt
Au3ZbjTWChOVb40wsp/5vNBmDwazsK/0N2bkPW0oAxj2sblZm//oWzfD73KjksVD
7mWur4gWi6RkDwRx/q6cJqp4p1IwAAkAnqG/T1JU/MoQs64hdKw6UHCUlSzj0/TK
ueW1oFokhyxjC5wTW/DqVDzgVp+xGz8lgw/QXGfF8swnQG2p4sfAlPifRfWDQkGS
Am2qG2L2JxOG1ZOVIt5w/XR6SOJ/u7NmX6vW2zGECMyeUfDfS1VMb9LAFty99j2b
tbsBw4pPhL7QI4kGuunK41JNSNtpyVgKnbK4g8TE4doCk12cKDG9XnVPMLlBBdMl
deF7erY4BazpmtGoyPC8YXnUXYUDoF3vCMbSvVj0gklc4hjp6ghpUvT1aC3LKK/+
ChsyEvFhgiPFl9ScqCuHYgj1lm9s6Y5Qx9uxODur0XliUXlo6cMT9r33YTdTX9JE
lUBanI6APExJp1oL1CCTWvK52Nk8F9OUxw5Wc3OBHmM4ffGD1vTGdLmTVA6Q3A3/
/nK7eu4vubm27382B1c8PcHRxCaXO0cpc+KY7Qw9/Bfj4jbkgwF8MnbaN1r31AtW
rR6IjziSShrtpPq89b5Tj7ZmAQC35M56X0ZXKX3Vq7VoHFxzDNmrw3fi5GrVdtUZ
jpaFDf6R0dhMEEipr4vaKFJKMVBkmTVH9IgUGOc5bIePvPIZnNbTZiGIRZ/yk9Yk
77o3xaOh4dLpRMqr3PM/buHcFC+xvbMsffNQ7ajXMBOmqcVsd5LNiYVwrZ6gFir3
hlem9N8oXD0Vf+kbB7qmNNgWkhWjVo7TjG0YtFOJHf5po6u+Xrt9SDzCVNnUbSAf
aA4y+j88gMkVi/uops7tRUpsYohaF0KyVED9RDMLzF+4wPJW54kYJhOD9MqIaqGJ
UaJwRaVgmEoj58lAzLiwNzYicesku+dkqHkEUkqsbQKXqhx8JDilK3YzwpikpXY7
iNZo7EnYuyCyYtSoiuarWanYIpODsyexU623Q6oGEzsPSTfiLZwa2XRNWqum6fop
IT71y+xgZ1h2l5PUay82n1zspStN4KHuHxm25K0vZcvT+oEW2j16OKKN4aiqYNbu
J5UT3ZljKsjY9nPzxE6b1ksvsacHSk31CXwYT34YrAMPWFQoWIqin5nBG3ha8SJ3
1R9V1SLwHeRpe2u2I265dCDFfGTjqa02aSTu6RmYwINgRcVj3ApAQbR8cFxM/ooX
gJiBEgG92cv3U7RkfNVknVB2zAtzUg7WMW+oMAJDu5ohx6Z74MKQBCDTC6lBUuTO
qrbT98VpfK6chMJfgIdawJ0fU5rJJSxVVQVOv61oUY6Ds3Rtod36XcN2GrEHnhcI
wJOIsPB+ZptE74hEo3oiTl9H2v6NK26soQHG9/kVOMFl60KGqHVMdDL3xAyDWZDP
vAvtMOAKvpOGZ7KQyzebMIfYY/v1Cxallc0XrFt/bpbqMxlJCx3AkSYnK4E/F7nz
DDF9OydzjIRrthEGJPHDGnBvEIKYNOYCFglKiXWxcYL3KnqOtjKL98A6HFSPEhTc
0PymGn/wBkSAsKUc6IvdEbrstlC+MaezqD9JAwHVoxDWHzg5g5B9O9DUnwPrpsUV
szWSXQ9+/qFxoXC18zpjHlvLj6CnnIeakifNMMeq6qR44SDNzEf0rrYcrpB/MOBz
OdhsYUyDzqmZBBqJwrYrxYnS6dKms+ZzKtOcJkQd9KMwvE5l4QV/c0o3jcTjW6aV
WxwiXmjTk7KPDrAsQJAZIn3RhuV9QKU2ykXEaqh0TRLX9qEVUr3F0RJlk8S0Qr1l
tklYF44ZbbS2qvpa8Hw3lA/qxtTiDUpUd966A1Tsgs1ld8ysEWrwPRtx6WWYAj4r
TBgmTS0tIP5eRr9CTP7myT40PDNJxEfmIw9ZjzrGNSBdgt2wpUzbps8K6seUXmHG
h3kldPRkMKKVecmiQ8oME8lMOB8MZwO4bALBM4+pHv/hBEpgkbHadTgKh7TsnmKE
dupqdm5Y5BqDo1ckgxen8KPdND2i6Z4EGso7ZtFNQqeXpENdN3aBguEBpMIOHn1U
uOLocuXg9r6JxmItuGmwvNUluXHKSFw2I4T6eHyQ12WcBvpY0sNlVy6rLxQazPGi
qV4Y30FG85Xye8w6gZwbJ3JGRQZ4R3JwqSHMXft2UxjsDJwhZv8+F5P6/upsPd30
HIiMy5FPsqq6CT2tQtb2ErGXSzf0Zi6IuC0g+bRmqlwGR7ah0igSGDBD/4iYdYwY
cbPAjxYpmPP5JeLQidQAbab4UrDvCSmRidoSMQus1vx3nZsGopQYqmgE4a/ioFHh
N0DWocY4E77NpFUDjpvl8iwZCwEkwHlMe4wp+JbiDCTQEp+IWCFgNrj4HXXi3bOi
13b/XvVNQSCwm9tKWdI1GKEriarfSNEcMLOjOZfzU80DggkkuaYq7VXEl2r6dkfY
t2QcKJuq8vVbqK7ZYCtTD1XzA2Lqwc88lT0HJcAArBukB4l+yZvSg1rEGg9Q8v8i
C7Kb2ZKfisHnKK1vxrG7HOYgq0AC6unVMUphVtNSaN7eZfwfzWKcGo+UBam38sed
vSfulRI0CLvA95YfCf+Yhl5Wk8NNP7bnngDnvZgFi95ai6aJqL5sDMgn3HmAHgMY
gi/0D2e9rQNafPi2He/TvZeX4hyx1N911s0ixjF3CM/k6E7nY175ykvkZo5s2L3x
ktp+swVsN8Hxfe6uxzTfgdPP3HSPiTGKwHBbqSsIWLTYv+4FYQzNyS4jpYjbMU0s
uQrWfn4cYHuC8Ef1Cg3Un5p3aHC/ZNwaI4gy0iTkx6GJK+UJzr9RLZcexl/arfQ1
5kt8+pOlIBV+4gAK0FYdmr1+mX7ZPagE1ZpBZXWS8q1pd+Au1fT2v+xqdQ7IjE06
s59VCHC4T/Bf67VqQCmMVOvQVof/FLXB1xv9ZOlNVngZ9yQyN7Z4iVnFiwG6u2Nu
KF0+f5KUX5q7cjWs45CmpSBZRqxEU1iNPc+k8piyp1Da86Zz4X9u/p3V4uQHvTUe
awfimd+/6TTVYo5S2hNxRHgnS62joBUYaXAM1zIVa5YZFPgPNBeWGY97tTX6f/6J
aRFnbYXeOb0cZhPB4JwsAb7xUqJBvZQWVmGbXkdgLtOb8TZNakrEZcc2+Ur9twjx
R1IFr1MyP2qE5CZ2DvgbbvEnG82aC4k2X5UPRjMrNSxl2jOBYeBrbhnnA35LbGz2
cO6S1ONfkqq/UANb0+BWDy50hxebKpbdRakoFIB0lYZh3QLAXTYymx37+OCxb1yf
g7W+X1IXNs2aHPaNcTWvnh0jUXDILLpVINntilIXQ8INpZz3Bs1htMxl7pE9SS2J
BiUXc1vhtzB1zZtxi056taXHkxUx9s/UVpxTTcOfDsaxj9ldk6Hd99gW8JLp2KFZ
fuku9bAlx3n2E4O8K8vcw3dYrCCdlQP8Sp8QRm+lMY1j6GYpRvLz/z4iSw6sUTz0
Undkk1JiP8p6RIsJH9q9e1MfIvFoNC/KT+MgHlHxxZUMyU8lZfH80LQPzUZyAUWS
xC0WvpfQ9P5oU2GobF71C4aK27AQ0SLN5eivM9vKJp/2JC1aDKxgWH1SNzsMit98
O6eE9s+qf0NVP+wHPg+JjMBMdcxH2BsWZcfgc0WPc5OU3VIcVWeddsEaviHpZiOE
V2MPEy9cmjT8cFxR9M5LZSidr6XKDcV/5nfkKNZNkFjnf5/IrUWax4AXfJgDZKRh
cKh8rtnLizbLhbTLDy/jU5zPrmUD/AGHJ9kkm1ms7FUqPb9S7UNZ+E22m3zXZHc8
z7o5Cva8qSB8u6f3tt9Dksp+k6WJUzc9E50TvBoG/7azPnePvXWC314PtY62jULQ
ITZjbS3efWiS0CnD5qXZXqhOZ4GDnHZKvhY21Yql4aZJhTFf/ezkYXEBNkMbsMoN
uKXuIoK1FFWhxhfptpZBzTTYpoUUofAaMxopLU4k0J4uh7B39L5RlpDkUUduxAOy
ywX4QVYpdx+GOv4CYRXiCsI+yhBTjES2+MNrd+BdYbVaVDuPgW/3JyHJn8Q0FO7H
R8w2JOUwGdeM5cYX6aD5VtiMFQPbO0ve4om+ge7U5N7BCujGOkpy9NjgdMdPcixO
KNNbDqenym+ldxiVnTb+oBcJeQcIy+OQwJ0kV9I2OmsVvyuB+A2nfUY2an17PfPM
z+XBTr9I4yejbZqF05JD+oDVczsS78dsZu2QdENp9cnz07KLhYk+j7dobh0TVjuA
Akwyk0VXbHo2BNiunMaG4a14WsUe9A1DCyR1A5jZRxc0qlJk7ebyogfhOmwLnNuH
vPvY1nOEwSlmkI2wWzg0KP+wA86gTnR5GQMBEt2PzUidd0OZBmj2DIWxsYnoyqTH
Mg9rlbKTNgGQgaEo6IAqTrkyx/y4c7sHEWJuH0Xed6RLGCyhzgesPgvJ84n5VFPi
7S1qiSeUWEmOAKg/6KpzYyNHkuU/v/BXArHVfvySGt50YbS43K5m8+FFc+FOwdiN
wmqa6vxHwI+unO4tHI3Jn6l0ejdTBlYQWpxTGw5odHvj9dbT+MsO+it98+r3uTEL
tO64cRdW8+DHsw7XG0kwLChbpYx2HSYoS4qigWo6aMQ0fklM9sktwfDH8xEeCwsT
/L/W0eNQEKJFIfxxbwodRxuex2P5xsFt6dRC38rRry4ULbgEbM9NKE+yBxiMeqKZ
MxSEK/RGfMqBQKF1Nx/Z/p3wQf1J6vDiWwC3modilNqwI5VVrn2pAk9r1+22hVNL
tNQpVnmdD2viq/wKKivk7PU6+cxu78fs26RYUR4OLeomd5O4a8qlooJSVdGUg+De
2VwteDyTceoc8AZJZ1sVyt84mjc0m6PwBlHgmu8orJdaEVaP63KyU07imm8E4DYT
wTV+6RKI8na++CBIWi3ybSozGay7EJrOoc/HOg0QFuXlST/YJBgMcP0PSStITngN
Yi3Ed/i7W5guwRKSKi0KUP7TADAU/fkT5gegpZHQdwZYPSjgqBgTWSA6uKQW82YX
ne6obTQgKhSlcRDqT3acur8Hi2n8Gftc2AkXOGmzY0T+D9VdgYYAUa2ruEAf3uZe
mnjQxHIZ/noPCKkjKQhPLm6+TLMX86+oRp+mPmh8gMDBnjau13SOi6HC2dnL9BZD
uv9msGfvHCLDM6YSEBFQI9c3p5dA+5066FRCE2po9uJhFb77zsuu1UHmpZL78RtA
UUwvp0+h8Q2warT65SKiiE9ramlHIwJgjZC7M1MMUG5eHcXcf3+hsDLzTAVA5Z+E
lOioAyYrzJvm9e1EYM7ViDuNn2L7DAJGoOG3K/Ai6W14MTyZpQOqOadsmktCvj1C
ETIEVA20gv35kgrqXxreqB6j9XRpwQBn7GP/W/DjEWDBwYzv8n7qK6v/hm7ZVRF4
7uAQ3v39d7aLgpKc+Lkeayx6Dp2nfG9j5RaVyjuxGALiE5pz4t8Hwxo2GKYdU9MO
Gtpn/5LDfM+aT1TIrKP0IvFPhxglju+yS5XUdjY8wjuP6jdR4/zyyKmPPP3XXWSW
hGzXK+9hXP0Z4VTdJxFhWuPKTIpJqJ4cODSCJJKmHtAYfFt+5jTznH8hPdsl9rTO
J0ZlR4Qsdsgpk3lQJ+HNuLRj2Xx+R++QNUm7NmYfEAD/O4yhD+VM9vfy8ZL194md
Wf1SWBEGGA5b5nlHM0ABhxkkCOYfl7/dq9ljODJGRMewdDjnAR/KrTSeVZe1r/bV
yxm0jUv3qTpEpL0PQOGYu+8qKzUVz9FnkIVKte08TOIl/pR6NNU1C7/gFsH5umq3
F3HN9D+SIHRH62+3qYBh0xMJTWnGUzzo3k6LnssrpRK7lVeYRwXeWNdBr7ldpF/y
LTdm4f/dOTOc91IVQwP2nGRs/hKPZIaLirjxjBqlOQgJRo66deQmMizi+ywQ3ehX
GthEs6+orSkf/Ql+bAZCTZiRMBp5j/m08uwSVUbplj1f5F5wWIdveZnWrCLyfJJO
YlUVmRbsvN8yAHn8ryV6KXwDCpKvoJmeuwlz2trAlXGUvgR//trGRFTGC4DU1QCb
wkf7w/KGxX5nphBMpZa6b7qURNC59+lNjonxe1KXbM5yxD+VqssElM1KVrrYTFj1
g+ommEn0Ru1owyCCHD3dPnOVOq5dYdmhlIZN+/WnLM6yhmSglEEvHfuz5/EGookk
tWnImbsx88RVlLYMg0+UzMqcDK1ddt8SOd28IMCDd1tYtegI/XBbGBjC4SW2kg9+
8lWl6DpzwK44IcwKrJnnPBeED/XZ82qE+jFVqtABpnLFaUUZZR7M4DjEC3fspnpj
B5UVIhazi/pJzlha9/ZMQ0niNFaOCFdqghqaS3XF8aFQZjZAqGWlC1KWLyQ9q/I9
KeuvJrqGNGVu3sEyrGSk1XLUyqRA+f6lVWOcaP/eIGCMH0SPcGoEXn+2PuJEq+ti
bqTQSo68gBq7y8mv7b5yeVZghYUy7pE1WIR9rC/OwnjS25fzJ0AnGfhbseO7MKfz
s0PMLOSwXKPNMvTdFMFxldIGqgUmuSiqG6aoHPVzYL4kJpdfiqxfKxBzAu7y9HN3
mY1Lpdx6FGQUxIqOplkleIM0CiwVl2nKzmoR4HcXxGXh2Qm1P9z1Hx6c5clrVA/r
mj0B9O8heIQTdmWm+/lDMV0QIroTHFWJYYyhGokRk7OnvsZ065IsUz0VRM9MPS4r
tID/LgSXzEzNjnBqvQ0d3d6tLxtnVZQTUYL+P7Q71A39zQ5lTC3kz00u61o1HRVq
8ADzMu5PtlqT3C/p1kj8VTa9iL9dxn/+UUqFYC5L157fzCPI/hx0u/tjytG/Fxcf
M+ABBQb5V2iFtlmVUXnfO6hj0+RMRNdBAUvyjh5jT0DtD/cTNDjr8XvvwooitU6Z
dGk3ZBXd6ibnkbCKID+jpaGdFXB4D3rsQqgyf7oDQqcEOAPAEi3YjZahO4ubnBZR
7GJh8FPaL6xwJbSmHmOU9PQT2l+fw+lJzFQvfo3hPpNUBp4uo93/BOBqt9P/yDZn
zaHaBRL/nC6Xx+z/QXZyslKsgTeyD3qKOcPB2HPqxgjP1bEjH0OloDhNz2QULXwc
sHRSb4noGhjjHnr0rsUpDxJ4FwmLgA/Eu7l3WJmUX3rm1Dhtf4OZGJU7AygHBDyL
BqqW6+S7VeCGhURCYG0QZUhJH5Hnctr/ich0nUXUoELtKFJjycaolFK47XRfKPbe
Ok3EyYgPX5qRQZowZ3xOdxAEIq3WRQlxm+7y/56BARDdnyzN7eqbmBbupQw/PVyh
FmsBNCikJaptTKZ7Jcdf85ToIIkkG6yx+HIN15OKj2n+AHWaXdkLOgzk8Rppd22c
3s/xosMPW8WjBCJMf7VGvNVLDi5pWJxvzSNgXgw7Wm/GD1IO0bhD9gMB37U2CXFv
9UWENSiBGkbn28EoBVVerV1nV4trZGnJ3AdczUsllSflBJrBHLmv74PH0edY8pwX
3hstV5lDXZKpvWvI5WYDiFOc18Aqp7PLFk3d6C8ox4LVRFjyOx1wUXNA++1jKtku
7gup3R2xBBEB8gCBkM0ZlyeQ2KbCTdjUsXTWrE3cWbhy1uc8By0e6IOCjNW6cT1U
yNgK4aEpfDuYCAf9ZZbJXe0eaTPkXYgR4QB96C6PcA/+1PXpdwEKaCK8PH6tDUt7
YgKbhVeR0sG9hpXUUywDfBn+3j3OBpBLYIyiRA6npQC8OsQ5LUTsNN6uaDWa40ZZ
q8qPybet2US2NgiM3ia3kPq14MXLE69yIRLym8EyqNNu6IZne51bK6moa118+6WW
puRlofIZZ3qXDJmobwCOcFqLKJwdN3uyuKTNGMH+zAlOtYel1pV5apU+ual1ua0H
RcFQF3y53vjz9LXjQ5pfpCPWJoo3J91cGcYoYjJQJ5UTzSdTTX+W+odGawEfHUuJ
YT73p7j8u06A4QwhxwZzc3JZkU3lcMJ/Fjubuz4vWJPKG0yhxVDUlV8ulOom4jqH
bpnk+eH7vYxX7PzoynZgawHmXa21SpR+RsC54TZ4qK7XuM1TU6NUoC0fnBwYX7mw
MFQwo6Wh2YKfCEqtJCv7hD6dDi3W4K/yzDh2RpqF6AkO6NWvzJrj4IliG277N9z6
Fkkh9ILBke97Py2ElIqsEHNZycjpZ4UcoHEEgEnASRRKn7aX81ORfK13HKat62D9
m1c7FZAbqQFHIkSObefPUuEmYGAN82in0wrHna4SYiEI01CLKNxQLeWTT9iedrMY
fR3Yr+RJzc0L0MaBzE92bwTpKSFqiIykDjda/RvBr/FbxT1/IM2b3FdR1XX2KT1E
zgjNVRyUp+U9wK9AVVQ4NQIkXsd1GFdrEUG5hwyLJ3+k3CE3ps6tuSdB0ijbRl/n
BZSdpMuoLJMeKcfVKWRErZ4R/L1A/oBufTSbWw72IB4VCMtnUPnWwkM+Riu/xulv
syba26O6Xj3hxvWboZJ8kIXqUjViazPSJRmg7h+5gSh2KR9/mqU1qxqhjb3TQoup
JKrE0OHzQw3SB4uR7I0HTWQ8f540nKU/1sFUaNUSAf+OoHYd+cvRMY8sxgX0GmZ7
DqQPImNfO6+Z8V9PWQlolWQawF5eCCXJ2Ieje1opAO3LL4/4RChYpjIHmCxBLEz7
PhkVwuEH69T817ow7pirKpMozPLOo25Yl0yz27AVNQH4pnxsQOKkIs5ox70O+ELm
Tuket7msTRN6jjl0tBufO/qqBCNACsFfBNC0gwn2mkLD2WLuUVqYCcVM2JuBfusO
98dd+pFaqK7aYtRfL8VpgHOQ5x55lKjqU1MafUIoPXmMgGhro9dCh+H5hTof8lVl
Ig4onlx3lDPXardo9SOp89NCm3DkKvbtxuVo0BbbM+UhLuHdi0lmQL40iWvHVjh+
sYbFNilMm7DeZsp/62JfBeDps7lzVe/GGcYS+sW/kA7KbedxqevckPW3n9q8sut3
cmuHmC7hrIB7ZcF9oCTVQ30JpM3tHN/4E9yljBhn4mtRv22+a5PKDOLmTvd6CBcJ
2wGdvX883Qlql3xam79xwJIQi5Hp5zXwFC4vCsZcPAVaRohqRpm3Lg2+vUggumDw
mTJh5XMSMc04EPE+CObdJmzlqDSc8/0V3PJbREw5SBIipSPXd7XgeCjRNdMTeejn
7LYnlWqHCYklqXhFD6qxj8ci8fefztEvz0kQuS9LqxFLdeY/Pzs7h7DTzA7fkJ/u
71sxo/TeSQ2JE5kiPUdJvpQOx/D5VLki2VgiXGUELxNFYz1+X8d7B78naun9odUk
hXkd3HpW/zC3msEgFMo6pDRPYDdC5l7oHPEIFqj1KjfXhCwQ9s2iJXsolg2TaTxd
DocvHgXqMntp/jFthtS905RzoKOiYxas1kcPqHGUaH/zKhp26i71Z+9o2/El7lJt
pBk6T9QJrJfSw5vsLQkEvSatiFeJoOzMFsHCh2kMEA5wJApgEmeWwWDiMrmmtV6O
RvCojNCv4JrbE1pTztygPVFtO1GSBP7Sgfa6uOgHfNiiCN0qy0q4FTwT4ibpQsDQ
lomRpzWEAqn8Rpt5Chpp96coVCP1uc8jQvXnZoAaiYfQHs7fMSxB/sg+PAwB3uJz
3yNfxbqGN2IBh5ziKNYv/2u3hWCFzPrj+seOOXil2Ebi9rmPg+vpYfOsefXpZrit
xZ+S+uOu0+j+BcPsIXARWPs8PeryNNZudd6ChWAq+IUzpAyOFcXU2aJK+/AngWi5
Qye6gLVAcKIJiuXtaD2sMn1wCoMOw8dbUA69QQjUYmcDUyyfXpzloMzFoa5xXFaV
kvHmJ8mY/Q24TFa/Gn3XWU4qmHbnV+Mw0oktB6npdQaRjs754uZiYpBtvN+CYopI
4G95FUT25s6KCWGp5Fv+RNkb13t2gZvBV1qiupoyO3di1spJx8ec4JV6AzqfBItM
r6JFBAEDcAVT1TKqqbAHi65jufP+pDbCL/DZUDqUHexVdspemYFe7Gt22DFyCqXA
qWh1yn2sg17jTVhycA/buI99emlBcvqWjj57ya7Ttrm/DReuHEejOvJqDOieNwUz
ybDydWSX7s5LVoDjyEKW+1iiGU7pCzo2582G0pDcVGucwvfqy3xoeMRTm1YAo6If
1+rZswQkwtI1VH/CvXtSpcRbcgaKg91jds6I5xd7d1rkEKW7mZmUoa3VnL/Qx9ai
IpjjeIK7trAzh3ZmUmu/YSWi8cO9mFXmgIi5VsaxMiLgCmBmmhG5vJxlFL26HhDY
5T2DVAQNMAslv2ewtydrbqjJs0ntS3APs+SqDleWtGT2obQE5fKtQDSxKMf6Ygbi
obwC8LnRViWuQ4gDZu4B6NpmEUE+V5SZKM0xXtTKZnukBK/qQc/M1uak4+0NcU4d
wK6kj3yhXsUd4C/B7VxXTHjDh9/VDqZrbLmu2ziZB7NSVgW/5VRg1RvG+lUT15n3
`protect END_PROTECTED
