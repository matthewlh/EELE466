`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
hRP+YjjVwaDW0gq//PJYDssfpeyBzsSAfxstgg1V7fUn9YSXokgp/W6w/i/UQ7wV
uiKdr2RhOZDvPst7UcMBMwdJf1MFbKc9LpuCgmmSjuZwwywPizJJRsxiXUe2JivW
ZlRWFMAnRAAcQj4o1xYspx3IBsidpSt/gtVeSE5QCrm6UILOGuXcq3/Rhp8nbkKS
589A2AHgA8mEyJI0ytHKh4gJsPNqsArNi6f70w23I+NuRef7VPYkbZ/Klf8RK+Kw
prBQ3GC33JlBzrdDgNci9U818zZfM13e83+UXJDxNfa+VKGmKN4MtbYv9/rBjwSm
ipGY9C+NZtu46Cfhtwjy0QAt2+2twCNOWggwTOQXZPL3MZHbI8cNemNUqqpJqbCz
YM0AvuGR2Gzel681XFw2m1BxpSuEK9SHD5u7VyL94TaNKZU/eRiombwiJUMMIpJr
khZo/lJwSn5tF55PqXo7zDbipedKYPsffRZRgN1b4N3HuPgW5kDC/POrUcxPAufz
bo6u4HnDIroUcQykhH8rpBV/DtZQgfqb6owN+jvjkpwx9Qh/MAAr01PUsJsjnZmC
yX5yunq5thDSHgwoYifecpVCoj8KkyBKZdRNI9NQpXWBcYSojCATh2zRWJhOVUMF
8t8pieuJ0mHSdwS4Qvc+beHqLs0pXZjCyhYFSbIXI4Q1cCpKrA/WhqEYXSesW64x
ghwAK6QfX+83k7Dk+otsiJFEAPhwRrmvBici2ZD4ueExZL9nxZGqJ/sJ71zQDL76
J1Q12rrtE2lVp25zhfgiEfp9bHFoVQiLj0N9CWbPOhg2h4dSmDZtvlqdq3ITFzKn
HU+VMduS93V7wGzxIoRpOkfkTeSxLxTQntT3eopcqe6/cAHGvVJ2IQbEwyU+Ae23
vFYg0Yxjc3bgpPmmsUhUbaovQzk5pydO8RcMt0//A03jFpmIaNlVpKK+0qfmRjKe
byNt9vi1An89CkxJLEOHEZlqIe5t0bB6pHQZOWIlON9rW2f/bD85+eYtTppbfmyl
Dj/7b9lPLP252FERPMmlnq/X6Cmpt9qL+r/B1+griJ/uoiuDZSfHw+4S0+ya74F5
2dXzNf6donUyuuM5Bb5jUOPykZ1tFHjTSP1RISULKypYhDGyxTLTVvIm/r2xrX7N
axdlU1uM81Z5Y321oRp3ochU23fF9aA6c1qE8XIzqqaA9VLXK+tTXZnqy5uK0EtB
EeM4T9ymZDGtZwKNs35nvvnsVO2SIt3+r4IplpanPLarEGXmMduGw7mAYEOKNLNB
mk5t7XzXJO5xdBOtP8zm2BFW7ck09OfooFFPT9RBGP0cVVCs52311Wh0dzvKxq1v
HMDRl/LoEyISI9cum3Bp9ZO/mEJWsLfO2vcQNSUkW4tiqI7B6n56eMqPge80u/uS
hhSixnyy9TdMHWAj//fy52/DLSjs+jCik/rl3bxJ1vaRkMoVkiHGGqG3gFxnom6r
TrOcHxds1p1Ya35nqDZT20pJc4hreC8niIvWph3jaCs=
`protect END_PROTECTED
