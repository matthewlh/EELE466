----------------------------------------------------------------------------------
--
-- Author(s):		David Keltgen
--					Matthew Handley
--
-- File:			lookup.vhd
--
-- Create Date:      03/17/2015
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.numeric_std.ALL;

entity lookup is 
	port(
		CLK				: in  STD_LOGIC;
		ADDRESS			: in  STD_LOGIC_VECTOR(15 downto 0);
		RESULT			: out STD_LOGIC_VECTOR(15 downto 0)
	);
	  
end entity;

architecture lookup_arch of lookup is

	begin
		--------------------------
		---- Signal Assigment ----
		--------------------------
		with ADDRESS select RESULT <=
			x"0000" when x"0000",
			x"FFFF" when x"0001",
			x"4000" when x"0002",
			x"1C72" when x"0003",
			x"1000" when x"0004",
			x"0A3D" when x"0005",
			x"071C" when x"0006",
			x"0539" when x"0007",
			x"0400" when x"0008",
			x"0329" when x"0009",
			x"028F" when x"000A",
			x"021E" when x"000B",
			x"01C7" when x"000C",
			x"0184" when x"000D",
			x"014E" when x"000E",
			x"0123" when x"000F",
			x"0100" when x"0010",
			x"00E3" when x"0011",
			x"00CA" when x"0012",
			x"00B6" when x"0013",
			x"00A4" when x"0014",
			x"0095" when x"0015",
			x"0087" when x"0016",
			x"007C" when x"0017",
			x"0072" when x"0018",
			x"0069" when x"0019",
			x"0061" when x"001A",
			x"005A" when x"001B",
			x"0054" when x"001C",
			x"004E" when x"001D",
			x"0049" when x"001E",
			x"0044" when x"001F",
			x"0040" when x"0020",
			x"003C" when x"0021",
			x"0039" when x"0022",
			x"0035" when x"0023",
			x"0033" when x"0024",
			x"0030" when x"0025",
			x"002D" when x"0026",
			x"002B" when x"0027",
			x"0029" when x"0028",
			x"0027" when x"0029",
			x"0025" when x"002A",
			x"0023" when x"002B",
			x"0022" when x"002C",
			x"0020" when x"002D",
			x"001F" when x"002E",
			x"001E" when x"002F",
			x"001C" when x"0030",
			x"001B" when x"0031",
			x"001A" when x"0032",
			x"0019" when x"0033",
			x"0018" when x"0034",
			x"0017" when x"0035",
			x"0016" when x"0036",
			x"0016" when x"0037",
			x"0015" when x"0038",
			x"0014" when x"0039",
			x"0013" when x"003A",
			x"0013" when x"003B",
			x"0012" when x"003C",
			x"0012" when x"003D",
			x"0011" when x"003E",
			x"0011" when x"003F",
			x"0010" when x"0040",
			x"0010" when x"0041",
			x"000F" when x"0042",
			x"000F" when x"0043",
			x"000E" when x"0044",
			x"000E" when x"0045",
			x"000D" when x"0046",
			x"000D" when x"0047",
			x"000D" when x"0048",
			x"000C" when x"0049",
			x"000C" when x"004A",
			x"000C" when x"004B",
			x"000B" when x"004C",
			x"000B" when x"004D",
			x"000B" when x"004E",
			x"000B" when x"004F",
			x"000A" when x"0050",
			x"000A" when x"0051",
			x"000A" when x"0052",
			x"000A" when x"0053",
			x"0009" when x"0054",
			x"0009" when x"0055",
			x"0009" when x"0056",
			x"0009" when x"0057",
			x"0008" when x"0058",
			x"0008" when x"0059",
			x"0008" when x"005A",
			x"0008" when x"005B",
			x"0008" when x"005C",
			x"0008" when x"005D",
			x"0007" when x"005E",
			x"0007" when x"005F",
			x"0007" when x"0060",
			x"0007" when x"0061",
			x"0007" when x"0062",
			x"0007" when x"0063",
			x"0007" when x"0064",
			x"0006" when x"0065",
			x"0006" when x"0066",
			x"0006" when x"0067",
			x"0006" when x"0068",
			x"0006" when x"0069",
			x"0006" when x"006A",
			x"0006" when x"006B",
			x"0006" when x"006C",
			x"0006" when x"006D",
			x"0005" when x"006E",
			x"0005" when x"006F",
			x"0005" when x"0070",
			x"0005" when x"0071",
			x"0005" when x"0072",
			x"0005" when x"0073",
			x"0005" when x"0074",
			x"0005" when x"0075",
			x"0005" when x"0076",
			x"0005" when x"0077",
			x"0005" when x"0078",
			x"0004" when x"0079",
			x"0004" when x"007A",
			x"0004" when x"007B",
			x"0004" when x"007C",
			x"0004" when x"007D",
			x"0004" when x"007E",
			x"0004" when x"007F",
			x"0004" when x"0080",
			x"0004" when x"0081",
			x"0004" when x"0082",
			x"0004" when x"0083",
			x"0004" when x"0084",
			x"0004" when x"0085",
			x"0004" when x"0086",
			x"0004" when x"0087",
			x"0004" when x"0088",
			x"0003" when x"0089",
			x"0003" when x"008A",
			x"0003" when x"008B",
			x"0003" when x"008C",
			x"0003" when x"008D",
			x"0003" when x"008E",
			x"0003" when x"008F",
			x"0003" when x"0090",
			x"0003" when x"0091",
			x"0003" when x"0092",
			x"0003" when x"0093",
			x"0003" when x"0094",
			x"0003" when x"0095",
			x"0003" when x"0096",
			x"0003" when x"0097",
			x"0003" when x"0098",
			x"0003" when x"0099",
			x"0003" when x"009A",
			x"0003" when x"009B",
			x"0003" when x"009C",
			x"0003" when x"009D",
			x"0003" when x"009E",
			x"0003" when x"009F",
			x"0003" when x"00A0",
			x"0003" when x"00A1",
			x"0002" when x"00A2",
			x"0002" when x"00A3",
			x"0002" when x"00A4",
			x"0002" when x"00A5",
			x"0002" when x"00A6",
			x"0002" when x"00A7",
			x"0002" when x"00A8",
			x"0002" when x"00A9",
			x"0002" when x"00AA",
			x"0002" when x"00AB",
			x"0002" when x"00AC",
			x"0002" when x"00AD",
			x"0002" when x"00AE",
			x"0002" when x"00AF",
			x"0002" when x"00B0",
			x"0002" when x"00B1",
			x"0002" when x"00B2",
			x"0002" when x"00B3",
			x"0002" when x"00B4",
			x"0002" when x"00B5",
			x"0002" when x"00B6",
			x"0002" when x"00B7",
			x"0002" when x"00B8",
			x"0002" when x"00B9",
			x"0002" when x"00BA",
			x"0002" when x"00BB",
			x"0002" when x"00BC",
			x"0002" when x"00BD",
			x"0002" when x"00BE",
			x"0002" when x"00BF",
			x"0002" when x"00C0",
			x"0002" when x"00C1",
			x"0002" when x"00C2",
			x"0002" when x"00C3",
			x"0002" when x"00C4",
			x"0002" when x"00C5",
			x"0002" when x"00C6",
			x"0002" when x"00C7",
			x"0002" when x"00C8",
			x"0002" when x"00C9",
			x"0002" when x"00CA",
			x"0002" when x"00CB",
			x"0002" when x"00CC",
			x"0002" when x"00CD",
			x"0002" when x"00CE",
			x"0002" when x"00CF",
			x"0002" when x"00D0",
			x"0002" when x"00D1",
			x"0001" when x"00D2",
			x"0001" when x"00D3",
			x"0001" when x"00D4",
			x"0001" when x"00D5",
			x"0001" when x"00D6",
			x"0001" when x"00D7",
			x"0001" when x"00D8",
			x"0001" when x"00D9",
			x"0001" when x"00DA",
			x"0001" when x"00DB",
			x"0001" when x"00DC",
			x"0001" when x"00DD",
			x"0001" when x"00DE",
			x"0001" when x"00DF",
			x"0001" when x"00E0",
			x"0001" when x"00E1",
			x"0001" when x"00E2",
			x"0001" when x"00E3",
			x"0001" when x"00E4",
			x"0001" when x"00E5",
			x"0001" when x"00E6",
			x"0001" when x"00E7",
			x"0001" when x"00E8",
			x"0001" when x"00E9",
			x"0001" when x"00EA",
			x"0001" when x"00EB",
			x"0001" when x"00EC",
			x"0001" when x"00ED",
			x"0001" when x"00EE",
			x"0001" when x"00EF",
			x"0001" when x"00F0",
			x"0001" when x"00F1",
			x"0001" when x"00F2",
			x"0001" when x"00F3",
			x"0001" when x"00F4",
			x"0001" when x"00F5",
			x"0001" when x"00F6",
			x"0001" when x"00F7",
			x"0001" when x"00F8",
			x"0001" when x"00F9",
			x"0001" when x"00FA",
			x"0001" when x"00FB",
			x"0001" when x"00FC",
			x"0001" when x"00FD",
			x"0001" when x"00FE",
			x"0001" when x"00FF",
			x"0001" when x"0100",
			x"0001" when x"0101",
			x"0001" when x"0102",
			x"0001" when x"0103",
			x"0001" when x"0104",
			x"0001" when x"0105",
			x"0001" when x"0106",
			x"0001" when x"0107",
			x"0001" when x"0108",
			x"0001" when x"0109",
			x"0001" when x"010A",
			x"0001" when x"010B",
			x"0001" when x"010C",
			x"0001" when x"010D",
			x"0001" when x"010E",
			x"0001" when x"010F",
			x"0001" when x"0110",
			x"0001" when x"0111",
			x"0001" when x"0112",
			x"0001" when x"0113",
			x"0001" when x"0114",
			x"0001" when x"0115",
			x"0001" when x"0116",
			x"0001" when x"0117",
			x"0001" when x"0118",
			x"0001" when x"0119",
			x"0001" when x"011A",
			x"0001" when x"011B",
			x"0001" when x"011C",
			x"0001" when x"011D",
			x"0001" when x"011E",
			x"0001" when x"011F",
			x"0001" when x"0120",
			x"0001" when x"0121",
			x"0001" when x"0122",
			x"0001" when x"0123",
			x"0001" when x"0124",
			x"0001" when x"0125",
			x"0001" when x"0126",
			x"0001" when x"0127",
			x"0001" when x"0128",
			x"0001" when x"0129",
			x"0001" when x"012A",
			x"0001" when x"012B",
			x"0001" when x"012C",
			x"0001" when x"012D",
			x"0001" when x"012E",
			x"0001" when x"012F",
			x"0001" when x"0130",
			x"0001" when x"0131",
			x"0001" when x"0132",
			x"0001" when x"0133",
			x"0001" when x"0134",
			x"0001" when x"0135",
			x"0001" when x"0136",
			x"0001" when x"0137",
			x"0001" when x"0138",
			x"0001" when x"0139",
			x"0001" when x"013A",
			x"0001" when x"013B",
			x"0001" when x"013C",
			x"0001" when x"013D",
			x"0001" when x"013E",
			x"0001" when x"013F",
			x"0001" when x"0140",
			x"0001" when x"0141",
			x"0001" when x"0142",
			x"0001" when x"0143",
			x"0001" when x"0144",
			x"0001" when x"0145",
			x"0001" when x"0146",
			x"0001" when x"0147",
			x"0001" when x"0148",
			x"0001" when x"0149",
			x"0001" when x"014A",
			x"0001" when x"014B",
			x"0001" when x"014C",
			x"0001" when x"014D",
			x"0001" when x"014E",
			x"0001" when x"014F",
			x"0001" when x"0150",
			x"0001" when x"0151",
			x"0001" when x"0152",
			x"0001" when x"0153",
			x"0001" when x"0154",
			x"0001" when x"0155",
			x"0001" when x"0156",
			x"0001" when x"0157",
			x"0001" when x"0158",
			x"0001" when x"0159",
			x"0001" when x"015A",
			x"0001" when x"015B",
			x"0001" when x"015C",
			x"0001" when x"015D",
			x"0001" when x"015E",
			x"0001" when x"015F",
			x"0001" when x"0160",
			x"0001" when x"0161",
			x"0001" when x"0162",
			x"0001" when x"0163",
			x"0001" when x"0164",
			x"0001" when x"0165",
			x"0001" when x"0166",
			x"0001" when x"0167",
			x"0001" when x"0168",
			x"0001" when x"0169",
			x"0001" when x"016A",
			x"0000" when x"016B",
			x"0000" when x"016C",
			x"0000" when x"016D",
			x"0000" when x"016E",
			x"0000" when x"016F",
			x"0000" when x"0170",
			x"0000" when x"0171",
			x"0000" when x"0172",
			x"0000" when x"0173",
			x"0000" when x"0174",
			x"0000" when x"0175",
			x"0000" when x"0176",
			x"0000" when x"0177",
			x"0000" when x"0178",
			x"0000" when x"0179",
			x"0000" when x"017A",
			x"0000" when x"017B",
			x"0000" when x"017C",
			x"0000" when x"017D",
			x"0000" when x"017E",
			x"0000" when x"017F",
			x"0000" when x"0180",
			x"0000" when x"0181",
			x"0000" when x"0182",
			x"0000" when x"0183",
			x"0000" when x"0184",
			x"0000" when x"0185",
			x"0000" when x"0186",
			x"0000" when x"0187",
			x"0000" when x"0188",
			x"0000" when x"0189",
			x"0000" when x"018A",
			x"0000" when x"018B",
			x"0000" when x"018C",
			x"0000" when x"018D",
			x"0000" when x"018E",
			x"0000" when x"018F",
			x"0000" when x"0190",
			x"0000" when x"0191",
			x"0000" when x"0192",
			x"0000" when x"0193",
			x"0000" when x"0194",
			x"0000" when x"0195",
			x"0000" when x"0196",
			x"0000" when x"0197",
			x"0000" when x"0198",
			x"0000" when x"0199",
			x"0000" when x"019A",
			x"0000" when x"019B",
			x"0000" when x"019C",
			x"0000" when x"019D",
			x"0000" when x"019E",
			x"0000" when x"019F",
			x"0000" when x"01A0",
			x"0000" when x"01A1",
			x"0000" when x"01A2",
			x"0000" when x"01A3",
			x"0000" when x"01A4",
			x"0000" when x"01A5",
			x"0000" when x"01A6",
			x"0000" when x"01A7",
			x"0000" when x"01A8",
			x"0000" when x"01A9",
			x"0000" when x"01AA",
			x"0000" when x"01AB",
			x"0000" when x"01AC",
			x"0000" when x"01AD",
			x"0000" when x"01AE",
			x"0000" when x"01AF",
			x"0000" when x"01B0",
			x"0000" when x"01B1",
			x"0000" when x"01B2",
			x"0000" when x"01B3",
			x"0000" when x"01B4",
			x"0000" when x"01B5",
			x"0000" when x"01B6",
			x"0000" when x"01B7",
			x"0000" when x"01B8",
			x"0000" when x"01B9",
			x"0000" when x"01BA",
			x"0000" when x"01BB",
			x"0000" when x"01BC",
			x"0000" when x"01BD",
			x"0000" when x"01BE",
			x"0000" when x"01BF",
			x"0000" when x"01C0",
			x"0000" when x"01C1",
			x"0000" when x"01C2",
			x"0000" when x"01C3",
			x"0000" when x"01C4",
			x"0000" when x"01C5",
			x"0000" when x"01C6",
			x"0000" when x"01C7",
			x"0000" when x"01C8",
			x"0000" when x"01C9",
			x"0000" when x"01CA",
			x"0000" when x"01CB",
			x"0000" when x"01CC",
			x"0000" when x"01CD",
			x"0000" when x"01CE",
			x"0000" when x"01CF",
			x"0000" when x"01D0",
			x"0000" when x"01D1",
			x"0000" when x"01D2",
			x"0000" when x"01D3",
			x"0000" when x"01D4",
			x"0000" when x"01D5",
			x"0000" when x"01D6",
			x"0000" when x"01D7",
			x"0000" when x"01D8",
			x"0000" when x"01D9",
			x"0000" when x"01DA",
			x"0000" when x"01DB",
			x"0000" when x"01DC",
			x"0000" when x"01DD",
			x"0000" when x"01DE",
			x"0000" when x"01DF",
			x"0000" when x"01E0",
			x"0000" when x"01E1",
			x"0000" when x"01E2",
			x"0000" when x"01E3",
			x"0000" when x"01E4",
			x"0000" when x"01E5",
			x"0000" when x"01E6",
			x"0000" when x"01E7",
			x"0000" when x"01E8",
			x"0000" when x"01E9",
			x"0000" when x"01EA",
			x"0000" when x"01EB",
			x"0000" when x"01EC",
			x"0000" when x"01ED",
			x"0000" when x"01EE",
			x"0000" when x"01EF",
			x"0000" when x"01F0",
			x"0000" when x"01F1",
			x"0000" when x"01F2",
			x"0000" when x"01F3",
			x"0000" when x"01F4",
			x"0000" when x"01F5",
			x"0000" when x"01F6",
			x"0000" when x"01F7",
			x"0000" when x"01F8",
			x"0000" when x"01F9",
			x"0000" when x"01FA",
			x"0000" when x"01FB",
			x"0000" when x"01FC",
			x"0000" when x"01FD",
			x"0000" when x"01FE",
			x"0000" when x"01FF",
			x"0000" when x"0200",
			x"0000" when x"0201",
			x"0000" when x"0202",
			x"0000" when x"0203",
			x"0000" when x"0204",
			x"0000" when x"0205",
			x"0000" when x"0206",
			x"0000" when x"0207",
			x"0000" when x"0208",
			x"0000" when x"0209",
			x"0000" when x"020A",
			x"0000" when x"020B",
			x"0000" when x"020C",
			x"0000" when x"020D",
			x"0000" when x"020E",
			x"0000" when x"020F",
			x"0000" when x"0210",
			x"0000" when x"0211",
			x"0000" when x"0212",
			x"0000" when x"0213",
			x"0000" when x"0214",
			x"0000" when x"0215",
			x"0000" when x"0216",
			x"0000" when x"0217",
			x"0000" when x"0218",
			x"0000" when x"0219",
			x"0000" when x"021A",
			x"0000" when x"021B",
			x"0000" when x"021C",
			x"0000" when x"021D",
			x"0000" when x"021E",
			x"0000" when x"021F",
			x"0000" when x"0220",
			x"0000" when x"0221",
			x"0000" when x"0222",
			x"0000" when x"0223",
			x"0000" when x"0224",
			x"0000" when x"0225",
			x"0000" when x"0226",
			x"0000" when x"0227",
			x"0000" when x"0228",
			x"0000" when x"0229",
			x"0000" when x"022A",
			x"0000" when x"022B",
			x"0000" when x"022C",
			x"0000" when x"022D",
			x"0000" when x"022E",
			x"0000" when x"022F",
			x"0000" when x"0230",
			x"0000" when x"0231",
			x"0000" when x"0232",
			x"0000" when x"0233",
			x"0000" when x"0234",
			x"0000" when x"0235",
			x"0000" when x"0236",
			x"0000" when x"0237",
			x"0000" when x"0238",
			x"0000" when x"0239",
			x"0000" when x"023A",
			x"0000" when x"023B",
			x"0000" when x"023C",
			x"0000" when x"023D",
			x"0000" when x"023E",
			x"0000" when x"023F",
			x"0000" when x"0240",
			x"0000" when x"0241",
			x"0000" when x"0242",
			x"0000" when x"0243",
			x"0000" when x"0244",
			x"0000" when x"0245",
			x"0000" when x"0246",
			x"0000" when x"0247",
			x"0000" when x"0248",
			x"0000" when x"0249",
			x"0000" when x"024A",
			x"0000" when x"024B",
			x"0000" when x"024C",
			x"0000" when x"024D",
			x"0000" when x"024E",
			x"0000" when x"024F",
			x"0000" when x"0250",
			x"0000" when x"0251",
			x"0000" when x"0252",
			x"0000" when x"0253",
			x"0000" when x"0254",
			x"0000" when x"0255",
			x"0000" when x"0256",
			x"0000" when x"0257",
			x"0000" when x"0258",
			x"0000" when x"0259",
			x"0000" when x"025A",
			x"0000" when x"025B",
			x"0000" when x"025C",
			x"0000" when x"025D",
			x"0000" when x"025E",
			x"0000" when x"025F",
			x"0000" when x"0260",
			x"0000" when x"0261",
			x"0000" when x"0262",
			x"0000" when x"0263",
			x"0000" when x"0264",
			x"0000" when x"0265",
			x"0000" when x"0266",
			x"0000" when x"0267",
			x"0000" when x"0268",
			x"0000" when x"0269",
			x"0000" when x"026A",
			x"0000" when x"026B",
			x"0000" when x"026C",
			x"0000" when x"026D",
			x"0000" when x"026E",
			x"0000" when x"026F",
			x"0000" when x"0270",
			x"0000" when x"0271",
			x"0000" when x"0272",
			x"0000" when x"0273",
			x"0000" when x"0274",
			x"0000" when x"0275",
			x"0000" when x"0276",
			x"0000" when x"0277",
			x"0000" when x"0278",
			x"0000" when x"0279",
			x"0000" when x"027A",
			x"0000" when x"027B",
			x"0000" when x"027C",
			x"0000" when x"027D",
			x"0000" when x"027E",
			x"0000" when x"027F",
			x"0000" when x"0280",
			x"0000" when x"0281",
			x"0000" when x"0282",
			x"0000" when x"0283",
			x"0000" when x"0284",
			x"0000" when x"0285",
			x"0000" when x"0286",
			x"0000" when x"0287",
			x"0000" when x"0288",
			x"0000" when x"0289",
			x"0000" when x"028A",
			x"0000" when x"028B",
			x"0000" when x"028C",
			x"0000" when x"028D",
			x"0000" when x"028E",
			x"0000" when x"028F",
			x"0000" when x"0290",
			x"0000" when x"0291",
			x"0000" when x"0292",
			x"0000" when x"0293",
			x"0000" when x"0294",
			x"0000" when x"0295",
			x"0000" when x"0296",
			x"0000" when x"0297",
			x"0000" when x"0298",
			x"0000" when x"0299",
			x"0000" when x"029A",
			x"0000" when x"029B",
			x"0000" when x"029C",
			x"0000" when x"029D",
			x"0000" when x"029E",
			x"0000" when x"029F",
			x"0000" when x"02A0",
			x"0000" when x"02A1",
			x"0000" when x"02A2",
			x"0000" when x"02A3",
			x"0000" when x"02A4",
			x"0000" when x"02A5",
			x"0000" when x"02A6",
			x"0000" when x"02A7",
			x"0000" when x"02A8",
			x"0000" when x"02A9",
			x"0000" when x"02AA",
			x"0000" when x"02AB",
			x"0000" when x"02AC",
			x"0000" when x"02AD",
			x"0000" when x"02AE",
			x"0000" when x"02AF",
			x"0000" when x"02B0",
			x"0000" when x"02B1",
			x"0000" when x"02B2",
			x"0000" when x"02B3",
			x"0000" when x"02B4",
			x"0000" when x"02B5",
			x"0000" when x"02B6",
			x"0000" when x"02B7",
			x"0000" when x"02B8",
			x"0000" when x"02B9",
			x"0000" when x"02BA",
			x"0000" when x"02BB",
			x"0000" when x"02BC",
			x"0000" when x"02BD",
			x"0000" when x"02BE",
			x"0000" when x"02BF",
			x"0000" when x"02C0",
			x"0000" when x"02C1",
			x"0000" when x"02C2",
			x"0000" when x"02C3",
			x"0000" when x"02C4",
			x"0000" when x"02C5",
			x"0000" when x"02C6",
			x"0000" when x"02C7",
			x"0000" when x"02C8",
			x"0000" when x"02C9",
			x"0000" when x"02CA",
			x"0000" when x"02CB",
			x"0000" when x"02CC",
			x"0000" when x"02CD",
			x"0000" when x"02CE",
			x"0000" when x"02CF",
			x"0000" when x"02D0",
			x"0000" when x"02D1",
			x"0000" when x"02D2",
			x"0000" when x"02D3",
			x"0000" when x"02D4",
			x"0000" when x"02D5",
			x"0000" when x"02D6",
			x"0000" when x"02D7",
			x"0000" when x"02D8",
			x"0000" when x"02D9",
			x"0000" when x"02DA",
			x"0000" when x"02DB",
			x"0000" when x"02DC",
			x"0000" when x"02DD",
			x"0000" when x"02DE",
			x"0000" when x"02DF",
			x"0000" when x"02E0",
			x"0000" when x"02E1",
			x"0000" when x"02E2",
			x"0000" when x"02E3",
			x"0000" when x"02E4",
			x"0000" when x"02E5",
			x"0000" when x"02E6",
			x"0000" when x"02E7",
			x"0000" when x"02E8",
			x"0000" when x"02E9",
			x"0000" when x"02EA",
			x"0000" when x"02EB",
			x"0000" when x"02EC",
			x"0000" when x"02ED",
			x"0000" when x"02EE",
			x"0000" when x"02EF",
			x"0000" when x"02F0",
			x"0000" when x"02F1",
			x"0000" when x"02F2",
			x"0000" when x"02F3",
			x"0000" when x"02F4",
			x"0000" when x"02F5",
			x"0000" when x"02F6",
			x"0000" when x"02F7",
			x"0000" when x"02F8",
			x"0000" when x"02F9",
			x"0000" when x"02FA",
			x"0000" when x"02FB",
			x"0000" when x"02FC",
			x"0000" when x"02FD",
			x"0000" when x"02FE",
			x"0000" when x"02FF",
			x"0000" when x"0300",
			x"0000" when x"0301",
			x"0000" when x"0302",
			x"0000" when x"0303",
			x"0000" when x"0304",
			x"0000" when x"0305",
			x"0000" when x"0306",
			x"0000" when x"0307",
			x"0000" when x"0308",
			x"0000" when x"0309",
			x"0000" when x"030A",
			x"0000" when x"030B",
			x"0000" when x"030C",
			x"0000" when x"030D",
			x"0000" when x"030E",
			x"0000" when x"030F",
			x"0000" when x"0310",
			x"0000" when x"0311",
			x"0000" when x"0312",
			x"0000" when x"0313",
			x"0000" when x"0314",
			x"0000" when x"0315",
			x"0000" when x"0316",
			x"0000" when x"0317",
			x"0000" when x"0318",
			x"0000" when x"0319",
			x"0000" when x"031A",
			x"0000" when x"031B",
			x"0000" when x"031C",
			x"0000" when x"031D",
			x"0000" when x"031E",
			x"0000" when x"031F",
			x"0000" when x"0320",
			x"0000" when x"0321",
			x"0000" when x"0322",
			x"0000" when x"0323",
			x"0000" when x"0324",
			x"0000" when x"0325",
			x"0000" when x"0326",
			x"0000" when x"0327",
			x"0000" when x"0328",
			x"0000" when x"0329",
			x"0000" when x"032A",
			x"0000" when x"032B",
			x"0000" when x"032C",
			x"0000" when x"032D",
			x"0000" when x"032E",
			x"0000" when x"032F",
			x"0000" when x"0330",
			x"0000" when x"0331",
			x"0000" when x"0332",
			x"0000" when x"0333",
			x"0000" when x"0334",
			x"0000" when x"0335",
			x"0000" when x"0336",
			x"0000" when x"0337",
			x"0000" when x"0338",
			x"0000" when x"0339",
			x"0000" when x"033A",
			x"0000" when x"033B",
			x"0000" when x"033C",
			x"0000" when x"033D",
			x"0000" when x"033E",
			x"0000" when x"033F",
			x"0000" when x"0340",
			x"0000" when x"0341",
			x"0000" when x"0342",
			x"0000" when x"0343",
			x"0000" when x"0344",
			x"0000" when x"0345",
			x"0000" when x"0346",
			x"0000" when x"0347",
			x"0000" when x"0348",
			x"0000" when x"0349",
			x"0000" when x"034A",
			x"0000" when x"034B",
			x"0000" when x"034C",
			x"0000" when x"034D",
			x"0000" when x"034E",
			x"0000" when x"034F",
			x"0000" when x"0350",
			x"0000" when x"0351",
			x"0000" when x"0352",
			x"0000" when x"0353",
			x"0000" when x"0354",
			x"0000" when x"0355",
			x"0000" when x"0356",
			x"0000" when x"0357",
			x"0000" when x"0358",
			x"0000" when x"0359",
			x"0000" when x"035A",
			x"0000" when x"035B",
			x"0000" when x"035C",
			x"0000" when x"035D",
			x"0000" when x"035E",
			x"0000" when x"035F",
			x"0000" when x"0360",
			x"0000" when x"0361",
			x"0000" when x"0362",
			x"0000" when x"0363",
			x"0000" when x"0364",
			x"0000" when x"0365",
			x"0000" when x"0366",
			x"0000" when x"0367",
			x"0000" when x"0368",
			x"0000" when x"0369",
			x"0000" when x"036A",
			x"0000" when x"036B",
			x"0000" when x"036C",
			x"0000" when x"036D",
			x"0000" when x"036E",
			x"0000" when x"036F",
			x"0000" when x"0370",
			x"0000" when x"0371",
			x"0000" when x"0372",
			x"0000" when x"0373",
			x"0000" when x"0374",
			x"0000" when x"0375",
			x"0000" when x"0376",
			x"0000" when x"0377",
			x"0000" when x"0378",
			x"0000" when x"0379",
			x"0000" when x"037A",
			x"0000" when x"037B",
			x"0000" when x"037C",
			x"0000" when x"037D",
			x"0000" when x"037E",
			x"0000" when x"037F",
			x"0000" when x"0380",
			x"0000" when x"0381",
			x"0000" when x"0382",
			x"0000" when x"0383",
			x"0000" when x"0384",
			x"0000" when x"0385",
			x"0000" when x"0386",
			x"0000" when x"0387",
			x"0000" when x"0388",
			x"0000" when x"0389",
			x"0000" when x"038A",
			x"0000" when x"038B",
			x"0000" when x"038C",
			x"0000" when x"038D",
			x"0000" when x"038E",
			x"0000" when x"038F",
			x"0000" when x"0390",
			x"0000" when x"0391",
			x"0000" when x"0392",
			x"0000" when x"0393",
			x"0000" when x"0394",
			x"0000" when x"0395",
			x"0000" when x"0396",
			x"0000" when x"0397",
			x"0000" when x"0398",
			x"0000" when x"0399",
			x"0000" when x"039A",
			x"0000" when x"039B",
			x"0000" when x"039C",
			x"0000" when x"039D",
			x"0000" when x"039E",
			x"0000" when x"039F",
			x"0000" when x"03A0",
			x"0000" when x"03A1",
			x"0000" when x"03A2",
			x"0000" when x"03A3",
			x"0000" when x"03A4",
			x"0000" when x"03A5",
			x"0000" when x"03A6",
			x"0000" when x"03A7",
			x"0000" when x"03A8",
			x"0000" when x"03A9",
			x"0000" when x"03AA",
			x"0000" when x"03AB",
			x"0000" when x"03AC",
			x"0000" when x"03AD",
			x"0000" when x"03AE",
			x"0000" when x"03AF",
			x"0000" when x"03B0",
			x"0000" when x"03B1",
			x"0000" when x"03B2",
			x"0000" when x"03B3",
			x"0000" when x"03B4",
			x"0000" when x"03B5",
			x"0000" when x"03B6",
			x"0000" when x"03B7",
			x"0000" when x"03B8",
			x"0000" when x"03B9",
			x"0000" when x"03BA",
			x"0000" when x"03BB",
			x"0000" when x"03BC",
			x"0000" when x"03BD",
			x"0000" when x"03BE",
			x"0000" when x"03BF",
			x"0000" when x"03C0",
			x"0000" when x"03C1",
			x"0000" when x"03C2",
			x"0000" when x"03C3",
			x"0000" when x"03C4",
			x"0000" when x"03C5",
			x"0000" when x"03C6",
			x"0000" when x"03C7",
			x"0000" when x"03C8",
			x"0000" when x"03C9",
			x"0000" when x"03CA",
			x"0000" when x"03CB",
			x"0000" when x"03CC",
			x"0000" when x"03CD",
			x"0000" when x"03CE",
			x"0000" when x"03CF",
			x"0000" when x"03D0",
			x"0000" when x"03D1",
			x"0000" when x"03D2",
			x"0000" when x"03D3",
			x"0000" when x"03D4",
			x"0000" when x"03D5",
			x"0000" when x"03D6",
			x"0000" when x"03D7",
			x"0000" when x"03D8",
			x"0000" when x"03D9",
			x"0000" when x"03DA",
			x"0000" when x"03DB",
			x"0000" when x"03DC",
			x"0000" when x"03DD",
			x"0000" when x"03DE",
			x"0000" when x"03DF",
			x"0000" when x"03E0",
			x"0000" when x"03E1",
			x"0000" when x"03E2",
			x"0000" when x"03E3",
			x"0000" when x"03E4",
			x"0000" when x"03E5",
			x"0000" when x"03E6",
			x"0000" when x"03E7",
			x"0000" when x"03E8",
			x"0000" when x"03E9",
			x"0000" when x"03EA",
			x"0000" when x"03EB",
			x"0000" when x"03EC",
			x"0000" when x"03ED",
			x"0000" when x"03EE",
			x"0000" when x"03EF",
			x"0000" when x"03F0",
			x"0000" when x"03F1",
			x"0000" when x"03F2",
			x"0000" when x"03F3",
			x"0000" when x"03F4",
			x"0000" when x"03F5",
			x"0000" when x"03F6",
			x"0000" when x"03F7",
			x"0000" when x"03F8",
			x"0000" when x"03F9",
			x"0000" when x"03FA",
			x"0000" when x"03FB",
			x"0000" when x"03FC",
			x"0000" when x"03FD",
			x"0000" when x"03FE",
			x"0000" when x"03FF",
			x"0000" when x"0400",
			x"0000" when x"0401",
			x"0000" when x"0402",
			x"0000" when x"0403",
			x"0000" when x"0404",
			x"0000" when x"0405",
			x"0000" when x"0406",
			x"0000" when x"0407",
			x"0000" when x"0408",
			x"0000" when x"0409",
			x"0000" when x"040A",
			x"0000" when x"040B",
			x"0000" when x"040C",
			x"0000" when x"040D",
			x"0000" when x"040E",
			x"0000" when x"040F",
			x"0000" when x"0410",
			x"0000" when x"0411",
			x"0000" when x"0412",
			x"0000" when x"0413",
			x"0000" when x"0414",
			x"0000" when x"0415",
			x"0000" when x"0416",
			x"0000" when x"0417",
			x"0000" when x"0418",
			x"0000" when x"0419",
			x"0000" when x"041A",
			x"0000" when x"041B",
			x"0000" when x"041C",
			x"0000" when x"041D",
			x"0000" when x"041E",
			x"0000" when x"041F",
			x"0000" when x"0420",
			x"0000" when x"0421",
			x"0000" when x"0422",
			x"0000" when x"0423",
			x"0000" when x"0424",
			x"0000" when x"0425",
			x"0000" when x"0426",
			x"0000" when x"0427",
			x"0000" when x"0428",
			x"0000" when x"0429",
			x"0000" when x"042A",
			x"0000" when x"042B",
			x"0000" when x"042C",
			x"0000" when x"042D",
			x"0000" when x"042E",
			x"0000" when x"042F",
			x"0000" when x"0430",
			x"0000" when x"0431",
			x"0000" when x"0432",
			x"0000" when x"0433",
			x"0000" when x"0434",
			x"0000" when x"0435",
			x"0000" when x"0436",
			x"0000" when x"0437",
			x"0000" when x"0438",
			x"0000" when x"0439",
			x"0000" when x"043A",
			x"0000" when x"043B",
			x"0000" when x"043C",
			x"0000" when x"043D",
			x"0000" when x"043E",
			x"0000" when x"043F",
			x"0000" when x"0440",
			x"0000" when x"0441",
			x"0000" when x"0442",
			x"0000" when x"0443",
			x"0000" when x"0444",
			x"0000" when x"0445",
			x"0000" when x"0446",
			x"0000" when x"0447",
			x"0000" when x"0448",
			x"0000" when x"0449",
			x"0000" when x"044A",
			x"0000" when x"044B",
			x"0000" when x"044C",
			x"0000" when x"044D",
			x"0000" when x"044E",
			x"0000" when x"044F",
			x"0000" when x"0450",
			x"0000" when x"0451",
			x"0000" when x"0452",
			x"0000" when x"0453",
			x"0000" when x"0454",
			x"0000" when x"0455",
			x"0000" when x"0456",
			x"0000" when x"0457",
			x"0000" when x"0458",
			x"0000" when x"0459",
			x"0000" when x"045A",
			x"0000" when x"045B",
			x"0000" when x"045C",
			x"0000" when x"045D",
			x"0000" when x"045E",
			x"0000" when x"045F",
			x"0000" when x"0460",
			x"0000" when x"0461",
			x"0000" when x"0462",
			x"0000" when x"0463",
			x"0000" when x"0464",
			x"0000" when x"0465",
			x"0000" when x"0466",
			x"0000" when x"0467",
			x"0000" when x"0468",
			x"0000" when x"0469",
			x"0000" when x"046A",
			x"0000" when x"046B",
			x"0000" when x"046C",
			x"0000" when x"046D",
			x"0000" when x"046E",
			x"0000" when x"046F",
			x"0000" when x"0470",
			x"0000" when x"0471",
			x"0000" when x"0472",
			x"0000" when x"0473",
			x"0000" when x"0474",
			x"0000" when x"0475",
			x"0000" when x"0476",
			x"0000" when x"0477",
			x"0000" when x"0478",
			x"0000" when x"0479",
			x"0000" when x"047A",
			x"0000" when x"047B",
			x"0000" when x"047C",
			x"0000" when x"047D",
			x"0000" when x"047E",
			x"0000" when x"047F",
			x"0000" when x"0480",
			x"0000" when x"0481",
			x"0000" when x"0482",
			x"0000" when x"0483",
			x"0000" when x"0484",
			x"0000" when x"0485",
			x"0000" when x"0486",
			x"0000" when x"0487",
			x"0000" when x"0488",
			x"0000" when x"0489",
			x"0000" when x"048A",
			x"0000" when x"048B",
			x"0000" when x"048C",
			x"0000" when x"048D",
			x"0000" when x"048E",
			x"0000" when x"048F",
			x"0000" when x"0490",
			x"0000" when x"0491",
			x"0000" when x"0492",
			x"0000" when x"0493",
			x"0000" when x"0494",
			x"0000" when x"0495",
			x"0000" when x"0496",
			x"0000" when x"0497",
			x"0000" when x"0498",
			x"0000" when x"0499",
			x"0000" when x"049A",
			x"0000" when x"049B",
			x"0000" when x"049C",
			x"0000" when x"049D",
			x"0000" when x"049E",
			x"0000" when x"049F",
			x"0000" when x"04A0",
			x"0000" when x"04A1",
			x"0000" when x"04A2",
			x"0000" when x"04A3",
			x"0000" when x"04A4",
			x"0000" when x"04A5",
			x"0000" when x"04A6",
			x"0000" when x"04A7",
			x"0000" when x"04A8",
			x"0000" when x"04A9",
			x"0000" when x"04AA",
			x"0000" when x"04AB",
			x"0000" when x"04AC",
			x"0000" when x"04AD",
			x"0000" when x"04AE",
			x"0000" when x"04AF",
			x"0000" when x"04B0",
			x"0000" when x"04B1",
			x"0000" when x"04B2",
			x"0000" when x"04B3",
			x"0000" when x"04B4",
			x"0000" when x"04B5",
			x"0000" when x"04B6",
			x"0000" when x"04B7",
			x"0000" when x"04B8",
			x"0000" when x"04B9",
			x"0000" when x"04BA",
			x"0000" when x"04BB",
			x"0000" when x"04BC",
			x"0000" when x"04BD",
			x"0000" when x"04BE",
			x"0000" when x"04BF",
			x"0000" when x"04C0",
			x"0000" when x"04C1",
			x"0000" when x"04C2",
			x"0000" when x"04C3",
			x"0000" when x"04C4",
			x"0000" when x"04C5",
			x"0000" when x"04C6",
			x"0000" when x"04C7",
			x"0000" when x"04C8",
			x"0000" when x"04C9",
			x"0000" when x"04CA",
			x"0000" when x"04CB",
			x"0000" when x"04CC",
			x"0000" when x"04CD",
			x"0000" when x"04CE",
			x"0000" when x"04CF",
			x"0000" when x"04D0",
			x"0000" when x"04D1",
			x"0000" when x"04D2",
			x"0000" when x"04D3",
			x"0000" when x"04D4",
			x"0000" when x"04D5",
			x"0000" when x"04D6",
			x"0000" when x"04D7",
			x"0000" when x"04D8",
			x"0000" when x"04D9",
			x"0000" when x"04DA",
			x"0000" when x"04DB",
			x"0000" when x"04DC",
			x"0000" when x"04DD",
			x"0000" when x"04DE",
			x"0000" when x"04DF",
			x"0000" when x"04E0",
			x"0000" when x"04E1",
			x"0000" when x"04E2",
			x"0000" when x"04E3",
			x"0000" when x"04E4",
			x"0000" when x"04E5",
			x"0000" when x"04E6",
			x"0000" when x"04E7",
			x"0000" when x"04E8",
			x"0000" when x"04E9",
			x"0000" when x"04EA",
			x"0000" when x"04EB",
			x"0000" when x"04EC",
			x"0000" when x"04ED",
			x"0000" when x"04EE",
			x"0000" when x"04EF",
			x"0000" when x"04F0",
			x"0000" when x"04F1",
			x"0000" when x"04F2",
			x"0000" when x"04F3",
			x"0000" when x"04F4",
			x"0000" when x"04F5",
			x"0000" when x"04F6",
			x"0000" when x"04F7",
			x"0000" when x"04F8",
			x"0000" when x"04F9",
			x"0000" when x"04FA",
			x"0000" when x"04FB",
			x"0000" when x"04FC",
			x"0000" when x"04FD",
			x"0000" when x"04FE",
			x"0000" when x"04FF",
			x"0000" when x"0500",
			x"0000" when x"0501",
			x"0000" when x"0502",
			x"0000" when x"0503",
			x"0000" when x"0504",
			x"0000" when x"0505",
			x"0000" when x"0506",
			x"0000" when x"0507",
			x"0000" when x"0508",
			x"0000" when x"0509",
			x"0000" when x"050A",
			x"0000" when x"050B",
			x"0000" when x"050C",
			x"0000" when x"050D",
			x"0000" when x"050E",
			x"0000" when x"050F",
			x"0000" when x"0510",
			x"0000" when x"0511",
			x"0000" when x"0512",
			x"0000" when x"0513",
			x"0000" when x"0514",
			x"0000" when x"0515",
			x"0000" when x"0516",
			x"0000" when x"0517",
			x"0000" when x"0518",
			x"0000" when x"0519",
			x"0000" when x"051A",
			x"0000" when x"051B",
			x"0000" when x"051C",
			x"0000" when x"051D",
			x"0000" when x"051E",
			x"0000" when x"051F",
			x"0000" when x"0520",
			x"0000" when x"0521",
			x"0000" when x"0522",
			x"0000" when x"0523",
			x"0000" when x"0524",
			x"0000" when x"0525",
			x"0000" when x"0526",
			x"0000" when x"0527",
			x"0000" when x"0528",
			x"0000" when x"0529",
			x"0000" when x"052A",
			x"0000" when x"052B",
			x"0000" when x"052C",
			x"0000" when x"052D",
			x"0000" when x"052E",
			x"0000" when x"052F",
			x"0000" when x"0530",
			x"0000" when x"0531",
			x"0000" when x"0532",
			x"0000" when x"0533",
			x"0000" when x"0534",
			x"0000" when x"0535",
			x"0000" when x"0536",
			x"0000" when x"0537",
			x"0000" when x"0538",
			x"0000" when x"0539",
			x"0000" when x"053A",
			x"0000" when x"053B",
			x"0000" when x"053C",
			x"0000" when x"053D",
			x"0000" when x"053E",
			x"0000" when x"053F",
			x"0000" when x"0540",
			x"0000" when x"0541",
			x"0000" when x"0542",
			x"0000" when x"0543",
			x"0000" when x"0544",
			x"0000" when x"0545",
			x"0000" when x"0546",
			x"0000" when x"0547",
			x"0000" when x"0548",
			x"0000" when x"0549",
			x"0000" when x"054A",
			x"0000" when x"054B",
			x"0000" when x"054C",
			x"0000" when x"054D",
			x"0000" when x"054E",
			x"0000" when x"054F",
			x"0000" when x"0550",
			x"0000" when x"0551",
			x"0000" when x"0552",
			x"0000" when x"0553",
			x"0000" when x"0554",
			x"0000" when x"0555",
			x"0000" when x"0556",
			x"0000" when x"0557",
			x"0000" when x"0558",
			x"0000" when x"0559",
			x"0000" when x"055A",
			x"0000" when x"055B",
			x"0000" when x"055C",
			x"0000" when x"055D",
			x"0000" when x"055E",
			x"0000" when x"055F",
			x"0000" when x"0560",
			x"0000" when x"0561",
			x"0000" when x"0562",
			x"0000" when x"0563",
			x"0000" when x"0564",
			x"0000" when x"0565",
			x"0000" when x"0566",
			x"0000" when x"0567",
			x"0000" when x"0568",
			x"0000" when x"0569",
			x"0000" when x"056A",
			x"0000" when x"056B",
			x"0000" when x"056C",
			x"0000" when x"056D",
			x"0000" when x"056E",
			x"0000" when x"056F",
			x"0000" when x"0570",
			x"0000" when x"0571",
			x"0000" when x"0572",
			x"0000" when x"0573",
			x"0000" when x"0574",
			x"0000" when x"0575",
			x"0000" when x"0576",
			x"0000" when x"0577",
			x"0000" when x"0578",
			x"0000" when x"0579",
			x"0000" when x"057A",
			x"0000" when x"057B",
			x"0000" when x"057C",
			x"0000" when x"057D",
			x"0000" when x"057E",
			x"0000" when x"057F",
			x"0000" when x"0580",
			x"0000" when x"0581",
			x"0000" when x"0582",
			x"0000" when x"0583",
			x"0000" when x"0584",
			x"0000" when x"0585",
			x"0000" when x"0586",
			x"0000" when x"0587",
			x"0000" when x"0588",
			x"0000" when x"0589",
			x"0000" when x"058A",
			x"0000" when x"058B",
			x"0000" when x"058C",
			x"0000" when x"058D",
			x"0000" when x"058E",
			x"0000" when x"058F",
			x"0000" when x"0590",
			x"0000" when x"0591",
			x"0000" when x"0592",
			x"0000" when x"0593",
			x"0000" when x"0594",
			x"0000" when x"0595",
			x"0000" when x"0596",
			x"0000" when x"0597",
			x"0000" when x"0598",
			x"0000" when x"0599",
			x"0000" when x"059A",
			x"0000" when x"059B",
			x"0000" when x"059C",
			x"0000" when x"059D",
			x"0000" when x"059E",
			x"0000" when x"059F",
			x"0000" when x"05A0",
			x"0000" when x"05A1",
			x"0000" when x"05A2",
			x"0000" when x"05A3",
			x"0000" when x"05A4",
			x"0000" when x"05A5",
			x"0000" when x"05A6",
			x"0000" when x"05A7",
			x"0000" when x"05A8",
			x"0000" when x"05A9",
			x"0000" when x"05AA",
			x"0000" when x"05AB",
			x"0000" when x"05AC",
			x"0000" when x"05AD",
			x"0000" when x"05AE",
			x"0000" when x"05AF",
			x"0000" when x"05B0",
			x"0000" when x"05B1",
			x"0000" when x"05B2",
			x"0000" when x"05B3",
			x"0000" when x"05B4",
			x"0000" when x"05B5",
			x"0000" when x"05B6",
			x"0000" when x"05B7",
			x"0000" when x"05B8",
			x"0000" when x"05B9",
			x"0000" when x"05BA",
			x"0000" when x"05BB",
			x"0000" when x"05BC",
			x"0000" when x"05BD",
			x"0000" when x"05BE",
			x"0000" when x"05BF",
			x"0000" when x"05C0",
			x"0000" when x"05C1",
			x"0000" when x"05C2",
			x"0000" when x"05C3",
			x"0000" when x"05C4",
			x"0000" when x"05C5",
			x"0000" when x"05C6",
			x"0000" when x"05C7",
			x"0000" when x"05C8",
			x"0000" when x"05C9",
			x"0000" when x"05CA",
			x"0000" when x"05CB",
			x"0000" when x"05CC",
			x"0000" when x"05CD",
			x"0000" when x"05CE",
			x"0000" when x"05CF",
			x"0000" when x"05D0",
			x"0000" when x"05D1",
			x"0000" when x"05D2",
			x"0000" when x"05D3",
			x"0000" when x"05D4",
			x"0000" when x"05D5",
			x"0000" when x"05D6",
			x"0000" when x"05D7",
			x"0000" when x"05D8",
			x"0000" when x"05D9",
			x"0000" when x"05DA",
			x"0000" when x"05DB",
			x"0000" when x"05DC",
			x"0000" when x"05DD",
			x"0000" when x"05DE",
			x"0000" when x"05DF",
			x"0000" when x"05E0",
			x"0000" when x"05E1",
			x"0000" when x"05E2",
			x"0000" when x"05E3",
			x"0000" when x"05E4",
			x"0000" when x"05E5",
			x"0000" when x"05E6",
			x"0000" when x"05E7",
			x"0000" when x"05E8",
			x"0000" when x"05E9",
			x"0000" when x"05EA",
			x"0000" when x"05EB",
			x"0000" when x"05EC",
			x"0000" when x"05ED",
			x"0000" when x"05EE",
			x"0000" when x"05EF",
			x"0000" when x"05F0",
			x"0000" when x"05F1",
			x"0000" when x"05F2",
			x"0000" when x"05F3",
			x"0000" when x"05F4",
			x"0000" when x"05F5",
			x"0000" when x"05F6",
			x"0000" when x"05F7",
			x"0000" when x"05F8",
			x"0000" when x"05F9",
			x"0000" when x"05FA",
			x"0000" when x"05FB",
			x"0000" when x"05FC",
			x"0000" when x"05FD",
			x"0000" when x"05FE",
			x"0000" when x"05FF",
			x"0000" when x"0600",
			x"0000" when x"0601",
			x"0000" when x"0602",
			x"0000" when x"0603",
			x"0000" when x"0604",
			x"0000" when x"0605",
			x"0000" when x"0606",
			x"0000" when x"0607",
			x"0000" when x"0608",
			x"0000" when x"0609",
			x"0000" when x"060A",
			x"0000" when x"060B",
			x"0000" when x"060C",
			x"0000" when x"060D",
			x"0000" when x"060E",
			x"0000" when x"060F",
			x"0000" when x"0610",
			x"0000" when x"0611",
			x"0000" when x"0612",
			x"0000" when x"0613",
			x"0000" when x"0614",
			x"0000" when x"0615",
			x"0000" when x"0616",
			x"0000" when x"0617",
			x"0000" when x"0618",
			x"0000" when x"0619",
			x"0000" when x"061A",
			x"0000" when x"061B",
			x"0000" when x"061C",
			x"0000" when x"061D",
			x"0000" when x"061E",
			x"0000" when x"061F",
			x"0000" when x"0620",
			x"0000" when x"0621",
			x"0000" when x"0622",
			x"0000" when x"0623",
			x"0000" when x"0624",
			x"0000" when x"0625",
			x"0000" when x"0626",
			x"0000" when x"0627",
			x"0000" when x"0628",
			x"0000" when x"0629",
			x"0000" when x"062A",
			x"0000" when x"062B",
			x"0000" when x"062C",
			x"0000" when x"062D",
			x"0000" when x"062E",
			x"0000" when x"062F",
			x"0000" when x"0630",
			x"0000" when x"0631",
			x"0000" when x"0632",
			x"0000" when x"0633",
			x"0000" when x"0634",
			x"0000" when x"0635",
			x"0000" when x"0636",
			x"0000" when x"0637",
			x"0000" when x"0638",
			x"0000" when x"0639",
			x"0000" when x"063A",
			x"0000" when x"063B",
			x"0000" when x"063C",
			x"0000" when x"063D",
			x"0000" when x"063E",
			x"0000" when x"063F",
			x"0000" when x"0640",
			x"0000" when x"0641",
			x"0000" when x"0642",
			x"0000" when x"0643",
			x"0000" when x"0644",
			x"0000" when x"0645",
			x"0000" when x"0646",
			x"0000" when x"0647",
			x"0000" when x"0648",
			x"0000" when x"0649",
			x"0000" when x"064A",
			x"0000" when x"064B",
			x"0000" when x"064C",
			x"0000" when x"064D",
			x"0000" when x"064E",
			x"0000" when x"064F",
			x"0000" when x"0650",
			x"0000" when x"0651",
			x"0000" when x"0652",
			x"0000" when x"0653",
			x"0000" when x"0654",
			x"0000" when x"0655",
			x"0000" when x"0656",
			x"0000" when x"0657",
			x"0000" when x"0658",
			x"0000" when x"0659",
			x"0000" when x"065A",
			x"0000" when x"065B",
			x"0000" when x"065C",
			x"0000" when x"065D",
			x"0000" when x"065E",
			x"0000" when x"065F",
			x"0000" when x"0660",
			x"0000" when x"0661",
			x"0000" when x"0662",
			x"0000" when x"0663",
			x"0000" when x"0664",
			x"0000" when x"0665",
			x"0000" when x"0666",
			x"0000" when x"0667",
			x"0000" when x"0668",
			x"0000" when x"0669",
			x"0000" when x"066A",
			x"0000" when x"066B",
			x"0000" when x"066C",
			x"0000" when x"066D",
			x"0000" when x"066E",
			x"0000" when x"066F",
			x"0000" when x"0670",
			x"0000" when x"0671",
			x"0000" when x"0672",
			x"0000" when x"0673",
			x"0000" when x"0674",
			x"0000" when x"0675",
			x"0000" when x"0676",
			x"0000" when x"0677",
			x"0000" when x"0678",
			x"0000" when x"0679",
			x"0000" when x"067A",
			x"0000" when x"067B",
			x"0000" when x"067C",
			x"0000" when x"067D",
			x"0000" when x"067E",
			x"0000" when x"067F",
			x"0000" when x"0680",
			x"0000" when x"0681",
			x"0000" when x"0682",
			x"0000" when x"0683",
			x"0000" when x"0684",
			x"0000" when x"0685",
			x"0000" when x"0686",
			x"0000" when x"0687",
			x"0000" when x"0688",
			x"0000" when x"0689",
			x"0000" when x"068A",
			x"0000" when x"068B",
			x"0000" when x"068C",
			x"0000" when x"068D",
			x"0000" when x"068E",
			x"0000" when x"068F",
			x"0000" when x"0690",
			x"0000" when x"0691",
			x"0000" when x"0692",
			x"0000" when x"0693",
			x"0000" when x"0694",
			x"0000" when x"0695",
			x"0000" when x"0696",
			x"0000" when x"0697",
			x"0000" when x"0698",
			x"0000" when x"0699",
			x"0000" when x"069A",
			x"0000" when x"069B",
			x"0000" when x"069C",
			x"0000" when x"069D",
			x"0000" when x"069E",
			x"0000" when x"069F",
			x"0000" when x"06A0",
			x"0000" when x"06A1",
			x"0000" when x"06A2",
			x"0000" when x"06A3",
			x"0000" when x"06A4",
			x"0000" when x"06A5",
			x"0000" when x"06A6",
			x"0000" when x"06A7",
			x"0000" when x"06A8",
			x"0000" when x"06A9",
			x"0000" when x"06AA",
			x"0000" when x"06AB",
			x"0000" when x"06AC",
			x"0000" when x"06AD",
			x"0000" when x"06AE",
			x"0000" when x"06AF",
			x"0000" when x"06B0",
			x"0000" when x"06B1",
			x"0000" when x"06B2",
			x"0000" when x"06B3",
			x"0000" when x"06B4",
			x"0000" when x"06B5",
			x"0000" when x"06B6",
			x"0000" when x"06B7",
			x"0000" when x"06B8",
			x"0000" when x"06B9",
			x"0000" when x"06BA",
			x"0000" when x"06BB",
			x"0000" when x"06BC",
			x"0000" when x"06BD",
			x"0000" when x"06BE",
			x"0000" when x"06BF",
			x"0000" when x"06C0",
			x"0000" when x"06C1",
			x"0000" when x"06C2",
			x"0000" when x"06C3",
			x"0000" when x"06C4",
			x"0000" when x"06C5",
			x"0000" when x"06C6",
			x"0000" when x"06C7",
			x"0000" when x"06C8",
			x"0000" when x"06C9",
			x"0000" when x"06CA",
			x"0000" when x"06CB",
			x"0000" when x"06CC",
			x"0000" when x"06CD",
			x"0000" when x"06CE",
			x"0000" when x"06CF",
			x"0000" when x"06D0",
			x"0000" when x"06D1",
			x"0000" when x"06D2",
			x"0000" when x"06D3",
			x"0000" when x"06D4",
			x"0000" when x"06D5",
			x"0000" when x"06D6",
			x"0000" when x"06D7",
			x"0000" when x"06D8",
			x"0000" when x"06D9",
			x"0000" when x"06DA",
			x"0000" when x"06DB",
			x"0000" when x"06DC",
			x"0000" when x"06DD",
			x"0000" when x"06DE",
			x"0000" when x"06DF",
			x"0000" when x"06E0",
			x"0000" when x"06E1",
			x"0000" when x"06E2",
			x"0000" when x"06E3",
			x"0000" when x"06E4",
			x"0000" when x"06E5",
			x"0000" when x"06E6",
			x"0000" when x"06E7",
			x"0000" when x"06E8",
			x"0000" when x"06E9",
			x"0000" when x"06EA",
			x"0000" when x"06EB",
			x"0000" when x"06EC",
			x"0000" when x"06ED",
			x"0000" when x"06EE",
			x"0000" when x"06EF",
			x"0000" when x"06F0",
			x"0000" when x"06F1",
			x"0000" when x"06F2",
			x"0000" when x"06F3",
			x"0000" when x"06F4",
			x"0000" when x"06F5",
			x"0000" when x"06F6",
			x"0000" when x"06F7",
			x"0000" when x"06F8",
			x"0000" when x"06F9",
			x"0000" when x"06FA",
			x"0000" when x"06FB",
			x"0000" when x"06FC",
			x"0000" when x"06FD",
			x"0000" when x"06FE",
			x"0000" when x"06FF",
			x"0000" when x"0700",
			x"0000" when x"0701",
			x"0000" when x"0702",
			x"0000" when x"0703",
			x"0000" when x"0704",
			x"0000" when x"0705",
			x"0000" when x"0706",
			x"0000" when x"0707",
			x"0000" when x"0708",
			x"0000" when x"0709",
			x"0000" when x"070A",
			x"0000" when x"070B",
			x"0000" when x"070C",
			x"0000" when x"070D",
			x"0000" when x"070E",
			x"0000" when x"070F",
			x"0000" when x"0710",
			x"0000" when x"0711",
			x"0000" when x"0712",
			x"0000" when x"0713",
			x"0000" when x"0714",
			x"0000" when x"0715",
			x"0000" when x"0716",
			x"0000" when x"0717",
			x"0000" when x"0718",
			x"0000" when x"0719",
			x"0000" when x"071A",
			x"0000" when x"071B",
			x"0000" when x"071C",
			x"0000" when x"071D",
			x"0000" when x"071E",
			x"0000" when x"071F",
			x"0000" when x"0720",
			x"0000" when x"0721",
			x"0000" when x"0722",
			x"0000" when x"0723",
			x"0000" when x"0724",
			x"0000" when x"0725",
			x"0000" when x"0726",
			x"0000" when x"0727",
			x"0000" when x"0728",
			x"0000" when x"0729",
			x"0000" when x"072A",
			x"0000" when x"072B",
			x"0000" when x"072C",
			x"0000" when x"072D",
			x"0000" when x"072E",
			x"0000" when x"072F",
			x"0000" when x"0730",
			x"0000" when x"0731",
			x"0000" when x"0732",
			x"0000" when x"0733",
			x"0000" when x"0734",
			x"0000" when x"0735",
			x"0000" when x"0736",
			x"0000" when x"0737",
			x"0000" when x"0738",
			x"0000" when x"0739",
			x"0000" when x"073A",
			x"0000" when x"073B",
			x"0000" when x"073C",
			x"0000" when x"073D",
			x"0000" when x"073E",
			x"0000" when x"073F",
			x"0000" when x"0740",
			x"0000" when x"0741",
			x"0000" when x"0742",
			x"0000" when x"0743",
			x"0000" when x"0744",
			x"0000" when x"0745",
			x"0000" when x"0746",
			x"0000" when x"0747",
			x"0000" when x"0748",
			x"0000" when x"0749",
			x"0000" when x"074A",
			x"0000" when x"074B",
			x"0000" when x"074C",
			x"0000" when x"074D",
			x"0000" when x"074E",
			x"0000" when x"074F",
			x"0000" when x"0750",
			x"0000" when x"0751",
			x"0000" when x"0752",
			x"0000" when x"0753",
			x"0000" when x"0754",
			x"0000" when x"0755",
			x"0000" when x"0756",
			x"0000" when x"0757",
			x"0000" when x"0758",
			x"0000" when x"0759",
			x"0000" when x"075A",
			x"0000" when x"075B",
			x"0000" when x"075C",
			x"0000" when x"075D",
			x"0000" when x"075E",
			x"0000" when x"075F",
			x"0000" when x"0760",
			x"0000" when x"0761",
			x"0000" when x"0762",
			x"0000" when x"0763",
			x"0000" when x"0764",
			x"0000" when x"0765",
			x"0000" when x"0766",
			x"0000" when x"0767",
			x"0000" when x"0768",
			x"0000" when x"0769",
			x"0000" when x"076A",
			x"0000" when x"076B",
			x"0000" when x"076C",
			x"0000" when x"076D",
			x"0000" when x"076E",
			x"0000" when x"076F",
			x"0000" when x"0770",
			x"0000" when x"0771",
			x"0000" when x"0772",
			x"0000" when x"0773",
			x"0000" when x"0774",
			x"0000" when x"0775",
			x"0000" when x"0776",
			x"0000" when x"0777",
			x"0000" when x"0778",
			x"0000" when x"0779",
			x"0000" when x"077A",
			x"0000" when x"077B",
			x"0000" when x"077C",
			x"0000" when x"077D",
			x"0000" when x"077E",
			x"0000" when x"077F",
			x"0000" when x"0780",
			x"0000" when x"0781",
			x"0000" when x"0782",
			x"0000" when x"0783",
			x"0000" when x"0784",
			x"0000" when x"0785",
			x"0000" when x"0786",
			x"0000" when x"0787",
			x"0000" when x"0788",
			x"0000" when x"0789",
			x"0000" when x"078A",
			x"0000" when x"078B",
			x"0000" when x"078C",
			x"0000" when x"078D",
			x"0000" when x"078E",
			x"0000" when x"078F",
			x"0000" when x"0790",
			x"0000" when x"0791",
			x"0000" when x"0792",
			x"0000" when x"0793",
			x"0000" when x"0794",
			x"0000" when x"0795",
			x"0000" when x"0796",
			x"0000" when x"0797",
			x"0000" when x"0798",
			x"0000" when x"0799",
			x"0000" when x"079A",
			x"0000" when x"079B",
			x"0000" when x"079C",
			x"0000" when x"079D",
			x"0000" when x"079E",
			x"0000" when x"079F",
			x"0000" when x"07A0",
			x"0000" when x"07A1",
			x"0000" when x"07A2",
			x"0000" when x"07A3",
			x"0000" when x"07A4",
			x"0000" when x"07A5",
			x"0000" when x"07A6",
			x"0000" when x"07A7",
			x"0000" when x"07A8",
			x"0000" when x"07A9",
			x"0000" when x"07AA",
			x"0000" when x"07AB",
			x"0000" when x"07AC",
			x"0000" when x"07AD",
			x"0000" when x"07AE",
			x"0000" when x"07AF",
			x"0000" when x"07B0",
			x"0000" when x"07B1",
			x"0000" when x"07B2",
			x"0000" when x"07B3",
			x"0000" when x"07B4",
			x"0000" when x"07B5",
			x"0000" when x"07B6",
			x"0000" when x"07B7",
			x"0000" when x"07B8",
			x"0000" when x"07B9",
			x"0000" when x"07BA",
			x"0000" when x"07BB",
			x"0000" when x"07BC",
			x"0000" when x"07BD",
			x"0000" when x"07BE",
			x"0000" when x"07BF",
			x"0000" when x"07C0",
			x"0000" when x"07C1",
			x"0000" when x"07C2",
			x"0000" when x"07C3",
			x"0000" when x"07C4",
			x"0000" when x"07C5",
			x"0000" when x"07C6",
			x"0000" when x"07C7",
			x"0000" when x"07C8",
			x"0000" when x"07C9",
			x"0000" when x"07CA",
			x"0000" when x"07CB",
			x"0000" when x"07CC",
			x"0000" when x"07CD",
			x"0000" when x"07CE",
			x"0000" when x"07CF",
			x"0000" when x"07D0",
			x"0000" when x"07D1",
			x"0000" when x"07D2",
			x"0000" when x"07D3",
			x"0000" when x"07D4",
			x"0000" when x"07D5",
			x"0000" when x"07D6",
			x"0000" when x"07D7",
			x"0000" when x"07D8",
			x"0000" when x"07D9",
			x"0000" when x"07DA",
			x"0000" when x"07DB",
			x"0000" when x"07DC",
			x"0000" when x"07DD",
			x"0000" when x"07DE",
			x"0000" when x"07DF",
			x"0000" when x"07E0",
			x"0000" when x"07E1",
			x"0000" when x"07E2",
			x"0000" when x"07E3",
			x"0000" when x"07E4",
			x"0000" when x"07E5",
			x"0000" when x"07E6",
			x"0000" when x"07E7",
			x"0000" when x"07E8",
			x"0000" when x"07E9",
			x"0000" when x"07EA",
			x"0000" when x"07EB",
			x"0000" when x"07EC",
			x"0000" when x"07ED",
			x"0000" when x"07EE",
			x"0000" when x"07EF",
			x"0000" when x"07F0",
			x"0000" when x"07F1",
			x"0000" when x"07F2",
			x"0000" when x"07F3",
			x"0000" when x"07F4",
			x"0000" when x"07F5",
			x"0000" when x"07F6",
			x"0000" when x"07F7",
			x"0000" when x"07F8",
			x"0000" when x"07F9",
			x"0000" when x"07FA",
			x"0000" when x"07FB",
			x"0000" when x"07FC",
			x"0000" when x"07FD",
			x"0000" when x"07FE",
			x"0000" when x"07FF",
			x"0000" when x"0800",
			x"0000" when x"0801",
			x"0000" when x"0802",
			x"0000" when x"0803",
			x"0000" when x"0804",
			x"0000" when x"0805",
			x"0000" when x"0806",
			x"0000" when x"0807",
			x"0000" when x"0808",
			x"0000" when x"0809",
			x"0000" when x"080A",
			x"0000" when x"080B",
			x"0000" when x"080C",
			x"0000" when x"080D",
			x"0000" when x"080E",
			x"0000" when x"080F",
			x"0000" when x"0810",
			x"0000" when x"0811",
			x"0000" when x"0812",
			x"0000" when x"0813",
			x"0000" when x"0814",
			x"0000" when x"0815",
			x"0000" when x"0816",
			x"0000" when x"0817",
			x"0000" when x"0818",
			x"0000" when x"0819",
			x"0000" when x"081A",
			x"0000" when x"081B",
			x"0000" when x"081C",
			x"0000" when x"081D",
			x"0000" when x"081E",
			x"0000" when x"081F",
			x"0000" when x"0820",
			x"0000" when x"0821",
			x"0000" when x"0822",
			x"0000" when x"0823",
			x"0000" when x"0824",
			x"0000" when x"0825",
			x"0000" when x"0826",
			x"0000" when x"0827",
			x"0000" when x"0828",
			x"0000" when x"0829",
			x"0000" when x"082A",
			x"0000" when x"082B",
			x"0000" when x"082C",
			x"0000" when x"082D",
			x"0000" when x"082E",
			x"0000" when x"082F",
			x"0000" when x"0830",
			x"0000" when x"0831",
			x"0000" when x"0832",
			x"0000" when x"0833",
			x"0000" when x"0834",
			x"0000" when x"0835",
			x"0000" when x"0836",
			x"0000" when x"0837",
			x"0000" when x"0838",
			x"0000" when x"0839",
			x"0000" when x"083A",
			x"0000" when x"083B",
			x"0000" when x"083C",
			x"0000" when x"083D",
			x"0000" when x"083E",
			x"0000" when x"083F",
			x"0000" when x"0840",
			x"0000" when x"0841",
			x"0000" when x"0842",
			x"0000" when x"0843",
			x"0000" when x"0844",
			x"0000" when x"0845",
			x"0000" when x"0846",
			x"0000" when x"0847",
			x"0000" when x"0848",
			x"0000" when x"0849",
			x"0000" when x"084A",
			x"0000" when x"084B",
			x"0000" when x"084C",
			x"0000" when x"084D",
			x"0000" when x"084E",
			x"0000" when x"084F",
			x"0000" when x"0850",
			x"0000" when x"0851",
			x"0000" when x"0852",
			x"0000" when x"0853",
			x"0000" when x"0854",
			x"0000" when x"0855",
			x"0000" when x"0856",
			x"0000" when x"0857",
			x"0000" when x"0858",
			x"0000" when x"0859",
			x"0000" when x"085A",
			x"0000" when x"085B",
			x"0000" when x"085C",
			x"0000" when x"085D",
			x"0000" when x"085E",
			x"0000" when x"085F",
			x"0000" when x"0860",
			x"0000" when x"0861",
			x"0000" when x"0862",
			x"0000" when x"0863",
			x"0000" when x"0864",
			x"0000" when x"0865",
			x"0000" when x"0866",
			x"0000" when x"0867",
			x"0000" when x"0868",
			x"0000" when x"0869",
			x"0000" when x"086A",
			x"0000" when x"086B",
			x"0000" when x"086C",
			x"0000" when x"086D",
			x"0000" when x"086E",
			x"0000" when x"086F",
			x"0000" when x"0870",
			x"0000" when x"0871",
			x"0000" when x"0872",
			x"0000" when x"0873",
			x"0000" when x"0874",
			x"0000" when x"0875",
			x"0000" when x"0876",
			x"0000" when x"0877",
			x"0000" when x"0878",
			x"0000" when x"0879",
			x"0000" when x"087A",
			x"0000" when x"087B",
			x"0000" when x"087C",
			x"0000" when x"087D",
			x"0000" when x"087E",
			x"0000" when x"087F",
			x"0000" when x"0880",
			x"0000" when x"0881",
			x"0000" when x"0882",
			x"0000" when x"0883",
			x"0000" when x"0884",
			x"0000" when x"0885",
			x"0000" when x"0886",
			x"0000" when x"0887",
			x"0000" when x"0888",
			x"0000" when x"0889",
			x"0000" when x"088A",
			x"0000" when x"088B",
			x"0000" when x"088C",
			x"0000" when x"088D",
			x"0000" when x"088E",
			x"0000" when x"088F",
			x"0000" when x"0890",
			x"0000" when x"0891",
			x"0000" when x"0892",
			x"0000" when x"0893",
			x"0000" when x"0894",
			x"0000" when x"0895",
			x"0000" when x"0896",
			x"0000" when x"0897",
			x"0000" when x"0898",
			x"0000" when x"0899",
			x"0000" when x"089A",
			x"0000" when x"089B",
			x"0000" when x"089C",
			x"0000" when x"089D",
			x"0000" when x"089E",
			x"0000" when x"089F",
			x"0000" when x"08A0",
			x"0000" when x"08A1",
			x"0000" when x"08A2",
			x"0000" when x"08A3",
			x"0000" when x"08A4",
			x"0000" when x"08A5",
			x"0000" when x"08A6",
			x"0000" when x"08A7",
			x"0000" when x"08A8",
			x"0000" when x"08A9",
			x"0000" when x"08AA",
			x"0000" when x"08AB",
			x"0000" when x"08AC",
			x"0000" when x"08AD",
			x"0000" when x"08AE",
			x"0000" when x"08AF",
			x"0000" when x"08B0",
			x"0000" when x"08B1",
			x"0000" when x"08B2",
			x"0000" when x"08B3",
			x"0000" when x"08B4",
			x"0000" when x"08B5",
			x"0000" when x"08B6",
			x"0000" when x"08B7",
			x"0000" when x"08B8",
			x"0000" when x"08B9",
			x"0000" when x"08BA",
			x"0000" when x"08BB",
			x"0000" when x"08BC",
			x"0000" when x"08BD",
			x"0000" when x"08BE",
			x"0000" when x"08BF",
			x"0000" when x"08C0",
			x"0000" when x"08C1",
			x"0000" when x"08C2",
			x"0000" when x"08C3",
			x"0000" when x"08C4",
			x"0000" when x"08C5",
			x"0000" when x"08C6",
			x"0000" when x"08C7",
			x"0000" when x"08C8",
			x"0000" when x"08C9",
			x"0000" when x"08CA",
			x"0000" when x"08CB",
			x"0000" when x"08CC",
			x"0000" when x"08CD",
			x"0000" when x"08CE",
			x"0000" when x"08CF",
			x"0000" when x"08D0",
			x"0000" when x"08D1",
			x"0000" when x"08D2",
			x"0000" when x"08D3",
			x"0000" when x"08D4",
			x"0000" when x"08D5",
			x"0000" when x"08D6",
			x"0000" when x"08D7",
			x"0000" when x"08D8",
			x"0000" when x"08D9",
			x"0000" when x"08DA",
			x"0000" when x"08DB",
			x"0000" when x"08DC",
			x"0000" when x"08DD",
			x"0000" when x"08DE",
			x"0000" when x"08DF",
			x"0000" when x"08E0",
			x"0000" when x"08E1",
			x"0000" when x"08E2",
			x"0000" when x"08E3",
			x"0000" when x"08E4",
			x"0000" when x"08E5",
			x"0000" when x"08E6",
			x"0000" when x"08E7",
			x"0000" when x"08E8",
			x"0000" when x"08E9",
			x"0000" when x"08EA",
			x"0000" when x"08EB",
			x"0000" when x"08EC",
			x"0000" when x"08ED",
			x"0000" when x"08EE",
			x"0000" when x"08EF",
			x"0000" when x"08F0",
			x"0000" when x"08F1",
			x"0000" when x"08F2",
			x"0000" when x"08F3",
			x"0000" when x"08F4",
			x"0000" when x"08F5",
			x"0000" when x"08F6",
			x"0000" when x"08F7",
			x"0000" when x"08F8",
			x"0000" when x"08F9",
			x"0000" when x"08FA",
			x"0000" when x"08FB",
			x"0000" when x"08FC",
			x"0000" when x"08FD",
			x"0000" when x"08FE",
			x"0000" when x"08FF",
			x"0000" when x"0900",
			x"0000" when x"0901",
			x"0000" when x"0902",
			x"0000" when x"0903",
			x"0000" when x"0904",
			x"0000" when x"0905",
			x"0000" when x"0906",
			x"0000" when x"0907",
			x"0000" when x"0908",
			x"0000" when x"0909",
			x"0000" when x"090A",
			x"0000" when x"090B",
			x"0000" when x"090C",
			x"0000" when x"090D",
			x"0000" when x"090E",
			x"0000" when x"090F",
			x"0000" when x"0910",
			x"0000" when x"0911",
			x"0000" when x"0912",
			x"0000" when x"0913",
			x"0000" when x"0914",
			x"0000" when x"0915",
			x"0000" when x"0916",
			x"0000" when x"0917",
			x"0000" when x"0918",
			x"0000" when x"0919",
			x"0000" when x"091A",
			x"0000" when x"091B",
			x"0000" when x"091C",
			x"0000" when x"091D",
			x"0000" when x"091E",
			x"0000" when x"091F",
			x"0000" when x"0920",
			x"0000" when x"0921",
			x"0000" when x"0922",
			x"0000" when x"0923",
			x"0000" when x"0924",
			x"0000" when x"0925",
			x"0000" when x"0926",
			x"0000" when x"0927",
			x"0000" when x"0928",
			x"0000" when x"0929",
			x"0000" when x"092A",
			x"0000" when x"092B",
			x"0000" when x"092C",
			x"0000" when x"092D",
			x"0000" when x"092E",
			x"0000" when x"092F",
			x"0000" when x"0930",
			x"0000" when x"0931",
			x"0000" when x"0932",
			x"0000" when x"0933",
			x"0000" when x"0934",
			x"0000" when x"0935",
			x"0000" when x"0936",
			x"0000" when x"0937",
			x"0000" when x"0938",
			x"0000" when x"0939",
			x"0000" when x"093A",
			x"0000" when x"093B",
			x"0000" when x"093C",
			x"0000" when x"093D",
			x"0000" when x"093E",
			x"0000" when x"093F",
			x"0000" when x"0940",
			x"0000" when x"0941",
			x"0000" when x"0942",
			x"0000" when x"0943",
			x"0000" when x"0944",
			x"0000" when x"0945",
			x"0000" when x"0946",
			x"0000" when x"0947",
			x"0000" when x"0948",
			x"0000" when x"0949",
			x"0000" when x"094A",
			x"0000" when x"094B",
			x"0000" when x"094C",
			x"0000" when x"094D",
			x"0000" when x"094E",
			x"0000" when x"094F",
			x"0000" when x"0950",
			x"0000" when x"0951",
			x"0000" when x"0952",
			x"0000" when x"0953",
			x"0000" when x"0954",
			x"0000" when x"0955",
			x"0000" when x"0956",
			x"0000" when x"0957",
			x"0000" when x"0958",
			x"0000" when x"0959",
			x"0000" when x"095A",
			x"0000" when x"095B",
			x"0000" when x"095C",
			x"0000" when x"095D",
			x"0000" when x"095E",
			x"0000" when x"095F",
			x"0000" when x"0960",
			x"0000" when x"0961",
			x"0000" when x"0962",
			x"0000" when x"0963",
			x"0000" when x"0964",
			x"0000" when x"0965",
			x"0000" when x"0966",
			x"0000" when x"0967",
			x"0000" when x"0968",
			x"0000" when x"0969",
			x"0000" when x"096A",
			x"0000" when x"096B",
			x"0000" when x"096C",
			x"0000" when x"096D",
			x"0000" when x"096E",
			x"0000" when x"096F",
			x"0000" when x"0970",
			x"0000" when x"0971",
			x"0000" when x"0972",
			x"0000" when x"0973",
			x"0000" when x"0974",
			x"0000" when x"0975",
			x"0000" when x"0976",
			x"0000" when x"0977",
			x"0000" when x"0978",
			x"0000" when x"0979",
			x"0000" when x"097A",
			x"0000" when x"097B",
			x"0000" when x"097C",
			x"0000" when x"097D",
			x"0000" when x"097E",
			x"0000" when x"097F",
			x"0000" when x"0980",
			x"0000" when x"0981",
			x"0000" when x"0982",
			x"0000" when x"0983",
			x"0000" when x"0984",
			x"0000" when x"0985",
			x"0000" when x"0986",
			x"0000" when x"0987",
			x"0000" when x"0988",
			x"0000" when x"0989",
			x"0000" when x"098A",
			x"0000" when x"098B",
			x"0000" when x"098C",
			x"0000" when x"098D",
			x"0000" when x"098E",
			x"0000" when x"098F",
			x"0000" when x"0990",
			x"0000" when x"0991",
			x"0000" when x"0992",
			x"0000" when x"0993",
			x"0000" when x"0994",
			x"0000" when x"0995",
			x"0000" when x"0996",
			x"0000" when x"0997",
			x"0000" when x"0998",
			x"0000" when x"0999",
			x"0000" when x"099A",
			x"0000" when x"099B",
			x"0000" when x"099C",
			x"0000" when x"099D",
			x"0000" when x"099E",
			x"0000" when x"099F",
			x"0000" when x"09A0",
			x"0000" when x"09A1",
			x"0000" when x"09A2",
			x"0000" when x"09A3",
			x"0000" when x"09A4",
			x"0000" when x"09A5",
			x"0000" when x"09A6",
			x"0000" when x"09A7",
			x"0000" when x"09A8",
			x"0000" when x"09A9",
			x"0000" when x"09AA",
			x"0000" when x"09AB",
			x"0000" when x"09AC",
			x"0000" when x"09AD",
			x"0000" when x"09AE",
			x"0000" when x"09AF",
			x"0000" when x"09B0",
			x"0000" when x"09B1",
			x"0000" when x"09B2",
			x"0000" when x"09B3",
			x"0000" when x"09B4",
			x"0000" when x"09B5",
			x"0000" when x"09B6",
			x"0000" when x"09B7",
			x"0000" when x"09B8",
			x"0000" when x"09B9",
			x"0000" when x"09BA",
			x"0000" when x"09BB",
			x"0000" when x"09BC",
			x"0000" when x"09BD",
			x"0000" when x"09BE",
			x"0000" when x"09BF",
			x"0000" when x"09C0",
			x"0000" when x"09C1",
			x"0000" when x"09C2",
			x"0000" when x"09C3",
			x"0000" when x"09C4",
			x"0000" when x"09C5",
			x"0000" when x"09C6",
			x"0000" when x"09C7",
			x"0000" when x"09C8",
			x"0000" when x"09C9",
			x"0000" when x"09CA",
			x"0000" when x"09CB",
			x"0000" when x"09CC",
			x"0000" when x"09CD",
			x"0000" when x"09CE",
			x"0000" when x"09CF",
			x"0000" when x"09D0",
			x"0000" when x"09D1",
			x"0000" when x"09D2",
			x"0000" when x"09D3",
			x"0000" when x"09D4",
			x"0000" when x"09D5",
			x"0000" when x"09D6",
			x"0000" when x"09D7",
			x"0000" when x"09D8",
			x"0000" when x"09D9",
			x"0000" when x"09DA",
			x"0000" when x"09DB",
			x"0000" when x"09DC",
			x"0000" when x"09DD",
			x"0000" when x"09DE",
			x"0000" when x"09DF",
			x"0000" when x"09E0",
			x"0000" when x"09E1",
			x"0000" when x"09E2",
			x"0000" when x"09E3",
			x"0000" when x"09E4",
			x"0000" when x"09E5",
			x"0000" when x"09E6",
			x"0000" when x"09E7",
			x"0000" when x"09E8",
			x"0000" when x"09E9",
			x"0000" when x"09EA",
			x"0000" when x"09EB",
			x"0000" when x"09EC",
			x"0000" when x"09ED",
			x"0000" when x"09EE",
			x"0000" when x"09EF",
			x"0000" when x"09F0",
			x"0000" when x"09F1",
			x"0000" when x"09F2",
			x"0000" when x"09F3",
			x"0000" when x"09F4",
			x"0000" when x"09F5",
			x"0000" when x"09F6",
			x"0000" when x"09F7",
			x"0000" when x"09F8",
			x"0000" when x"09F9",
			x"0000" when x"09FA",
			x"0000" when x"09FB",
			x"0000" when x"09FC",
			x"0000" when x"09FD",
			x"0000" when x"09FE",
			x"0000" when x"09FF",
			x"0000" when x"0A00",
			x"0000" when x"0A01",
			x"0000" when x"0A02",
			x"0000" when x"0A03",
			x"0000" when x"0A04",
			x"0000" when x"0A05",
			x"0000" when x"0A06",
			x"0000" when x"0A07",
			x"0000" when x"0A08",
			x"0000" when x"0A09",
			x"0000" when x"0A0A",
			x"0000" when x"0A0B",
			x"0000" when x"0A0C",
			x"0000" when x"0A0D",
			x"0000" when x"0A0E",
			x"0000" when x"0A0F",
			x"0000" when x"0A10",
			x"0000" when x"0A11",
			x"0000" when x"0A12",
			x"0000" when x"0A13",
			x"0000" when x"0A14",
			x"0000" when x"0A15",
			x"0000" when x"0A16",
			x"0000" when x"0A17",
			x"0000" when x"0A18",
			x"0000" when x"0A19",
			x"0000" when x"0A1A",
			x"0000" when x"0A1B",
			x"0000" when x"0A1C",
			x"0000" when x"0A1D",
			x"0000" when x"0A1E",
			x"0000" when x"0A1F",
			x"0000" when x"0A20",
			x"0000" when x"0A21",
			x"0000" when x"0A22",
			x"0000" when x"0A23",
			x"0000" when x"0A24",
			x"0000" when x"0A25",
			x"0000" when x"0A26",
			x"0000" when x"0A27",
			x"0000" when x"0A28",
			x"0000" when x"0A29",
			x"0000" when x"0A2A",
			x"0000" when x"0A2B",
			x"0000" when x"0A2C",
			x"0000" when x"0A2D",
			x"0000" when x"0A2E",
			x"0000" when x"0A2F",
			x"0000" when x"0A30",
			x"0000" when x"0A31",
			x"0000" when x"0A32",
			x"0000" when x"0A33",
			x"0000" when x"0A34",
			x"0000" when x"0A35",
			x"0000" when x"0A36",
			x"0000" when x"0A37",
			x"0000" when x"0A38",
			x"0000" when x"0A39",
			x"0000" when x"0A3A",
			x"0000" when x"0A3B",
			x"0000" when x"0A3C",
			x"0000" when x"0A3D",
			x"0000" when x"0A3E",
			x"0000" when x"0A3F",
			x"0000" when x"0A40",
			x"0000" when x"0A41",
			x"0000" when x"0A42",
			x"0000" when x"0A43",
			x"0000" when x"0A44",
			x"0000" when x"0A45",
			x"0000" when x"0A46",
			x"0000" when x"0A47",
			x"0000" when x"0A48",
			x"0000" when x"0A49",
			x"0000" when x"0A4A",
			x"0000" when x"0A4B",
			x"0000" when x"0A4C",
			x"0000" when x"0A4D",
			x"0000" when x"0A4E",
			x"0000" when x"0A4F",
			x"0000" when x"0A50",
			x"0000" when x"0A51",
			x"0000" when x"0A52",
			x"0000" when x"0A53",
			x"0000" when x"0A54",
			x"0000" when x"0A55",
			x"0000" when x"0A56",
			x"0000" when x"0A57",
			x"0000" when x"0A58",
			x"0000" when x"0A59",
			x"0000" when x"0A5A",
			x"0000" when x"0A5B",
			x"0000" when x"0A5C",
			x"0000" when x"0A5D",
			x"0000" when x"0A5E",
			x"0000" when x"0A5F",
			x"0000" when x"0A60",
			x"0000" when x"0A61",
			x"0000" when x"0A62",
			x"0000" when x"0A63",
			x"0000" when x"0A64",
			x"0000" when x"0A65",
			x"0000" when x"0A66",
			x"0000" when x"0A67",
			x"0000" when x"0A68",
			x"0000" when x"0A69",
			x"0000" when x"0A6A",
			x"0000" when x"0A6B",
			x"0000" when x"0A6C",
			x"0000" when x"0A6D",
			x"0000" when x"0A6E",
			x"0000" when x"0A6F",
			x"0000" when x"0A70",
			x"0000" when x"0A71",
			x"0000" when x"0A72",
			x"0000" when x"0A73",
			x"0000" when x"0A74",
			x"0000" when x"0A75",
			x"0000" when x"0A76",
			x"0000" when x"0A77",
			x"0000" when x"0A78",
			x"0000" when x"0A79",
			x"0000" when x"0A7A",
			x"0000" when x"0A7B",
			x"0000" when x"0A7C",
			x"0000" when x"0A7D",
			x"0000" when x"0A7E",
			x"0000" when x"0A7F",
			x"0000" when x"0A80",
			x"0000" when x"0A81",
			x"0000" when x"0A82",
			x"0000" when x"0A83",
			x"0000" when x"0A84",
			x"0000" when x"0A85",
			x"0000" when x"0A86",
			x"0000" when x"0A87",
			x"0000" when x"0A88",
			x"0000" when x"0A89",
			x"0000" when x"0A8A",
			x"0000" when x"0A8B",
			x"0000" when x"0A8C",
			x"0000" when x"0A8D",
			x"0000" when x"0A8E",
			x"0000" when x"0A8F",
			x"0000" when x"0A90",
			x"0000" when x"0A91",
			x"0000" when x"0A92",
			x"0000" when x"0A93",
			x"0000" when x"0A94",
			x"0000" when x"0A95",
			x"0000" when x"0A96",
			x"0000" when x"0A97",
			x"0000" when x"0A98",
			x"0000" when x"0A99",
			x"0000" when x"0A9A",
			x"0000" when x"0A9B",
			x"0000" when x"0A9C",
			x"0000" when x"0A9D",
			x"0000" when x"0A9E",
			x"0000" when x"0A9F",
			x"0000" when x"0AA0",
			x"0000" when x"0AA1",
			x"0000" when x"0AA2",
			x"0000" when x"0AA3",
			x"0000" when x"0AA4",
			x"0000" when x"0AA5",
			x"0000" when x"0AA6",
			x"0000" when x"0AA7",
			x"0000" when x"0AA8",
			x"0000" when x"0AA9",
			x"0000" when x"0AAA",
			x"0000" when x"0AAB",
			x"0000" when x"0AAC",
			x"0000" when x"0AAD",
			x"0000" when x"0AAE",
			x"0000" when x"0AAF",
			x"0000" when x"0AB0",
			x"0000" when x"0AB1",
			x"0000" when x"0AB2",
			x"0000" when x"0AB3",
			x"0000" when x"0AB4",
			x"0000" when x"0AB5",
			x"0000" when x"0AB6",
			x"0000" when x"0AB7",
			x"0000" when x"0AB8",
			x"0000" when x"0AB9",
			x"0000" when x"0ABA",
			x"0000" when x"0ABB",
			x"0000" when x"0ABC",
			x"0000" when x"0ABD",
			x"0000" when x"0ABE",
			x"0000" when x"0ABF",
			x"0000" when x"0AC0",
			x"0000" when x"0AC1",
			x"0000" when x"0AC2",
			x"0000" when x"0AC3",
			x"0000" when x"0AC4",
			x"0000" when x"0AC5",
			x"0000" when x"0AC6",
			x"0000" when x"0AC7",
			x"0000" when x"0AC8",
			x"0000" when x"0AC9",
			x"0000" when x"0ACA",
			x"0000" when x"0ACB",
			x"0000" when x"0ACC",
			x"0000" when x"0ACD",
			x"0000" when x"0ACE",
			x"0000" when x"0ACF",
			x"0000" when x"0AD0",
			x"0000" when x"0AD1",
			x"0000" when x"0AD2",
			x"0000" when x"0AD3",
			x"0000" when x"0AD4",
			x"0000" when x"0AD5",
			x"0000" when x"0AD6",
			x"0000" when x"0AD7",
			x"0000" when x"0AD8",
			x"0000" when x"0AD9",
			x"0000" when x"0ADA",
			x"0000" when x"0ADB",
			x"0000" when x"0ADC",
			x"0000" when x"0ADD",
			x"0000" when x"0ADE",
			x"0000" when x"0ADF",
			x"0000" when x"0AE0",
			x"0000" when x"0AE1",
			x"0000" when x"0AE2",
			x"0000" when x"0AE3",
			x"0000" when x"0AE4",
			x"0000" when x"0AE5",
			x"0000" when x"0AE6",
			x"0000" when x"0AE7",
			x"0000" when x"0AE8",
			x"0000" when x"0AE9",
			x"0000" when x"0AEA",
			x"0000" when x"0AEB",
			x"0000" when x"0AEC",
			x"0000" when x"0AED",
			x"0000" when x"0AEE",
			x"0000" when x"0AEF",
			x"0000" when x"0AF0",
			x"0000" when x"0AF1",
			x"0000" when x"0AF2",
			x"0000" when x"0AF3",
			x"0000" when x"0AF4",
			x"0000" when x"0AF5",
			x"0000" when x"0AF6",
			x"0000" when x"0AF7",
			x"0000" when x"0AF8",
			x"0000" when x"0AF9",
			x"0000" when x"0AFA",
			x"0000" when x"0AFB",
			x"0000" when x"0AFC",
			x"0000" when x"0AFD",
			x"0000" when x"0AFE",
			x"0000" when x"0AFF",
			x"0000" when x"0B00",
			x"0000" when x"0B01",
			x"0000" when x"0B02",
			x"0000" when x"0B03",
			x"0000" when x"0B04",
			x"0000" when x"0B05",
			x"0000" when x"0B06",
			x"0000" when x"0B07",
			x"0000" when x"0B08",
			x"0000" when x"0B09",
			x"0000" when x"0B0A",
			x"0000" when x"0B0B",
			x"0000" when x"0B0C",
			x"0000" when x"0B0D",
			x"0000" when x"0B0E",
			x"0000" when x"0B0F",
			x"0000" when x"0B10",
			x"0000" when x"0B11",
			x"0000" when x"0B12",
			x"0000" when x"0B13",
			x"0000" when x"0B14",
			x"0000" when x"0B15",
			x"0000" when x"0B16",
			x"0000" when x"0B17",
			x"0000" when x"0B18",
			x"0000" when x"0B19",
			x"0000" when x"0B1A",
			x"0000" when x"0B1B",
			x"0000" when x"0B1C",
			x"0000" when x"0B1D",
			x"0000" when x"0B1E",
			x"0000" when x"0B1F",
			x"0000" when x"0B20",
			x"0000" when x"0B21",
			x"0000" when x"0B22",
			x"0000" when x"0B23",
			x"0000" when x"0B24",
			x"0000" when x"0B25",
			x"0000" when x"0B26",
			x"0000" when x"0B27",
			x"0000" when x"0B28",
			x"0000" when x"0B29",
			x"0000" when x"0B2A",
			x"0000" when x"0B2B",
			x"0000" when x"0B2C",
			x"0000" when x"0B2D",
			x"0000" when x"0B2E",
			x"0000" when x"0B2F",
			x"0000" when x"0B30",
			x"0000" when x"0B31",
			x"0000" when x"0B32",
			x"0000" when x"0B33",
			x"0000" when x"0B34",
			x"0000" when x"0B35",
			x"0000" when x"0B36",
			x"0000" when x"0B37",
			x"0000" when x"0B38",
			x"0000" when x"0B39",
			x"0000" when x"0B3A",
			x"0000" when x"0B3B",
			x"0000" when x"0B3C",
			x"0000" when x"0B3D",
			x"0000" when x"0B3E",
			x"0000" when x"0B3F",
			x"0000" when x"0B40",
			x"0000" when x"0B41",
			x"0000" when x"0B42",
			x"0000" when x"0B43",
			x"0000" when x"0B44",
			x"0000" when x"0B45",
			x"0000" when x"0B46",
			x"0000" when x"0B47",
			x"0000" when x"0B48",
			x"0000" when x"0B49",
			x"0000" when x"0B4A",
			x"0000" when x"0B4B",
			x"0000" when x"0B4C",
			x"0000" when x"0B4D",
			x"0000" when x"0B4E",
			x"0000" when x"0B4F",
			x"0000" when x"0B50",
			x"0000" when x"0B51",
			x"0000" when x"0B52",
			x"0000" when x"0B53",
			x"0000" when x"0B54",
			x"0000" when x"0B55",
			x"0000" when x"0B56",
			x"0000" when x"0B57",
			x"0000" when x"0B58",
			x"0000" when x"0B59",
			x"0000" when x"0B5A",
			x"0000" when x"0B5B",
			x"0000" when x"0B5C",
			x"0000" when x"0B5D",
			x"0000" when x"0B5E",
			x"0000" when x"0B5F",
			x"0000" when x"0B60",
			x"0000" when x"0B61",
			x"0000" when x"0B62",
			x"0000" when x"0B63",
			x"0000" when x"0B64",
			x"0000" when x"0B65",
			x"0000" when x"0B66",
			x"0000" when x"0B67",
			x"0000" when x"0B68",
			x"0000" when x"0B69",
			x"0000" when x"0B6A",
			x"0000" when x"0B6B",
			x"0000" when x"0B6C",
			x"0000" when x"0B6D",
			x"0000" when x"0B6E",
			x"0000" when x"0B6F",
			x"0000" when x"0B70",
			x"0000" when x"0B71",
			x"0000" when x"0B72",
			x"0000" when x"0B73",
			x"0000" when x"0B74",
			x"0000" when x"0B75",
			x"0000" when x"0B76",
			x"0000" when x"0B77",
			x"0000" when x"0B78",
			x"0000" when x"0B79",
			x"0000" when x"0B7A",
			x"0000" when x"0B7B",
			x"0000" when x"0B7C",
			x"0000" when x"0B7D",
			x"0000" when x"0B7E",
			x"0000" when x"0B7F",
			x"0000" when x"0B80",
			x"0000" when x"0B81",
			x"0000" when x"0B82",
			x"0000" when x"0B83",
			x"0000" when x"0B84",
			x"0000" when x"0B85",
			x"0000" when x"0B86",
			x"0000" when x"0B87",
			x"0000" when x"0B88",
			x"0000" when x"0B89",
			x"0000" when x"0B8A",
			x"0000" when x"0B8B",
			x"0000" when x"0B8C",
			x"0000" when x"0B8D",
			x"0000" when x"0B8E",
			x"0000" when x"0B8F",
			x"0000" when x"0B90",
			x"0000" when x"0B91",
			x"0000" when x"0B92",
			x"0000" when x"0B93",
			x"0000" when x"0B94",
			x"0000" when x"0B95",
			x"0000" when x"0B96",
			x"0000" when x"0B97",
			x"0000" when x"0B98",
			x"0000" when x"0B99",
			x"0000" when x"0B9A",
			x"0000" when x"0B9B",
			x"0000" when x"0B9C",
			x"0000" when x"0B9D",
			x"0000" when x"0B9E",
			x"0000" when x"0B9F",
			x"0000" when x"0BA0",
			x"0000" when x"0BA1",
			x"0000" when x"0BA2",
			x"0000" when x"0BA3",
			x"0000" when x"0BA4",
			x"0000" when x"0BA5",
			x"0000" when x"0BA6",
			x"0000" when x"0BA7",
			x"0000" when x"0BA8",
			x"0000" when x"0BA9",
			x"0000" when x"0BAA",
			x"0000" when x"0BAB",
			x"0000" when x"0BAC",
			x"0000" when x"0BAD",
			x"0000" when x"0BAE",
			x"0000" when x"0BAF",
			x"0000" when x"0BB0",
			x"0000" when x"0BB1",
			x"0000" when x"0BB2",
			x"0000" when x"0BB3",
			x"0000" when x"0BB4",
			x"0000" when x"0BB5",
			x"0000" when x"0BB6",
			x"0000" when x"0BB7",
			x"0000" when x"0BB8",
			x"0000" when x"0BB9",
			x"0000" when x"0BBA",
			x"0000" when x"0BBB",
			x"0000" when x"0BBC",
			x"0000" when x"0BBD",
			x"0000" when x"0BBE",
			x"0000" when x"0BBF",
			x"0000" when x"0BC0",
			x"0000" when x"0BC1",
			x"0000" when x"0BC2",
			x"0000" when x"0BC3",
			x"0000" when x"0BC4",
			x"0000" when x"0BC5",
			x"0000" when x"0BC6",
			x"0000" when x"0BC7",
			x"0000" when x"0BC8",
			x"0000" when x"0BC9",
			x"0000" when x"0BCA",
			x"0000" when x"0BCB",
			x"0000" when x"0BCC",
			x"0000" when x"0BCD",
			x"0000" when x"0BCE",
			x"0000" when x"0BCF",
			x"0000" when x"0BD0",
			x"0000" when x"0BD1",
			x"0000" when x"0BD2",
			x"0000" when x"0BD3",
			x"0000" when x"0BD4",
			x"0000" when x"0BD5",
			x"0000" when x"0BD6",
			x"0000" when x"0BD7",
			x"0000" when x"0BD8",
			x"0000" when x"0BD9",
			x"0000" when x"0BDA",
			x"0000" when x"0BDB",
			x"0000" when x"0BDC",
			x"0000" when x"0BDD",
			x"0000" when x"0BDE",
			x"0000" when x"0BDF",
			x"0000" when x"0BE0",
			x"0000" when x"0BE1",
			x"0000" when x"0BE2",
			x"0000" when x"0BE3",
			x"0000" when x"0BE4",
			x"0000" when x"0BE5",
			x"0000" when x"0BE6",
			x"0000" when x"0BE7",
			x"0000" when x"0BE8",
			x"0000" when x"0BE9",
			x"0000" when x"0BEA",
			x"0000" when x"0BEB",
			x"0000" when x"0BEC",
			x"0000" when x"0BED",
			x"0000" when x"0BEE",
			x"0000" when x"0BEF",
			x"0000" when x"0BF0",
			x"0000" when x"0BF1",
			x"0000" when x"0BF2",
			x"0000" when x"0BF3",
			x"0000" when x"0BF4",
			x"0000" when x"0BF5",
			x"0000" when x"0BF6",
			x"0000" when x"0BF7",
			x"0000" when x"0BF8",
			x"0000" when x"0BF9",
			x"0000" when x"0BFA",
			x"0000" when x"0BFB",
			x"0000" when x"0BFC",
			x"0000" when x"0BFD",
			x"0000" when x"0BFE",
			x"0000" when x"0BFF",
			x"0000" when x"0C00",
			x"0000" when x"0C01",
			x"0000" when x"0C02",
			x"0000" when x"0C03",
			x"0000" when x"0C04",
			x"0000" when x"0C05",
			x"0000" when x"0C06",
			x"0000" when x"0C07",
			x"0000" when x"0C08",
			x"0000" when x"0C09",
			x"0000" when x"0C0A",
			x"0000" when x"0C0B",
			x"0000" when x"0C0C",
			x"0000" when x"0C0D",
			x"0000" when x"0C0E",
			x"0000" when x"0C0F",
			x"0000" when x"0C10",
			x"0000" when x"0C11",
			x"0000" when x"0C12",
			x"0000" when x"0C13",
			x"0000" when x"0C14",
			x"0000" when x"0C15",
			x"0000" when x"0C16",
			x"0000" when x"0C17",
			x"0000" when x"0C18",
			x"0000" when x"0C19",
			x"0000" when x"0C1A",
			x"0000" when x"0C1B",
			x"0000" when x"0C1C",
			x"0000" when x"0C1D",
			x"0000" when x"0C1E",
			x"0000" when x"0C1F",
			x"0000" when x"0C20",
			x"0000" when x"0C21",
			x"0000" when x"0C22",
			x"0000" when x"0C23",
			x"0000" when x"0C24",
			x"0000" when x"0C25",
			x"0000" when x"0C26",
			x"0000" when x"0C27",
			x"0000" when x"0C28",
			x"0000" when x"0C29",
			x"0000" when x"0C2A",
			x"0000" when x"0C2B",
			x"0000" when x"0C2C",
			x"0000" when x"0C2D",
			x"0000" when x"0C2E",
			x"0000" when x"0C2F",
			x"0000" when x"0C30",
			x"0000" when x"0C31",
			x"0000" when x"0C32",
			x"0000" when x"0C33",
			x"0000" when x"0C34",
			x"0000" when x"0C35",
			x"0000" when x"0C36",
			x"0000" when x"0C37",
			x"0000" when x"0C38",
			x"0000" when x"0C39",
			x"0000" when x"0C3A",
			x"0000" when x"0C3B",
			x"0000" when x"0C3C",
			x"0000" when x"0C3D",
			x"0000" when x"0C3E",
			x"0000" when x"0C3F",
			x"0000" when x"0C40",
			x"0000" when x"0C41",
			x"0000" when x"0C42",
			x"0000" when x"0C43",
			x"0000" when x"0C44",
			x"0000" when x"0C45",
			x"0000" when x"0C46",
			x"0000" when x"0C47",
			x"0000" when x"0C48",
			x"0000" when x"0C49",
			x"0000" when x"0C4A",
			x"0000" when x"0C4B",
			x"0000" when x"0C4C",
			x"0000" when x"0C4D",
			x"0000" when x"0C4E",
			x"0000" when x"0C4F",
			x"0000" when x"0C50",
			x"0000" when x"0C51",
			x"0000" when x"0C52",
			x"0000" when x"0C53",
			x"0000" when x"0C54",
			x"0000" when x"0C55",
			x"0000" when x"0C56",
			x"0000" when x"0C57",
			x"0000" when x"0C58",
			x"0000" when x"0C59",
			x"0000" when x"0C5A",
			x"0000" when x"0C5B",
			x"0000" when x"0C5C",
			x"0000" when x"0C5D",
			x"0000" when x"0C5E",
			x"0000" when x"0C5F",
			x"0000" when x"0C60",
			x"0000" when x"0C61",
			x"0000" when x"0C62",
			x"0000" when x"0C63",
			x"0000" when x"0C64",
			x"0000" when x"0C65",
			x"0000" when x"0C66",
			x"0000" when x"0C67",
			x"0000" when x"0C68",
			x"0000" when x"0C69",
			x"0000" when x"0C6A",
			x"0000" when x"0C6B",
			x"0000" when x"0C6C",
			x"0000" when x"0C6D",
			x"0000" when x"0C6E",
			x"0000" when x"0C6F",
			x"0000" when x"0C70",
			x"0000" when x"0C71",
			x"0000" when x"0C72",
			x"0000" when x"0C73",
			x"0000" when x"0C74",
			x"0000" when x"0C75",
			x"0000" when x"0C76",
			x"0000" when x"0C77",
			x"0000" when x"0C78",
			x"0000" when x"0C79",
			x"0000" when x"0C7A",
			x"0000" when x"0C7B",
			x"0000" when x"0C7C",
			x"0000" when x"0C7D",
			x"0000" when x"0C7E",
			x"0000" when x"0C7F",
			x"0000" when x"0C80",
			x"0000" when x"0C81",
			x"0000" when x"0C82",
			x"0000" when x"0C83",
			x"0000" when x"0C84",
			x"0000" when x"0C85",
			x"0000" when x"0C86",
			x"0000" when x"0C87",
			x"0000" when x"0C88",
			x"0000" when x"0C89",
			x"0000" when x"0C8A",
			x"0000" when x"0C8B",
			x"0000" when x"0C8C",
			x"0000" when x"0C8D",
			x"0000" when x"0C8E",
			x"0000" when x"0C8F",
			x"0000" when x"0C90",
			x"0000" when x"0C91",
			x"0000" when x"0C92",
			x"0000" when x"0C93",
			x"0000" when x"0C94",
			x"0000" when x"0C95",
			x"0000" when x"0C96",
			x"0000" when x"0C97",
			x"0000" when x"0C98",
			x"0000" when x"0C99",
			x"0000" when x"0C9A",
			x"0000" when x"0C9B",
			x"0000" when x"0C9C",
			x"0000" when x"0C9D",
			x"0000" when x"0C9E",
			x"0000" when x"0C9F",
			x"0000" when x"0CA0",
			x"0000" when x"0CA1",
			x"0000" when x"0CA2",
			x"0000" when x"0CA3",
			x"0000" when x"0CA4",
			x"0000" when x"0CA5",
			x"0000" when x"0CA6",
			x"0000" when x"0CA7",
			x"0000" when x"0CA8",
			x"0000" when x"0CA9",
			x"0000" when x"0CAA",
			x"0000" when x"0CAB",
			x"0000" when x"0CAC",
			x"0000" when x"0CAD",
			x"0000" when x"0CAE",
			x"0000" when x"0CAF",
			x"0000" when x"0CB0",
			x"0000" when x"0CB1",
			x"0000" when x"0CB2",
			x"0000" when x"0CB3",
			x"0000" when x"0CB4",
			x"0000" when x"0CB5",
			x"0000" when x"0CB6",
			x"0000" when x"0CB7",
			x"0000" when x"0CB8",
			x"0000" when x"0CB9",
			x"0000" when x"0CBA",
			x"0000" when x"0CBB",
			x"0000" when x"0CBC",
			x"0000" when x"0CBD",
			x"0000" when x"0CBE",
			x"0000" when x"0CBF",
			x"0000" when x"0CC0",
			x"0000" when x"0CC1",
			x"0000" when x"0CC2",
			x"0000" when x"0CC3",
			x"0000" when x"0CC4",
			x"0000" when x"0CC5",
			x"0000" when x"0CC6",
			x"0000" when x"0CC7",
			x"0000" when x"0CC8",
			x"0000" when x"0CC9",
			x"0000" when x"0CCA",
			x"0000" when x"0CCB",
			x"0000" when x"0CCC",
			x"0000" when x"0CCD",
			x"0000" when x"0CCE",
			x"0000" when x"0CCF",
			x"0000" when x"0CD0",
			x"0000" when x"0CD1",
			x"0000" when x"0CD2",
			x"0000" when x"0CD3",
			x"0000" when x"0CD4",
			x"0000" when x"0CD5",
			x"0000" when x"0CD6",
			x"0000" when x"0CD7",
			x"0000" when x"0CD8",
			x"0000" when x"0CD9",
			x"0000" when x"0CDA",
			x"0000" when x"0CDB",
			x"0000" when x"0CDC",
			x"0000" when x"0CDD",
			x"0000" when x"0CDE",
			x"0000" when x"0CDF",
			x"0000" when x"0CE0",
			x"0000" when x"0CE1",
			x"0000" when x"0CE2",
			x"0000" when x"0CE3",
			x"0000" when x"0CE4",
			x"0000" when x"0CE5",
			x"0000" when x"0CE6",
			x"0000" when x"0CE7",
			x"0000" when x"0CE8",
			x"0000" when x"0CE9",
			x"0000" when x"0CEA",
			x"0000" when x"0CEB",
			x"0000" when x"0CEC",
			x"0000" when x"0CED",
			x"0000" when x"0CEE",
			x"0000" when x"0CEF",
			x"0000" when x"0CF0",
			x"0000" when x"0CF1",
			x"0000" when x"0CF2",
			x"0000" when x"0CF3",
			x"0000" when x"0CF4",
			x"0000" when x"0CF5",
			x"0000" when x"0CF6",
			x"0000" when x"0CF7",
			x"0000" when x"0CF8",
			x"0000" when x"0CF9",
			x"0000" when x"0CFA",
			x"0000" when x"0CFB",
			x"0000" when x"0CFC",
			x"0000" when x"0CFD",
			x"0000" when x"0CFE",
			x"0000" when x"0CFF",
			x"0000" when x"0D00",
			x"0000" when x"0D01",
			x"0000" when x"0D02",
			x"0000" when x"0D03",
			x"0000" when x"0D04",
			x"0000" when x"0D05",
			x"0000" when x"0D06",
			x"0000" when x"0D07",
			x"0000" when x"0D08",
			x"0000" when x"0D09",
			x"0000" when x"0D0A",
			x"0000" when x"0D0B",
			x"0000" when x"0D0C",
			x"0000" when x"0D0D",
			x"0000" when x"0D0E",
			x"0000" when x"0D0F",
			x"0000" when x"0D10",
			x"0000" when x"0D11",
			x"0000" when x"0D12",
			x"0000" when x"0D13",
			x"0000" when x"0D14",
			x"0000" when x"0D15",
			x"0000" when x"0D16",
			x"0000" when x"0D17",
			x"0000" when x"0D18",
			x"0000" when x"0D19",
			x"0000" when x"0D1A",
			x"0000" when x"0D1B",
			x"0000" when x"0D1C",
			x"0000" when x"0D1D",
			x"0000" when x"0D1E",
			x"0000" when x"0D1F",
			x"0000" when x"0D20",
			x"0000" when x"0D21",
			x"0000" when x"0D22",
			x"0000" when x"0D23",
			x"0000" when x"0D24",
			x"0000" when x"0D25",
			x"0000" when x"0D26",
			x"0000" when x"0D27",
			x"0000" when x"0D28",
			x"0000" when x"0D29",
			x"0000" when x"0D2A",
			x"0000" when x"0D2B",
			x"0000" when x"0D2C",
			x"0000" when x"0D2D",
			x"0000" when x"0D2E",
			x"0000" when x"0D2F",
			x"0000" when x"0D30",
			x"0000" when x"0D31",
			x"0000" when x"0D32",
			x"0000" when x"0D33",
			x"0000" when x"0D34",
			x"0000" when x"0D35",
			x"0000" when x"0D36",
			x"0000" when x"0D37",
			x"0000" when x"0D38",
			x"0000" when x"0D39",
			x"0000" when x"0D3A",
			x"0000" when x"0D3B",
			x"0000" when x"0D3C",
			x"0000" when x"0D3D",
			x"0000" when x"0D3E",
			x"0000" when x"0D3F",
			x"0000" when x"0D40",
			x"0000" when x"0D41",
			x"0000" when x"0D42",
			x"0000" when x"0D43",
			x"0000" when x"0D44",
			x"0000" when x"0D45",
			x"0000" when x"0D46",
			x"0000" when x"0D47",
			x"0000" when x"0D48",
			x"0000" when x"0D49",
			x"0000" when x"0D4A",
			x"0000" when x"0D4B",
			x"0000" when x"0D4C",
			x"0000" when x"0D4D",
			x"0000" when x"0D4E",
			x"0000" when x"0D4F",
			x"0000" when x"0D50",
			x"0000" when x"0D51",
			x"0000" when x"0D52",
			x"0000" when x"0D53",
			x"0000" when x"0D54",
			x"0000" when x"0D55",
			x"0000" when x"0D56",
			x"0000" when x"0D57",
			x"0000" when x"0D58",
			x"0000" when x"0D59",
			x"0000" when x"0D5A",
			x"0000" when x"0D5B",
			x"0000" when x"0D5C",
			x"0000" when x"0D5D",
			x"0000" when x"0D5E",
			x"0000" when x"0D5F",
			x"0000" when x"0D60",
			x"0000" when x"0D61",
			x"0000" when x"0D62",
			x"0000" when x"0D63",
			x"0000" when x"0D64",
			x"0000" when x"0D65",
			x"0000" when x"0D66",
			x"0000" when x"0D67",
			x"0000" when x"0D68",
			x"0000" when x"0D69",
			x"0000" when x"0D6A",
			x"0000" when x"0D6B",
			x"0000" when x"0D6C",
			x"0000" when x"0D6D",
			x"0000" when x"0D6E",
			x"0000" when x"0D6F",
			x"0000" when x"0D70",
			x"0000" when x"0D71",
			x"0000" when x"0D72",
			x"0000" when x"0D73",
			x"0000" when x"0D74",
			x"0000" when x"0D75",
			x"0000" when x"0D76",
			x"0000" when x"0D77",
			x"0000" when x"0D78",
			x"0000" when x"0D79",
			x"0000" when x"0D7A",
			x"0000" when x"0D7B",
			x"0000" when x"0D7C",
			x"0000" when x"0D7D",
			x"0000" when x"0D7E",
			x"0000" when x"0D7F",
			x"0000" when x"0D80",
			x"0000" when x"0D81",
			x"0000" when x"0D82",
			x"0000" when x"0D83",
			x"0000" when x"0D84",
			x"0000" when x"0D85",
			x"0000" when x"0D86",
			x"0000" when x"0D87",
			x"0000" when x"0D88",
			x"0000" when x"0D89",
			x"0000" when x"0D8A",
			x"0000" when x"0D8B",
			x"0000" when x"0D8C",
			x"0000" when x"0D8D",
			x"0000" when x"0D8E",
			x"0000" when x"0D8F",
			x"0000" when x"0D90",
			x"0000" when x"0D91",
			x"0000" when x"0D92",
			x"0000" when x"0D93",
			x"0000" when x"0D94",
			x"0000" when x"0D95",
			x"0000" when x"0D96",
			x"0000" when x"0D97",
			x"0000" when x"0D98",
			x"0000" when x"0D99",
			x"0000" when x"0D9A",
			x"0000" when x"0D9B",
			x"0000" when x"0D9C",
			x"0000" when x"0D9D",
			x"0000" when x"0D9E",
			x"0000" when x"0D9F",
			x"0000" when x"0DA0",
			x"0000" when x"0DA1",
			x"0000" when x"0DA2",
			x"0000" when x"0DA3",
			x"0000" when x"0DA4",
			x"0000" when x"0DA5",
			x"0000" when x"0DA6",
			x"0000" when x"0DA7",
			x"0000" when x"0DA8",
			x"0000" when x"0DA9",
			x"0000" when x"0DAA",
			x"0000" when x"0DAB",
			x"0000" when x"0DAC",
			x"0000" when x"0DAD",
			x"0000" when x"0DAE",
			x"0000" when x"0DAF",
			x"0000" when x"0DB0",
			x"0000" when x"0DB1",
			x"0000" when x"0DB2",
			x"0000" when x"0DB3",
			x"0000" when x"0DB4",
			x"0000" when x"0DB5",
			x"0000" when x"0DB6",
			x"0000" when x"0DB7",
			x"0000" when x"0DB8",
			x"0000" when x"0DB9",
			x"0000" when x"0DBA",
			x"0000" when x"0DBB",
			x"0000" when x"0DBC",
			x"0000" when x"0DBD",
			x"0000" when x"0DBE",
			x"0000" when x"0DBF",
			x"0000" when x"0DC0",
			x"0000" when x"0DC1",
			x"0000" when x"0DC2",
			x"0000" when x"0DC3",
			x"0000" when x"0DC4",
			x"0000" when x"0DC5",
			x"0000" when x"0DC6",
			x"0000" when x"0DC7",
			x"0000" when x"0DC8",
			x"0000" when x"0DC9",
			x"0000" when x"0DCA",
			x"0000" when x"0DCB",
			x"0000" when x"0DCC",
			x"0000" when x"0DCD",
			x"0000" when x"0DCE",
			x"0000" when x"0DCF",
			x"0000" when x"0DD0",
			x"0000" when x"0DD1",
			x"0000" when x"0DD2",
			x"0000" when x"0DD3",
			x"0000" when x"0DD4",
			x"0000" when x"0DD5",
			x"0000" when x"0DD6",
			x"0000" when x"0DD7",
			x"0000" when x"0DD8",
			x"0000" when x"0DD9",
			x"0000" when x"0DDA",
			x"0000" when x"0DDB",
			x"0000" when x"0DDC",
			x"0000" when x"0DDD",
			x"0000" when x"0DDE",
			x"0000" when x"0DDF",
			x"0000" when x"0DE0",
			x"0000" when x"0DE1",
			x"0000" when x"0DE2",
			x"0000" when x"0DE3",
			x"0000" when x"0DE4",
			x"0000" when x"0DE5",
			x"0000" when x"0DE6",
			x"0000" when x"0DE7",
			x"0000" when x"0DE8",
			x"0000" when x"0DE9",
			x"0000" when x"0DEA",
			x"0000" when x"0DEB",
			x"0000" when x"0DEC",
			x"0000" when x"0DED",
			x"0000" when x"0DEE",
			x"0000" when x"0DEF",
			x"0000" when x"0DF0",
			x"0000" when x"0DF1",
			x"0000" when x"0DF2",
			x"0000" when x"0DF3",
			x"0000" when x"0DF4",
			x"0000" when x"0DF5",
			x"0000" when x"0DF6",
			x"0000" when x"0DF7",
			x"0000" when x"0DF8",
			x"0000" when x"0DF9",
			x"0000" when x"0DFA",
			x"0000" when x"0DFB",
			x"0000" when x"0DFC",
			x"0000" when x"0DFD",
			x"0000" when x"0DFE",
			x"0000" when x"0DFF",
			x"0000" when x"0E00",
			x"0000" when x"0E01",
			x"0000" when x"0E02",
			x"0000" when x"0E03",
			x"0000" when x"0E04",
			x"0000" when x"0E05",
			x"0000" when x"0E06",
			x"0000" when x"0E07",
			x"0000" when x"0E08",
			x"0000" when x"0E09",
			x"0000" when x"0E0A",
			x"0000" when x"0E0B",
			x"0000" when x"0E0C",
			x"0000" when x"0E0D",
			x"0000" when x"0E0E",
			x"0000" when x"0E0F",
			x"0000" when x"0E10",
			x"0000" when x"0E11",
			x"0000" when x"0E12",
			x"0000" when x"0E13",
			x"0000" when x"0E14",
			x"0000" when x"0E15",
			x"0000" when x"0E16",
			x"0000" when x"0E17",
			x"0000" when x"0E18",
			x"0000" when x"0E19",
			x"0000" when x"0E1A",
			x"0000" when x"0E1B",
			x"0000" when x"0E1C",
			x"0000" when x"0E1D",
			x"0000" when x"0E1E",
			x"0000" when x"0E1F",
			x"0000" when x"0E20",
			x"0000" when x"0E21",
			x"0000" when x"0E22",
			x"0000" when x"0E23",
			x"0000" when x"0E24",
			x"0000" when x"0E25",
			x"0000" when x"0E26",
			x"0000" when x"0E27",
			x"0000" when x"0E28",
			x"0000" when x"0E29",
			x"0000" when x"0E2A",
			x"0000" when x"0E2B",
			x"0000" when x"0E2C",
			x"0000" when x"0E2D",
			x"0000" when x"0E2E",
			x"0000" when x"0E2F",
			x"0000" when x"0E30",
			x"0000" when x"0E31",
			x"0000" when x"0E32",
			x"0000" when x"0E33",
			x"0000" when x"0E34",
			x"0000" when x"0E35",
			x"0000" when x"0E36",
			x"0000" when x"0E37",
			x"0000" when x"0E38",
			x"0000" when x"0E39",
			x"0000" when x"0E3A",
			x"0000" when x"0E3B",
			x"0000" when x"0E3C",
			x"0000" when x"0E3D",
			x"0000" when x"0E3E",
			x"0000" when x"0E3F",
			x"0000" when x"0E40",
			x"0000" when x"0E41",
			x"0000" when x"0E42",
			x"0000" when x"0E43",
			x"0000" when x"0E44",
			x"0000" when x"0E45",
			x"0000" when x"0E46",
			x"0000" when x"0E47",
			x"0000" when x"0E48",
			x"0000" when x"0E49",
			x"0000" when x"0E4A",
			x"0000" when x"0E4B",
			x"0000" when x"0E4C",
			x"0000" when x"0E4D",
			x"0000" when x"0E4E",
			x"0000" when x"0E4F",
			x"0000" when x"0E50",
			x"0000" when x"0E51",
			x"0000" when x"0E52",
			x"0000" when x"0E53",
			x"0000" when x"0E54",
			x"0000" when x"0E55",
			x"0000" when x"0E56",
			x"0000" when x"0E57",
			x"0000" when x"0E58",
			x"0000" when x"0E59",
			x"0000" when x"0E5A",
			x"0000" when x"0E5B",
			x"0000" when x"0E5C",
			x"0000" when x"0E5D",
			x"0000" when x"0E5E",
			x"0000" when x"0E5F",
			x"0000" when x"0E60",
			x"0000" when x"0E61",
			x"0000" when x"0E62",
			x"0000" when x"0E63",
			x"0000" when x"0E64",
			x"0000" when x"0E65",
			x"0000" when x"0E66",
			x"0000" when x"0E67",
			x"0000" when x"0E68",
			x"0000" when x"0E69",
			x"0000" when x"0E6A",
			x"0000" when x"0E6B",
			x"0000" when x"0E6C",
			x"0000" when x"0E6D",
			x"0000" when x"0E6E",
			x"0000" when x"0E6F",
			x"0000" when x"0E70",
			x"0000" when x"0E71",
			x"0000" when x"0E72",
			x"0000" when x"0E73",
			x"0000" when x"0E74",
			x"0000" when x"0E75",
			x"0000" when x"0E76",
			x"0000" when x"0E77",
			x"0000" when x"0E78",
			x"0000" when x"0E79",
			x"0000" when x"0E7A",
			x"0000" when x"0E7B",
			x"0000" when x"0E7C",
			x"0000" when x"0E7D",
			x"0000" when x"0E7E",
			x"0000" when x"0E7F",
			x"0000" when x"0E80",
			x"0000" when x"0E81",
			x"0000" when x"0E82",
			x"0000" when x"0E83",
			x"0000" when x"0E84",
			x"0000" when x"0E85",
			x"0000" when x"0E86",
			x"0000" when x"0E87",
			x"0000" when x"0E88",
			x"0000" when x"0E89",
			x"0000" when x"0E8A",
			x"0000" when x"0E8B",
			x"0000" when x"0E8C",
			x"0000" when x"0E8D",
			x"0000" when x"0E8E",
			x"0000" when x"0E8F",
			x"0000" when x"0E90",
			x"0000" when x"0E91",
			x"0000" when x"0E92",
			x"0000" when x"0E93",
			x"0000" when x"0E94",
			x"0000" when x"0E95",
			x"0000" when x"0E96",
			x"0000" when x"0E97",
			x"0000" when x"0E98",
			x"0000" when x"0E99",
			x"0000" when x"0E9A",
			x"0000" when x"0E9B",
			x"0000" when x"0E9C",
			x"0000" when x"0E9D",
			x"0000" when x"0E9E",
			x"0000" when x"0E9F",
			x"0000" when x"0EA0",
			x"0000" when x"0EA1",
			x"0000" when x"0EA2",
			x"0000" when x"0EA3",
			x"0000" when x"0EA4",
			x"0000" when x"0EA5",
			x"0000" when x"0EA6",
			x"0000" when x"0EA7",
			x"0000" when x"0EA8",
			x"0000" when x"0EA9",
			x"0000" when x"0EAA",
			x"0000" when x"0EAB",
			x"0000" when x"0EAC",
			x"0000" when x"0EAD",
			x"0000" when x"0EAE",
			x"0000" when x"0EAF",
			x"0000" when x"0EB0",
			x"0000" when x"0EB1",
			x"0000" when x"0EB2",
			x"0000" when x"0EB3",
			x"0000" when x"0EB4",
			x"0000" when x"0EB5",
			x"0000" when x"0EB6",
			x"0000" when x"0EB7",
			x"0000" when x"0EB8",
			x"0000" when x"0EB9",
			x"0000" when x"0EBA",
			x"0000" when x"0EBB",
			x"0000" when x"0EBC",
			x"0000" when x"0EBD",
			x"0000" when x"0EBE",
			x"0000" when x"0EBF",
			x"0000" when x"0EC0",
			x"0000" when x"0EC1",
			x"0000" when x"0EC2",
			x"0000" when x"0EC3",
			x"0000" when x"0EC4",
			x"0000" when x"0EC5",
			x"0000" when x"0EC6",
			x"0000" when x"0EC7",
			x"0000" when x"0EC8",
			x"0000" when x"0EC9",
			x"0000" when x"0ECA",
			x"0000" when x"0ECB",
			x"0000" when x"0ECC",
			x"0000" when x"0ECD",
			x"0000" when x"0ECE",
			x"0000" when x"0ECF",
			x"0000" when x"0ED0",
			x"0000" when x"0ED1",
			x"0000" when x"0ED2",
			x"0000" when x"0ED3",
			x"0000" when x"0ED4",
			x"0000" when x"0ED5",
			x"0000" when x"0ED6",
			x"0000" when x"0ED7",
			x"0000" when x"0ED8",
			x"0000" when x"0ED9",
			x"0000" when x"0EDA",
			x"0000" when x"0EDB",
			x"0000" when x"0EDC",
			x"0000" when x"0EDD",
			x"0000" when x"0EDE",
			x"0000" when x"0EDF",
			x"0000" when x"0EE0",
			x"0000" when x"0EE1",
			x"0000" when x"0EE2",
			x"0000" when x"0EE3",
			x"0000" when x"0EE4",
			x"0000" when x"0EE5",
			x"0000" when x"0EE6",
			x"0000" when x"0EE7",
			x"0000" when x"0EE8",
			x"0000" when x"0EE9",
			x"0000" when x"0EEA",
			x"0000" when x"0EEB",
			x"0000" when x"0EEC",
			x"0000" when x"0EED",
			x"0000" when x"0EEE",
			x"0000" when x"0EEF",
			x"0000" when x"0EF0",
			x"0000" when x"0EF1",
			x"0000" when x"0EF2",
			x"0000" when x"0EF3",
			x"0000" when x"0EF4",
			x"0000" when x"0EF5",
			x"0000" when x"0EF6",
			x"0000" when x"0EF7",
			x"0000" when x"0EF8",
			x"0000" when x"0EF9",
			x"0000" when x"0EFA",
			x"0000" when x"0EFB",
			x"0000" when x"0EFC",
			x"0000" when x"0EFD",
			x"0000" when x"0EFE",
			x"0000" when x"0EFF",
			x"0000" when x"0F00",
			x"0000" when x"0F01",
			x"0000" when x"0F02",
			x"0000" when x"0F03",
			x"0000" when x"0F04",
			x"0000" when x"0F05",
			x"0000" when x"0F06",
			x"0000" when x"0F07",
			x"0000" when x"0F08",
			x"0000" when x"0F09",
			x"0000" when x"0F0A",
			x"0000" when x"0F0B",
			x"0000" when x"0F0C",
			x"0000" when x"0F0D",
			x"0000" when x"0F0E",
			x"0000" when x"0F0F",
			x"0000" when x"0F10",
			x"0000" when x"0F11",
			x"0000" when x"0F12",
			x"0000" when x"0F13",
			x"0000" when x"0F14",
			x"0000" when x"0F15",
			x"0000" when x"0F16",
			x"0000" when x"0F17",
			x"0000" when x"0F18",
			x"0000" when x"0F19",
			x"0000" when x"0F1A",
			x"0000" when x"0F1B",
			x"0000" when x"0F1C",
			x"0000" when x"0F1D",
			x"0000" when x"0F1E",
			x"0000" when x"0F1F",
			x"0000" when x"0F20",
			x"0000" when x"0F21",
			x"0000" when x"0F22",
			x"0000" when x"0F23",
			x"0000" when x"0F24",
			x"0000" when x"0F25",
			x"0000" when x"0F26",
			x"0000" when x"0F27",
			x"0000" when x"0F28",
			x"0000" when x"0F29",
			x"0000" when x"0F2A",
			x"0000" when x"0F2B",
			x"0000" when x"0F2C",
			x"0000" when x"0F2D",
			x"0000" when x"0F2E",
			x"0000" when x"0F2F",
			x"0000" when x"0F30",
			x"0000" when x"0F31",
			x"0000" when x"0F32",
			x"0000" when x"0F33",
			x"0000" when x"0F34",
			x"0000" when x"0F35",
			x"0000" when x"0F36",
			x"0000" when x"0F37",
			x"0000" when x"0F38",
			x"0000" when x"0F39",
			x"0000" when x"0F3A",
			x"0000" when x"0F3B",
			x"0000" when x"0F3C",
			x"0000" when x"0F3D",
			x"0000" when x"0F3E",
			x"0000" when x"0F3F",
			x"0000" when x"0F40",
			x"0000" when x"0F41",
			x"0000" when x"0F42",
			x"0000" when x"0F43",
			x"0000" when x"0F44",
			x"0000" when x"0F45",
			x"0000" when x"0F46",
			x"0000" when x"0F47",
			x"0000" when x"0F48",
			x"0000" when x"0F49",
			x"0000" when x"0F4A",
			x"0000" when x"0F4B",
			x"0000" when x"0F4C",
			x"0000" when x"0F4D",
			x"0000" when x"0F4E",
			x"0000" when x"0F4F",
			x"0000" when x"0F50",
			x"0000" when x"0F51",
			x"0000" when x"0F52",
			x"0000" when x"0F53",
			x"0000" when x"0F54",
			x"0000" when x"0F55",
			x"0000" when x"0F56",
			x"0000" when x"0F57",
			x"0000" when x"0F58",
			x"0000" when x"0F59",
			x"0000" when x"0F5A",
			x"0000" when x"0F5B",
			x"0000" when x"0F5C",
			x"0000" when x"0F5D",
			x"0000" when x"0F5E",
			x"0000" when x"0F5F",
			x"0000" when x"0F60",
			x"0000" when x"0F61",
			x"0000" when x"0F62",
			x"0000" when x"0F63",
			x"0000" when x"0F64",
			x"0000" when x"0F65",
			x"0000" when x"0F66",
			x"0000" when x"0F67",
			x"0000" when x"0F68",
			x"0000" when x"0F69",
			x"0000" when x"0F6A",
			x"0000" when x"0F6B",
			x"0000" when x"0F6C",
			x"0000" when x"0F6D",
			x"0000" when x"0F6E",
			x"0000" when x"0F6F",
			x"0000" when x"0F70",
			x"0000" when x"0F71",
			x"0000" when x"0F72",
			x"0000" when x"0F73",
			x"0000" when x"0F74",
			x"0000" when x"0F75",
			x"0000" when x"0F76",
			x"0000" when x"0F77",
			x"0000" when x"0F78",
			x"0000" when x"0F79",
			x"0000" when x"0F7A",
			x"0000" when x"0F7B",
			x"0000" when x"0F7C",
			x"0000" when x"0F7D",
			x"0000" when x"0F7E",
			x"0000" when x"0F7F",
			x"0000" when x"0F80",
			x"0000" when x"0F81",
			x"0000" when x"0F82",
			x"0000" when x"0F83",
			x"0000" when x"0F84",
			x"0000" when x"0F85",
			x"0000" when x"0F86",
			x"0000" when x"0F87",
			x"0000" when x"0F88",
			x"0000" when x"0F89",
			x"0000" when x"0F8A",
			x"0000" when x"0F8B",
			x"0000" when x"0F8C",
			x"0000" when x"0F8D",
			x"0000" when x"0F8E",
			x"0000" when x"0F8F",
			x"0000" when x"0F90",
			x"0000" when x"0F91",
			x"0000" when x"0F92",
			x"0000" when x"0F93",
			x"0000" when x"0F94",
			x"0000" when x"0F95",
			x"0000" when x"0F96",
			x"0000" when x"0F97",
			x"0000" when x"0F98",
			x"0000" when x"0F99",
			x"0000" when x"0F9A",
			x"0000" when x"0F9B",
			x"0000" when x"0F9C",
			x"0000" when x"0F9D",
			x"0000" when x"0F9E",
			x"0000" when x"0F9F",
			x"0000" when x"0FA0",
			x"0000" when x"0FA1",
			x"0000" when x"0FA2",
			x"0000" when x"0FA3",
			x"0000" when x"0FA4",
			x"0000" when x"0FA5",
			x"0000" when x"0FA6",
			x"0000" when x"0FA7",
			x"0000" when x"0FA8",
			x"0000" when x"0FA9",
			x"0000" when x"0FAA",
			x"0000" when x"0FAB",
			x"0000" when x"0FAC",
			x"0000" when x"0FAD",
			x"0000" when x"0FAE",
			x"0000" when x"0FAF",
			x"0000" when x"0FB0",
			x"0000" when x"0FB1",
			x"0000" when x"0FB2",
			x"0000" when x"0FB3",
			x"0000" when x"0FB4",
			x"0000" when x"0FB5",
			x"0000" when x"0FB6",
			x"0000" when x"0FB7",
			x"0000" when x"0FB8",
			x"0000" when x"0FB9",
			x"0000" when x"0FBA",
			x"0000" when x"0FBB",
			x"0000" when x"0FBC",
			x"0000" when x"0FBD",
			x"0000" when x"0FBE",
			x"0000" when x"0FBF",
			x"0000" when x"0FC0",
			x"0000" when x"0FC1",
			x"0000" when x"0FC2",
			x"0000" when x"0FC3",
			x"0000" when x"0FC4",
			x"0000" when x"0FC5",
			x"0000" when x"0FC6",
			x"0000" when x"0FC7",
			x"0000" when x"0FC8",
			x"0000" when x"0FC9",
			x"0000" when x"0FCA",
			x"0000" when x"0FCB",
			x"0000" when x"0FCC",
			x"0000" when x"0FCD",
			x"0000" when x"0FCE",
			x"0000" when x"0FCF",
			x"0000" when x"0FD0",
			x"0000" when x"0FD1",
			x"0000" when x"0FD2",
			x"0000" when x"0FD3",
			x"0000" when x"0FD4",
			x"0000" when x"0FD5",
			x"0000" when x"0FD6",
			x"0000" when x"0FD7",
			x"0000" when x"0FD8",
			x"0000" when x"0FD9",
			x"0000" when x"0FDA",
			x"0000" when x"0FDB",
			x"0000" when x"0FDC",
			x"0000" when x"0FDD",
			x"0000" when x"0FDE",
			x"0000" when x"0FDF",
			x"0000" when x"0FE0",
			x"0000" when x"0FE1",
			x"0000" when x"0FE2",
			x"0000" when x"0FE3",
			x"0000" when x"0FE4",
			x"0000" when x"0FE5",
			x"0000" when x"0FE6",
			x"0000" when x"0FE7",
			x"0000" when x"0FE8",
			x"0000" when x"0FE9",
			x"0000" when x"0FEA",
			x"0000" when x"0FEB",
			x"0000" when x"0FEC",
			x"0000" when x"0FED",
			x"0000" when x"0FEE",
			x"0000" when x"0FEF",
			x"0000" when x"0FF0",
			x"0000" when x"0FF1",
			x"0000" when x"0FF2",
			x"0000" when x"0FF3",
			x"0000" when x"0FF4",
			x"0000" when x"0FF5",
			x"0000" when x"0FF6",
			x"0000" when x"0FF7",
			x"0000" when x"0FF8",
			x"0000" when x"0FF9",
			x"0000" when x"0FFA",
			x"0000" when x"0FFB",
			x"0000" when x"0FFC",
			x"0000" when x"0FFD",
			x"0000" when x"0FFE",
			x"0000" when x"0FFF",
			x"0000" when x"1000",
			x"0000" when x"1001",
			x"0000" when x"1002",
			x"0000" when x"1003",
			x"0000" when x"1004",
			x"0000" when x"1005",
			x"0000" when x"1006",
			x"0000" when x"1007",
			x"0000" when x"1008",
			x"0000" when x"1009",
			x"0000" when x"100A",
			x"0000" when x"100B",
			x"0000" when x"100C",
			x"0000" when x"100D",
			x"0000" when x"100E",
			x"0000" when x"100F",
			x"0000" when x"1010",
			x"0000" when x"1011",
			x"0000" when x"1012",
			x"0000" when x"1013",
			x"0000" when x"1014",
			x"0000" when x"1015",
			x"0000" when x"1016",
			x"0000" when x"1017",
			x"0000" when x"1018",
			x"0000" when x"1019",
			x"0000" when x"101A",
			x"0000" when x"101B",
			x"0000" when x"101C",
			x"0000" when x"101D",
			x"0000" when x"101E",
			x"0000" when x"101F",
			x"0000" when x"1020",
			x"0000" when x"1021",
			x"0000" when x"1022",
			x"0000" when x"1023",
			x"0000" when x"1024",
			x"0000" when x"1025",
			x"0000" when x"1026",
			x"0000" when x"1027",
			x"0000" when x"1028",
			x"0000" when x"1029",
			x"0000" when x"102A",
			x"0000" when x"102B",
			x"0000" when x"102C",
			x"0000" when x"102D",
			x"0000" when x"102E",
			x"0000" when x"102F",
			x"0000" when x"1030",
			x"0000" when x"1031",
			x"0000" when x"1032",
			x"0000" when x"1033",
			x"0000" when x"1034",
			x"0000" when x"1035",
			x"0000" when x"1036",
			x"0000" when x"1037",
			x"0000" when x"1038",
			x"0000" when x"1039",
			x"0000" when x"103A",
			x"0000" when x"103B",
			x"0000" when x"103C",
			x"0000" when x"103D",
			x"0000" when x"103E",
			x"0000" when x"103F",
			x"0000" when x"1040",
			x"0000" when x"1041",
			x"0000" when x"1042",
			x"0000" when x"1043",
			x"0000" when x"1044",
			x"0000" when x"1045",
			x"0000" when x"1046",
			x"0000" when x"1047",
			x"0000" when x"1048",
			x"0000" when x"1049",
			x"0000" when x"104A",
			x"0000" when x"104B",
			x"0000" when x"104C",
			x"0000" when x"104D",
			x"0000" when x"104E",
			x"0000" when x"104F",
			x"0000" when x"1050",
			x"0000" when x"1051",
			x"0000" when x"1052",
			x"0000" when x"1053",
			x"0000" when x"1054",
			x"0000" when x"1055",
			x"0000" when x"1056",
			x"0000" when x"1057",
			x"0000" when x"1058",
			x"0000" when x"1059",
			x"0000" when x"105A",
			x"0000" when x"105B",
			x"0000" when x"105C",
			x"0000" when x"105D",
			x"0000" when x"105E",
			x"0000" when x"105F",
			x"0000" when x"1060",
			x"0000" when x"1061",
			x"0000" when x"1062",
			x"0000" when x"1063",
			x"0000" when x"1064",
			x"0000" when x"1065",
			x"0000" when x"1066",
			x"0000" when x"1067",
			x"0000" when x"1068",
			x"0000" when x"1069",
			x"0000" when x"106A",
			x"0000" when x"106B",
			x"0000" when x"106C",
			x"0000" when x"106D",
			x"0000" when x"106E",
			x"0000" when x"106F",
			x"0000" when x"1070",
			x"0000" when x"1071",
			x"0000" when x"1072",
			x"0000" when x"1073",
			x"0000" when x"1074",
			x"0000" when x"1075",
			x"0000" when x"1076",
			x"0000" when x"1077",
			x"0000" when x"1078",
			x"0000" when x"1079",
			x"0000" when x"107A",
			x"0000" when x"107B",
			x"0000" when x"107C",
			x"0000" when x"107D",
			x"0000" when x"107E",
			x"0000" when x"107F",
			x"0000" when x"1080",
			x"0000" when x"1081",
			x"0000" when x"1082",
			x"0000" when x"1083",
			x"0000" when x"1084",
			x"0000" when x"1085",
			x"0000" when x"1086",
			x"0000" when x"1087",
			x"0000" when x"1088",
			x"0000" when x"1089",
			x"0000" when x"108A",
			x"0000" when x"108B",
			x"0000" when x"108C",
			x"0000" when x"108D",
			x"0000" when x"108E",
			x"0000" when x"108F",
			x"0000" when x"1090",
			x"0000" when x"1091",
			x"0000" when x"1092",
			x"0000" when x"1093",
			x"0000" when x"1094",
			x"0000" when x"1095",
			x"0000" when x"1096",
			x"0000" when x"1097",
			x"0000" when x"1098",
			x"0000" when x"1099",
			x"0000" when x"109A",
			x"0000" when x"109B",
			x"0000" when x"109C",
			x"0000" when x"109D",
			x"0000" when x"109E",
			x"0000" when x"109F",
			x"0000" when x"10A0",
			x"0000" when x"10A1",
			x"0000" when x"10A2",
			x"0000" when x"10A3",
			x"0000" when x"10A4",
			x"0000" when x"10A5",
			x"0000" when x"10A6",
			x"0000" when x"10A7",
			x"0000" when x"10A8",
			x"0000" when x"10A9",
			x"0000" when x"10AA",
			x"0000" when x"10AB",
			x"0000" when x"10AC",
			x"0000" when x"10AD",
			x"0000" when x"10AE",
			x"0000" when x"10AF",
			x"0000" when x"10B0",
			x"0000" when x"10B1",
			x"0000" when x"10B2",
			x"0000" when x"10B3",
			x"0000" when x"10B4",
			x"0000" when x"10B5",
			x"0000" when x"10B6",
			x"0000" when x"10B7",
			x"0000" when x"10B8",
			x"0000" when x"10B9",
			x"0000" when x"10BA",
			x"0000" when x"10BB",
			x"0000" when x"10BC",
			x"0000" when x"10BD",
			x"0000" when x"10BE",
			x"0000" when x"10BF",
			x"0000" when x"10C0",
			x"0000" when x"10C1",
			x"0000" when x"10C2",
			x"0000" when x"10C3",
			x"0000" when x"10C4",
			x"0000" when x"10C5",
			x"0000" when x"10C6",
			x"0000" when x"10C7",
			x"0000" when x"10C8",
			x"0000" when x"10C9",
			x"0000" when x"10CA",
			x"0000" when x"10CB",
			x"0000" when x"10CC",
			x"0000" when x"10CD",
			x"0000" when x"10CE",
			x"0000" when x"10CF",
			x"0000" when x"10D0",
			x"0000" when x"10D1",
			x"0000" when x"10D2",
			x"0000" when x"10D3",
			x"0000" when x"10D4",
			x"0000" when x"10D5",
			x"0000" when x"10D6",
			x"0000" when x"10D7",
			x"0000" when x"10D8",
			x"0000" when x"10D9",
			x"0000" when x"10DA",
			x"0000" when x"10DB",
			x"0000" when x"10DC",
			x"0000" when x"10DD",
			x"0000" when x"10DE",
			x"0000" when x"10DF",
			x"0000" when x"10E0",
			x"0000" when x"10E1",
			x"0000" when x"10E2",
			x"0000" when x"10E3",
			x"0000" when x"10E4",
			x"0000" when x"10E5",
			x"0000" when x"10E6",
			x"0000" when x"10E7",
			x"0000" when x"10E8",
			x"0000" when x"10E9",
			x"0000" when x"10EA",
			x"0000" when x"10EB",
			x"0000" when x"10EC",
			x"0000" when x"10ED",
			x"0000" when x"10EE",
			x"0000" when x"10EF",
			x"0000" when x"10F0",
			x"0000" when x"10F1",
			x"0000" when x"10F2",
			x"0000" when x"10F3",
			x"0000" when x"10F4",
			x"0000" when x"10F5",
			x"0000" when x"10F6",
			x"0000" when x"10F7",
			x"0000" when x"10F8",
			x"0000" when x"10F9",
			x"0000" when x"10FA",
			x"0000" when x"10FB",
			x"0000" when x"10FC",
			x"0000" when x"10FD",
			x"0000" when x"10FE",
			x"0000" when x"10FF",
			x"0000" when x"1100",
			x"0000" when x"1101",
			x"0000" when x"1102",
			x"0000" when x"1103",
			x"0000" when x"1104",
			x"0000" when x"1105",
			x"0000" when x"1106",
			x"0000" when x"1107",
			x"0000" when x"1108",
			x"0000" when x"1109",
			x"0000" when x"110A",
			x"0000" when x"110B",
			x"0000" when x"110C",
			x"0000" when x"110D",
			x"0000" when x"110E",
			x"0000" when x"110F",
			x"0000" when x"1110",
			x"0000" when x"1111",
			x"0000" when x"1112",
			x"0000" when x"1113",
			x"0000" when x"1114",
			x"0000" when x"1115",
			x"0000" when x"1116",
			x"0000" when x"1117",
			x"0000" when x"1118",
			x"0000" when x"1119",
			x"0000" when x"111A",
			x"0000" when x"111B",
			x"0000" when x"111C",
			x"0000" when x"111D",
			x"0000" when x"111E",
			x"0000" when x"111F",
			x"0000" when x"1120",
			x"0000" when x"1121",
			x"0000" when x"1122",
			x"0000" when x"1123",
			x"0000" when x"1124",
			x"0000" when x"1125",
			x"0000" when x"1126",
			x"0000" when x"1127",
			x"0000" when x"1128",
			x"0000" when x"1129",
			x"0000" when x"112A",
			x"0000" when x"112B",
			x"0000" when x"112C",
			x"0000" when x"112D",
			x"0000" when x"112E",
			x"0000" when x"112F",
			x"0000" when x"1130",
			x"0000" when x"1131",
			x"0000" when x"1132",
			x"0000" when x"1133",
			x"0000" when x"1134",
			x"0000" when x"1135",
			x"0000" when x"1136",
			x"0000" when x"1137",
			x"0000" when x"1138",
			x"0000" when x"1139",
			x"0000" when x"113A",
			x"0000" when x"113B",
			x"0000" when x"113C",
			x"0000" when x"113D",
			x"0000" when x"113E",
			x"0000" when x"113F",
			x"0000" when x"1140",
			x"0000" when x"1141",
			x"0000" when x"1142",
			x"0000" when x"1143",
			x"0000" when x"1144",
			x"0000" when x"1145",
			x"0000" when x"1146",
			x"0000" when x"1147",
			x"0000" when x"1148",
			x"0000" when x"1149",
			x"0000" when x"114A",
			x"0000" when x"114B",
			x"0000" when x"114C",
			x"0000" when x"114D",
			x"0000" when x"114E",
			x"0000" when x"114F",
			x"0000" when x"1150",
			x"0000" when x"1151",
			x"0000" when x"1152",
			x"0000" when x"1153",
			x"0000" when x"1154",
			x"0000" when x"1155",
			x"0000" when x"1156",
			x"0000" when x"1157",
			x"0000" when x"1158",
			x"0000" when x"1159",
			x"0000" when x"115A",
			x"0000" when x"115B",
			x"0000" when x"115C",
			x"0000" when x"115D",
			x"0000" when x"115E",
			x"0000" when x"115F",
			x"0000" when x"1160",
			x"0000" when x"1161",
			x"0000" when x"1162",
			x"0000" when x"1163",
			x"0000" when x"1164",
			x"0000" when x"1165",
			x"0000" when x"1166",
			x"0000" when x"1167",
			x"0000" when x"1168",
			x"0000" when x"1169",
			x"0000" when x"116A",
			x"0000" when x"116B",
			x"0000" when x"116C",
			x"0000" when x"116D",
			x"0000" when x"116E",
			x"0000" when x"116F",
			x"0000" when x"1170",
			x"0000" when x"1171",
			x"0000" when x"1172",
			x"0000" when x"1173",
			x"0000" when x"1174",
			x"0000" when x"1175",
			x"0000" when x"1176",
			x"0000" when x"1177",
			x"0000" when x"1178",
			x"0000" when x"1179",
			x"0000" when x"117A",
			x"0000" when x"117B",
			x"0000" when x"117C",
			x"0000" when x"117D",
			x"0000" when x"117E",
			x"0000" when x"117F",
			x"0000" when x"1180",
			x"0000" when x"1181",
			x"0000" when x"1182",
			x"0000" when x"1183",
			x"0000" when x"1184",
			x"0000" when x"1185",
			x"0000" when x"1186",
			x"0000" when x"1187",
			x"0000" when x"1188",
			x"0000" when x"1189",
			x"0000" when x"118A",
			x"0000" when x"118B",
			x"0000" when x"118C",
			x"0000" when x"118D",
			x"0000" when x"118E",
			x"0000" when x"118F",
			x"0000" when x"1190",
			x"0000" when x"1191",
			x"0000" when x"1192",
			x"0000" when x"1193",
			x"0000" when x"1194",
			x"0000" when x"1195",
			x"0000" when x"1196",
			x"0000" when x"1197",
			x"0000" when x"1198",
			x"0000" when x"1199",
			x"0000" when x"119A",
			x"0000" when x"119B",
			x"0000" when x"119C",
			x"0000" when x"119D",
			x"0000" when x"119E",
			x"0000" when x"119F",
			x"0000" when x"11A0",
			x"0000" when x"11A1",
			x"0000" when x"11A2",
			x"0000" when x"11A3",
			x"0000" when x"11A4",
			x"0000" when x"11A5",
			x"0000" when x"11A6",
			x"0000" when x"11A7",
			x"0000" when x"11A8",
			x"0000" when x"11A9",
			x"0000" when x"11AA",
			x"0000" when x"11AB",
			x"0000" when x"11AC",
			x"0000" when x"11AD",
			x"0000" when x"11AE",
			x"0000" when x"11AF",
			x"0000" when x"11B0",
			x"0000" when x"11B1",
			x"0000" when x"11B2",
			x"0000" when x"11B3",
			x"0000" when x"11B4",
			x"0000" when x"11B5",
			x"0000" when x"11B6",
			x"0000" when x"11B7",
			x"0000" when x"11B8",
			x"0000" when x"11B9",
			x"0000" when x"11BA",
			x"0000" when x"11BB",
			x"0000" when x"11BC",
			x"0000" when x"11BD",
			x"0000" when x"11BE",
			x"0000" when x"11BF",
			x"0000" when x"11C0",
			x"0000" when x"11C1",
			x"0000" when x"11C2",
			x"0000" when x"11C3",
			x"0000" when x"11C4",
			x"0000" when x"11C5",
			x"0000" when x"11C6",
			x"0000" when x"11C7",
			x"0000" when x"11C8",
			x"0000" when x"11C9",
			x"0000" when x"11CA",
			x"0000" when x"11CB",
			x"0000" when x"11CC",
			x"0000" when x"11CD",
			x"0000" when x"11CE",
			x"0000" when x"11CF",
			x"0000" when x"11D0",
			x"0000" when x"11D1",
			x"0000" when x"11D2",
			x"0000" when x"11D3",
			x"0000" when x"11D4",
			x"0000" when x"11D5",
			x"0000" when x"11D6",
			x"0000" when x"11D7",
			x"0000" when x"11D8",
			x"0000" when x"11D9",
			x"0000" when x"11DA",
			x"0000" when x"11DB",
			x"0000" when x"11DC",
			x"0000" when x"11DD",
			x"0000" when x"11DE",
			x"0000" when x"11DF",
			x"0000" when x"11E0",
			x"0000" when x"11E1",
			x"0000" when x"11E2",
			x"0000" when x"11E3",
			x"0000" when x"11E4",
			x"0000" when x"11E5",
			x"0000" when x"11E6",
			x"0000" when x"11E7",
			x"0000" when x"11E8",
			x"0000" when x"11E9",
			x"0000" when x"11EA",
			x"0000" when x"11EB",
			x"0000" when x"11EC",
			x"0000" when x"11ED",
			x"0000" when x"11EE",
			x"0000" when x"11EF",
			x"0000" when x"11F0",
			x"0000" when x"11F1",
			x"0000" when x"11F2",
			x"0000" when x"11F3",
			x"0000" when x"11F4",
			x"0000" when x"11F5",
			x"0000" when x"11F6",
			x"0000" when x"11F7",
			x"0000" when x"11F8",
			x"0000" when x"11F9",
			x"0000" when x"11FA",
			x"0000" when x"11FB",
			x"0000" when x"11FC",
			x"0000" when x"11FD",
			x"0000" when x"11FE",
			x"0000" when x"11FF",
			x"0000" when x"1200",
			x"0000" when x"1201",
			x"0000" when x"1202",
			x"0000" when x"1203",
			x"0000" when x"1204",
			x"0000" when x"1205",
			x"0000" when x"1206",
			x"0000" when x"1207",
			x"0000" when x"1208",
			x"0000" when x"1209",
			x"0000" when x"120A",
			x"0000" when x"120B",
			x"0000" when x"120C",
			x"0000" when x"120D",
			x"0000" when x"120E",
			x"0000" when x"120F",
			x"0000" when x"1210",
			x"0000" when x"1211",
			x"0000" when x"1212",
			x"0000" when x"1213",
			x"0000" when x"1214",
			x"0000" when x"1215",
			x"0000" when x"1216",
			x"0000" when x"1217",
			x"0000" when x"1218",
			x"0000" when x"1219",
			x"0000" when x"121A",
			x"0000" when x"121B",
			x"0000" when x"121C",
			x"0000" when x"121D",
			x"0000" when x"121E",
			x"0000" when x"121F",
			x"0000" when x"1220",
			x"0000" when x"1221",
			x"0000" when x"1222",
			x"0000" when x"1223",
			x"0000" when x"1224",
			x"0000" when x"1225",
			x"0000" when x"1226",
			x"0000" when x"1227",
			x"0000" when x"1228",
			x"0000" when x"1229",
			x"0000" when x"122A",
			x"0000" when x"122B",
			x"0000" when x"122C",
			x"0000" when x"122D",
			x"0000" when x"122E",
			x"0000" when x"122F",
			x"0000" when x"1230",
			x"0000" when x"1231",
			x"0000" when x"1232",
			x"0000" when x"1233",
			x"0000" when x"1234",
			x"0000" when x"1235",
			x"0000" when x"1236",
			x"0000" when x"1237",
			x"0000" when x"1238",
			x"0000" when x"1239",
			x"0000" when x"123A",
			x"0000" when x"123B",
			x"0000" when x"123C",
			x"0000" when x"123D",
			x"0000" when x"123E",
			x"0000" when x"123F",
			x"0000" when x"1240",
			x"0000" when x"1241",
			x"0000" when x"1242",
			x"0000" when x"1243",
			x"0000" when x"1244",
			x"0000" when x"1245",
			x"0000" when x"1246",
			x"0000" when x"1247",
			x"0000" when x"1248",
			x"0000" when x"1249",
			x"0000" when x"124A",
			x"0000" when x"124B",
			x"0000" when x"124C",
			x"0000" when x"124D",
			x"0000" when x"124E",
			x"0000" when x"124F",
			x"0000" when x"1250",
			x"0000" when x"1251",
			x"0000" when x"1252",
			x"0000" when x"1253",
			x"0000" when x"1254",
			x"0000" when x"1255",
			x"0000" when x"1256",
			x"0000" when x"1257",
			x"0000" when x"1258",
			x"0000" when x"1259",
			x"0000" when x"125A",
			x"0000" when x"125B",
			x"0000" when x"125C",
			x"0000" when x"125D",
			x"0000" when x"125E",
			x"0000" when x"125F",
			x"0000" when x"1260",
			x"0000" when x"1261",
			x"0000" when x"1262",
			x"0000" when x"1263",
			x"0000" when x"1264",
			x"0000" when x"1265",
			x"0000" when x"1266",
			x"0000" when x"1267",
			x"0000" when x"1268",
			x"0000" when x"1269",
			x"0000" when x"126A",
			x"0000" when x"126B",
			x"0000" when x"126C",
			x"0000" when x"126D",
			x"0000" when x"126E",
			x"0000" when x"126F",
			x"0000" when x"1270",
			x"0000" when x"1271",
			x"0000" when x"1272",
			x"0000" when x"1273",
			x"0000" when x"1274",
			x"0000" when x"1275",
			x"0000" when x"1276",
			x"0000" when x"1277",
			x"0000" when x"1278",
			x"0000" when x"1279",
			x"0000" when x"127A",
			x"0000" when x"127B",
			x"0000" when x"127C",
			x"0000" when x"127D",
			x"0000" when x"127E",
			x"0000" when x"127F",
			x"0000" when x"1280",
			x"0000" when x"1281",
			x"0000" when x"1282",
			x"0000" when x"1283",
			x"0000" when x"1284",
			x"0000" when x"1285",
			x"0000" when x"1286",
			x"0000" when x"1287",
			x"0000" when x"1288",
			x"0000" when x"1289",
			x"0000" when x"128A",
			x"0000" when x"128B",
			x"0000" when x"128C",
			x"0000" when x"128D",
			x"0000" when x"128E",
			x"0000" when x"128F",
			x"0000" when x"1290",
			x"0000" when x"1291",
			x"0000" when x"1292",
			x"0000" when x"1293",
			x"0000" when x"1294",
			x"0000" when x"1295",
			x"0000" when x"1296",
			x"0000" when x"1297",
			x"0000" when x"1298",
			x"0000" when x"1299",
			x"0000" when x"129A",
			x"0000" when x"129B",
			x"0000" when x"129C",
			x"0000" when x"129D",
			x"0000" when x"129E",
			x"0000" when x"129F",
			x"0000" when x"12A0",
			x"0000" when x"12A1",
			x"0000" when x"12A2",
			x"0000" when x"12A3",
			x"0000" when x"12A4",
			x"0000" when x"12A5",
			x"0000" when x"12A6",
			x"0000" when x"12A7",
			x"0000" when x"12A8",
			x"0000" when x"12A9",
			x"0000" when x"12AA",
			x"0000" when x"12AB",
			x"0000" when x"12AC",
			x"0000" when x"12AD",
			x"0000" when x"12AE",
			x"0000" when x"12AF",
			x"0000" when x"12B0",
			x"0000" when x"12B1",
			x"0000" when x"12B2",
			x"0000" when x"12B3",
			x"0000" when x"12B4",
			x"0000" when x"12B5",
			x"0000" when x"12B6",
			x"0000" when x"12B7",
			x"0000" when x"12B8",
			x"0000" when x"12B9",
			x"0000" when x"12BA",
			x"0000" when x"12BB",
			x"0000" when x"12BC",
			x"0000" when x"12BD",
			x"0000" when x"12BE",
			x"0000" when x"12BF",
			x"0000" when x"12C0",
			x"0000" when x"12C1",
			x"0000" when x"12C2",
			x"0000" when x"12C3",
			x"0000" when x"12C4",
			x"0000" when x"12C5",
			x"0000" when x"12C6",
			x"0000" when x"12C7",
			x"0000" when x"12C8",
			x"0000" when x"12C9",
			x"0000" when x"12CA",
			x"0000" when x"12CB",
			x"0000" when x"12CC",
			x"0000" when x"12CD",
			x"0000" when x"12CE",
			x"0000" when x"12CF",
			x"0000" when x"12D0",
			x"0000" when x"12D1",
			x"0000" when x"12D2",
			x"0000" when x"12D3",
			x"0000" when x"12D4",
			x"0000" when x"12D5",
			x"0000" when x"12D6",
			x"0000" when x"12D7",
			x"0000" when x"12D8",
			x"0000" when x"12D9",
			x"0000" when x"12DA",
			x"0000" when x"12DB",
			x"0000" when x"12DC",
			x"0000" when x"12DD",
			x"0000" when x"12DE",
			x"0000" when x"12DF",
			x"0000" when x"12E0",
			x"0000" when x"12E1",
			x"0000" when x"12E2",
			x"0000" when x"12E3",
			x"0000" when x"12E4",
			x"0000" when x"12E5",
			x"0000" when x"12E6",
			x"0000" when x"12E7",
			x"0000" when x"12E8",
			x"0000" when x"12E9",
			x"0000" when x"12EA",
			x"0000" when x"12EB",
			x"0000" when x"12EC",
			x"0000" when x"12ED",
			x"0000" when x"12EE",
			x"0000" when x"12EF",
			x"0000" when x"12F0",
			x"0000" when x"12F1",
			x"0000" when x"12F2",
			x"0000" when x"12F3",
			x"0000" when x"12F4",
			x"0000" when x"12F5",
			x"0000" when x"12F6",
			x"0000" when x"12F7",
			x"0000" when x"12F8",
			x"0000" when x"12F9",
			x"0000" when x"12FA",
			x"0000" when x"12FB",
			x"0000" when x"12FC",
			x"0000" when x"12FD",
			x"0000" when x"12FE",
			x"0000" when x"12FF",
			x"0000" when x"1300",
			x"0000" when x"1301",
			x"0000" when x"1302",
			x"0000" when x"1303",
			x"0000" when x"1304",
			x"0000" when x"1305",
			x"0000" when x"1306",
			x"0000" when x"1307",
			x"0000" when x"1308",
			x"0000" when x"1309",
			x"0000" when x"130A",
			x"0000" when x"130B",
			x"0000" when x"130C",
			x"0000" when x"130D",
			x"0000" when x"130E",
			x"0000" when x"130F",
			x"0000" when x"1310",
			x"0000" when x"1311",
			x"0000" when x"1312",
			x"0000" when x"1313",
			x"0000" when x"1314",
			x"0000" when x"1315",
			x"0000" when x"1316",
			x"0000" when x"1317",
			x"0000" when x"1318",
			x"0000" when x"1319",
			x"0000" when x"131A",
			x"0000" when x"131B",
			x"0000" when x"131C",
			x"0000" when x"131D",
			x"0000" when x"131E",
			x"0000" when x"131F",
			x"0000" when x"1320",
			x"0000" when x"1321",
			x"0000" when x"1322",
			x"0000" when x"1323",
			x"0000" when x"1324",
			x"0000" when x"1325",
			x"0000" when x"1326",
			x"0000" when x"1327",
			x"0000" when x"1328",
			x"0000" when x"1329",
			x"0000" when x"132A",
			x"0000" when x"132B",
			x"0000" when x"132C",
			x"0000" when x"132D",
			x"0000" when x"132E",
			x"0000" when x"132F",
			x"0000" when x"1330",
			x"0000" when x"1331",
			x"0000" when x"1332",
			x"0000" when x"1333",
			x"0000" when x"1334",
			x"0000" when x"1335",
			x"0000" when x"1336",
			x"0000" when x"1337",
			x"0000" when x"1338",
			x"0000" when x"1339",
			x"0000" when x"133A",
			x"0000" when x"133B",
			x"0000" when x"133C",
			x"0000" when x"133D",
			x"0000" when x"133E",
			x"0000" when x"133F",
			x"0000" when x"1340",
			x"0000" when x"1341",
			x"0000" when x"1342",
			x"0000" when x"1343",
			x"0000" when x"1344",
			x"0000" when x"1345",
			x"0000" when x"1346",
			x"0000" when x"1347",
			x"0000" when x"1348",
			x"0000" when x"1349",
			x"0000" when x"134A",
			x"0000" when x"134B",
			x"0000" when x"134C",
			x"0000" when x"134D",
			x"0000" when x"134E",
			x"0000" when x"134F",
			x"0000" when x"1350",
			x"0000" when x"1351",
			x"0000" when x"1352",
			x"0000" when x"1353",
			x"0000" when x"1354",
			x"0000" when x"1355",
			x"0000" when x"1356",
			x"0000" when x"1357",
			x"0000" when x"1358",
			x"0000" when x"1359",
			x"0000" when x"135A",
			x"0000" when x"135B",
			x"0000" when x"135C",
			x"0000" when x"135D",
			x"0000" when x"135E",
			x"0000" when x"135F",
			x"0000" when x"1360",
			x"0000" when x"1361",
			x"0000" when x"1362",
			x"0000" when x"1363",
			x"0000" when x"1364",
			x"0000" when x"1365",
			x"0000" when x"1366",
			x"0000" when x"1367",
			x"0000" when x"1368",
			x"0000" when x"1369",
			x"0000" when x"136A",
			x"0000" when x"136B",
			x"0000" when x"136C",
			x"0000" when x"136D",
			x"0000" when x"136E",
			x"0000" when x"136F",
			x"0000" when x"1370",
			x"0000" when x"1371",
			x"0000" when x"1372",
			x"0000" when x"1373",
			x"0000" when x"1374",
			x"0000" when x"1375",
			x"0000" when x"1376",
			x"0000" when x"1377",
			x"0000" when x"1378",
			x"0000" when x"1379",
			x"0000" when x"137A",
			x"0000" when x"137B",
			x"0000" when x"137C",
			x"0000" when x"137D",
			x"0000" when x"137E",
			x"0000" when x"137F",
			x"0000" when x"1380",
			x"0000" when x"1381",
			x"0000" when x"1382",
			x"0000" when x"1383",
			x"0000" when x"1384",
			x"0000" when x"1385",
			x"0000" when x"1386",
			x"0000" when x"1387",
			x"0000" when x"1388",
			x"0000" when x"1389",
			x"0000" when x"138A",
			x"0000" when x"138B",
			x"0000" when x"138C",
			x"0000" when x"138D",
			x"0000" when x"138E",
			x"0000" when x"138F",
			x"0000" when x"1390",
			x"0000" when x"1391",
			x"0000" when x"1392",
			x"0000" when x"1393",
			x"0000" when x"1394",
			x"0000" when x"1395",
			x"0000" when x"1396",
			x"0000" when x"1397",
			x"0000" when x"1398",
			x"0000" when x"1399",
			x"0000" when x"139A",
			x"0000" when x"139B",
			x"0000" when x"139C",
			x"0000" when x"139D",
			x"0000" when x"139E",
			x"0000" when x"139F",
			x"0000" when x"13A0",
			x"0000" when x"13A1",
			x"0000" when x"13A2",
			x"0000" when x"13A3",
			x"0000" when x"13A4",
			x"0000" when x"13A5",
			x"0000" when x"13A6",
			x"0000" when x"13A7",
			x"0000" when x"13A8",
			x"0000" when x"13A9",
			x"0000" when x"13AA",
			x"0000" when x"13AB",
			x"0000" when x"13AC",
			x"0000" when x"13AD",
			x"0000" when x"13AE",
			x"0000" when x"13AF",
			x"0000" when x"13B0",
			x"0000" when x"13B1",
			x"0000" when x"13B2",
			x"0000" when x"13B3",
			x"0000" when x"13B4",
			x"0000" when x"13B5",
			x"0000" when x"13B6",
			x"0000" when x"13B7",
			x"0000" when x"13B8",
			x"0000" when x"13B9",
			x"0000" when x"13BA",
			x"0000" when x"13BB",
			x"0000" when x"13BC",
			x"0000" when x"13BD",
			x"0000" when x"13BE",
			x"0000" when x"13BF",
			x"0000" when x"13C0",
			x"0000" when x"13C1",
			x"0000" when x"13C2",
			x"0000" when x"13C3",
			x"0000" when x"13C4",
			x"0000" when x"13C5",
			x"0000" when x"13C6",
			x"0000" when x"13C7",
			x"0000" when x"13C8",
			x"0000" when x"13C9",
			x"0000" when x"13CA",
			x"0000" when x"13CB",
			x"0000" when x"13CC",
			x"0000" when x"13CD",
			x"0000" when x"13CE",
			x"0000" when x"13CF",
			x"0000" when x"13D0",
			x"0000" when x"13D1",
			x"0000" when x"13D2",
			x"0000" when x"13D3",
			x"0000" when x"13D4",
			x"0000" when x"13D5",
			x"0000" when x"13D6",
			x"0000" when x"13D7",
			x"0000" when x"13D8",
			x"0000" when x"13D9",
			x"0000" when x"13DA",
			x"0000" when x"13DB",
			x"0000" when x"13DC",
			x"0000" when x"13DD",
			x"0000" when x"13DE",
			x"0000" when x"13DF",
			x"0000" when x"13E0",
			x"0000" when x"13E1",
			x"0000" when x"13E2",
			x"0000" when x"13E3",
			x"0000" when x"13E4",
			x"0000" when x"13E5",
			x"0000" when x"13E6",
			x"0000" when x"13E7",
			x"0000" when x"13E8",
			x"0000" when x"13E9",
			x"0000" when x"13EA",
			x"0000" when x"13EB",
			x"0000" when x"13EC",
			x"0000" when x"13ED",
			x"0000" when x"13EE",
			x"0000" when x"13EF",
			x"0000" when x"13F0",
			x"0000" when x"13F1",
			x"0000" when x"13F2",
			x"0000" when x"13F3",
			x"0000" when x"13F4",
			x"0000" when x"13F5",
			x"0000" when x"13F6",
			x"0000" when x"13F7",
			x"0000" when x"13F8",
			x"0000" when x"13F9",
			x"0000" when x"13FA",
			x"0000" when x"13FB",
			x"0000" when x"13FC",
			x"0000" when x"13FD",
			x"0000" when x"13FE",
			x"0000" when x"13FF",
			x"0000" when x"1400",
			x"0000" when x"1401",
			x"0000" when x"1402",
			x"0000" when x"1403",
			x"0000" when x"1404",
			x"0000" when x"1405",
			x"0000" when x"1406",
			x"0000" when x"1407",
			x"0000" when x"1408",
			x"0000" when x"1409",
			x"0000" when x"140A",
			x"0000" when x"140B",
			x"0000" when x"140C",
			x"0000" when x"140D",
			x"0000" when x"140E",
			x"0000" when x"140F",
			x"0000" when x"1410",
			x"0000" when x"1411",
			x"0000" when x"1412",
			x"0000" when x"1413",
			x"0000" when x"1414",
			x"0000" when x"1415",
			x"0000" when x"1416",
			x"0000" when x"1417",
			x"0000" when x"1418",
			x"0000" when x"1419",
			x"0000" when x"141A",
			x"0000" when x"141B",
			x"0000" when x"141C",
			x"0000" when x"141D",
			x"0000" when x"141E",
			x"0000" when x"141F",
			x"0000" when x"1420",
			x"0000" when x"1421",
			x"0000" when x"1422",
			x"0000" when x"1423",
			x"0000" when x"1424",
			x"0000" when x"1425",
			x"0000" when x"1426",
			x"0000" when x"1427",
			x"0000" when x"1428",
			x"0000" when x"1429",
			x"0000" when x"142A",
			x"0000" when x"142B",
			x"0000" when x"142C",
			x"0000" when x"142D",
			x"0000" when x"142E",
			x"0000" when x"142F",
			x"0000" when x"1430",
			x"0000" when x"1431",
			x"0000" when x"1432",
			x"0000" when x"1433",
			x"0000" when x"1434",
			x"0000" when x"1435",
			x"0000" when x"1436",
			x"0000" when x"1437",
			x"0000" when x"1438",
			x"0000" when x"1439",
			x"0000" when x"143A",
			x"0000" when x"143B",
			x"0000" when x"143C",
			x"0000" when x"143D",
			x"0000" when x"143E",
			x"0000" when x"143F",
			x"0000" when x"1440",
			x"0000" when x"1441",
			x"0000" when x"1442",
			x"0000" when x"1443",
			x"0000" when x"1444",
			x"0000" when x"1445",
			x"0000" when x"1446",
			x"0000" when x"1447",
			x"0000" when x"1448",
			x"0000" when x"1449",
			x"0000" when x"144A",
			x"0000" when x"144B",
			x"0000" when x"144C",
			x"0000" when x"144D",
			x"0000" when x"144E",
			x"0000" when x"144F",
			x"0000" when x"1450",
			x"0000" when x"1451",
			x"0000" when x"1452",
			x"0000" when x"1453",
			x"0000" when x"1454",
			x"0000" when x"1455",
			x"0000" when x"1456",
			x"0000" when x"1457",
			x"0000" when x"1458",
			x"0000" when x"1459",
			x"0000" when x"145A",
			x"0000" when x"145B",
			x"0000" when x"145C",
			x"0000" when x"145D",
			x"0000" when x"145E",
			x"0000" when x"145F",
			x"0000" when x"1460",
			x"0000" when x"1461",
			x"0000" when x"1462",
			x"0000" when x"1463",
			x"0000" when x"1464",
			x"0000" when x"1465",
			x"0000" when x"1466",
			x"0000" when x"1467",
			x"0000" when x"1468",
			x"0000" when x"1469",
			x"0000" when x"146A",
			x"0000" when x"146B",
			x"0000" when x"146C",
			x"0000" when x"146D",
			x"0000" when x"146E",
			x"0000" when x"146F",
			x"0000" when x"1470",
			x"0000" when x"1471",
			x"0000" when x"1472",
			x"0000" when x"1473",
			x"0000" when x"1474",
			x"0000" when x"1475",
			x"0000" when x"1476",
			x"0000" when x"1477",
			x"0000" when x"1478",
			x"0000" when x"1479",
			x"0000" when x"147A",
			x"0000" when x"147B",
			x"0000" when x"147C",
			x"0000" when x"147D",
			x"0000" when x"147E",
			x"0000" when x"147F",
			x"0000" when x"1480",
			x"0000" when x"1481",
			x"0000" when x"1482",
			x"0000" when x"1483",
			x"0000" when x"1484",
			x"0000" when x"1485",
			x"0000" when x"1486",
			x"0000" when x"1487",
			x"0000" when x"1488",
			x"0000" when x"1489",
			x"0000" when x"148A",
			x"0000" when x"148B",
			x"0000" when x"148C",
			x"0000" when x"148D",
			x"0000" when x"148E",
			x"0000" when x"148F",
			x"0000" when x"1490",
			x"0000" when x"1491",
			x"0000" when x"1492",
			x"0000" when x"1493",
			x"0000" when x"1494",
			x"0000" when x"1495",
			x"0000" when x"1496",
			x"0000" when x"1497",
			x"0000" when x"1498",
			x"0000" when x"1499",
			x"0000" when x"149A",
			x"0000" when x"149B",
			x"0000" when x"149C",
			x"0000" when x"149D",
			x"0000" when x"149E",
			x"0000" when x"149F",
			x"0000" when x"14A0",
			x"0000" when x"14A1",
			x"0000" when x"14A2",
			x"0000" when x"14A3",
			x"0000" when x"14A4",
			x"0000" when x"14A5",
			x"0000" when x"14A6",
			x"0000" when x"14A7",
			x"0000" when x"14A8",
			x"0000" when x"14A9",
			x"0000" when x"14AA",
			x"0000" when x"14AB",
			x"0000" when x"14AC",
			x"0000" when x"14AD",
			x"0000" when x"14AE",
			x"0000" when x"14AF",
			x"0000" when x"14B0",
			x"0000" when x"14B1",
			x"0000" when x"14B2",
			x"0000" when x"14B3",
			x"0000" when x"14B4",
			x"0000" when x"14B5",
			x"0000" when x"14B6",
			x"0000" when x"14B7",
			x"0000" when x"14B8",
			x"0000" when x"14B9",
			x"0000" when x"14BA",
			x"0000" when x"14BB",
			x"0000" when x"14BC",
			x"0000" when x"14BD",
			x"0000" when x"14BE",
			x"0000" when x"14BF",
			x"0000" when x"14C0",
			x"0000" when x"14C1",
			x"0000" when x"14C2",
			x"0000" when x"14C3",
			x"0000" when x"14C4",
			x"0000" when x"14C5",
			x"0000" when x"14C6",
			x"0000" when x"14C7",
			x"0000" when x"14C8",
			x"0000" when x"14C9",
			x"0000" when x"14CA",
			x"0000" when x"14CB",
			x"0000" when x"14CC",
			x"0000" when x"14CD",
			x"0000" when x"14CE",
			x"0000" when x"14CF",
			x"0000" when x"14D0",
			x"0000" when x"14D1",
			x"0000" when x"14D2",
			x"0000" when x"14D3",
			x"0000" when x"14D4",
			x"0000" when x"14D5",
			x"0000" when x"14D6",
			x"0000" when x"14D7",
			x"0000" when x"14D8",
			x"0000" when x"14D9",
			x"0000" when x"14DA",
			x"0000" when x"14DB",
			x"0000" when x"14DC",
			x"0000" when x"14DD",
			x"0000" when x"14DE",
			x"0000" when x"14DF",
			x"0000" when x"14E0",
			x"0000" when x"14E1",
			x"0000" when x"14E2",
			x"0000" when x"14E3",
			x"0000" when x"14E4",
			x"0000" when x"14E5",
			x"0000" when x"14E6",
			x"0000" when x"14E7",
			x"0000" when x"14E8",
			x"0000" when x"14E9",
			x"0000" when x"14EA",
			x"0000" when x"14EB",
			x"0000" when x"14EC",
			x"0000" when x"14ED",
			x"0000" when x"14EE",
			x"0000" when x"14EF",
			x"0000" when x"14F0",
			x"0000" when x"14F1",
			x"0000" when x"14F2",
			x"0000" when x"14F3",
			x"0000" when x"14F4",
			x"0000" when x"14F5",
			x"0000" when x"14F6",
			x"0000" when x"14F7",
			x"0000" when x"14F8",
			x"0000" when x"14F9",
			x"0000" when x"14FA",
			x"0000" when x"14FB",
			x"0000" when x"14FC",
			x"0000" when x"14FD",
			x"0000" when x"14FE",
			x"0000" when x"14FF",
			x"0000" when x"1500",
			x"0000" when x"1501",
			x"0000" when x"1502",
			x"0000" when x"1503",
			x"0000" when x"1504",
			x"0000" when x"1505",
			x"0000" when x"1506",
			x"0000" when x"1507",
			x"0000" when x"1508",
			x"0000" when x"1509",
			x"0000" when x"150A",
			x"0000" when x"150B",
			x"0000" when x"150C",
			x"0000" when x"150D",
			x"0000" when x"150E",
			x"0000" when x"150F",
			x"0000" when x"1510",
			x"0000" when x"1511",
			x"0000" when x"1512",
			x"0000" when x"1513",
			x"0000" when x"1514",
			x"0000" when x"1515",
			x"0000" when x"1516",
			x"0000" when x"1517",
			x"0000" when x"1518",
			x"0000" when x"1519",
			x"0000" when x"151A",
			x"0000" when x"151B",
			x"0000" when x"151C",
			x"0000" when x"151D",
			x"0000" when x"151E",
			x"0000" when x"151F",
			x"0000" when x"1520",
			x"0000" when x"1521",
			x"0000" when x"1522",
			x"0000" when x"1523",
			x"0000" when x"1524",
			x"0000" when x"1525",
			x"0000" when x"1526",
			x"0000" when x"1527",
			x"0000" when x"1528",
			x"0000" when x"1529",
			x"0000" when x"152A",
			x"0000" when x"152B",
			x"0000" when x"152C",
			x"0000" when x"152D",
			x"0000" when x"152E",
			x"0000" when x"152F",
			x"0000" when x"1530",
			x"0000" when x"1531",
			x"0000" when x"1532",
			x"0000" when x"1533",
			x"0000" when x"1534",
			x"0000" when x"1535",
			x"0000" when x"1536",
			x"0000" when x"1537",
			x"0000" when x"1538",
			x"0000" when x"1539",
			x"0000" when x"153A",
			x"0000" when x"153B",
			x"0000" when x"153C",
			x"0000" when x"153D",
			x"0000" when x"153E",
			x"0000" when x"153F",
			x"0000" when x"1540",
			x"0000" when x"1541",
			x"0000" when x"1542",
			x"0000" when x"1543",
			x"0000" when x"1544",
			x"0000" when x"1545",
			x"0000" when x"1546",
			x"0000" when x"1547",
			x"0000" when x"1548",
			x"0000" when x"1549",
			x"0000" when x"154A",
			x"0000" when x"154B",
			x"0000" when x"154C",
			x"0000" when x"154D",
			x"0000" when x"154E",
			x"0000" when x"154F",
			x"0000" when x"1550",
			x"0000" when x"1551",
			x"0000" when x"1552",
			x"0000" when x"1553",
			x"0000" when x"1554",
			x"0000" when x"1555",
			x"0000" when x"1556",
			x"0000" when x"1557",
			x"0000" when x"1558",
			x"0000" when x"1559",
			x"0000" when x"155A",
			x"0000" when x"155B",
			x"0000" when x"155C",
			x"0000" when x"155D",
			x"0000" when x"155E",
			x"0000" when x"155F",
			x"0000" when x"1560",
			x"0000" when x"1561",
			x"0000" when x"1562",
			x"0000" when x"1563",
			x"0000" when x"1564",
			x"0000" when x"1565",
			x"0000" when x"1566",
			x"0000" when x"1567",
			x"0000" when x"1568",
			x"0000" when x"1569",
			x"0000" when x"156A",
			x"0000" when x"156B",
			x"0000" when x"156C",
			x"0000" when x"156D",
			x"0000" when x"156E",
			x"0000" when x"156F",
			x"0000" when x"1570",
			x"0000" when x"1571",
			x"0000" when x"1572",
			x"0000" when x"1573",
			x"0000" when x"1574",
			x"0000" when x"1575",
			x"0000" when x"1576",
			x"0000" when x"1577",
			x"0000" when x"1578",
			x"0000" when x"1579",
			x"0000" when x"157A",
			x"0000" when x"157B",
			x"0000" when x"157C",
			x"0000" when x"157D",
			x"0000" when x"157E",
			x"0000" when x"157F",
			x"0000" when x"1580",
			x"0000" when x"1581",
			x"0000" when x"1582",
			x"0000" when x"1583",
			x"0000" when x"1584",
			x"0000" when x"1585",
			x"0000" when x"1586",
			x"0000" when x"1587",
			x"0000" when x"1588",
			x"0000" when x"1589",
			x"0000" when x"158A",
			x"0000" when x"158B",
			x"0000" when x"158C",
			x"0000" when x"158D",
			x"0000" when x"158E",
			x"0000" when x"158F",
			x"0000" when x"1590",
			x"0000" when x"1591",
			x"0000" when x"1592",
			x"0000" when x"1593",
			x"0000" when x"1594",
			x"0000" when x"1595",
			x"0000" when x"1596",
			x"0000" when x"1597",
			x"0000" when x"1598",
			x"0000" when x"1599",
			x"0000" when x"159A",
			x"0000" when x"159B",
			x"0000" when x"159C",
			x"0000" when x"159D",
			x"0000" when x"159E",
			x"0000" when x"159F",
			x"0000" when x"15A0",
			x"0000" when x"15A1",
			x"0000" when x"15A2",
			x"0000" when x"15A3",
			x"0000" when x"15A4",
			x"0000" when x"15A5",
			x"0000" when x"15A6",
			x"0000" when x"15A7",
			x"0000" when x"15A8",
			x"0000" when x"15A9",
			x"0000" when x"15AA",
			x"0000" when x"15AB",
			x"0000" when x"15AC",
			x"0000" when x"15AD",
			x"0000" when x"15AE",
			x"0000" when x"15AF",
			x"0000" when x"15B0",
			x"0000" when x"15B1",
			x"0000" when x"15B2",
			x"0000" when x"15B3",
			x"0000" when x"15B4",
			x"0000" when x"15B5",
			x"0000" when x"15B6",
			x"0000" when x"15B7",
			x"0000" when x"15B8",
			x"0000" when x"15B9",
			x"0000" when x"15BA",
			x"0000" when x"15BB",
			x"0000" when x"15BC",
			x"0000" when x"15BD",
			x"0000" when x"15BE",
			x"0000" when x"15BF",
			x"0000" when x"15C0",
			x"0000" when x"15C1",
			x"0000" when x"15C2",
			x"0000" when x"15C3",
			x"0000" when x"15C4",
			x"0000" when x"15C5",
			x"0000" when x"15C6",
			x"0000" when x"15C7",
			x"0000" when x"15C8",
			x"0000" when x"15C9",
			x"0000" when x"15CA",
			x"0000" when x"15CB",
			x"0000" when x"15CC",
			x"0000" when x"15CD",
			x"0000" when x"15CE",
			x"0000" when x"15CF",
			x"0000" when x"15D0",
			x"0000" when x"15D1",
			x"0000" when x"15D2",
			x"0000" when x"15D3",
			x"0000" when x"15D4",
			x"0000" when x"15D5",
			x"0000" when x"15D6",
			x"0000" when x"15D7",
			x"0000" when x"15D8",
			x"0000" when x"15D9",
			x"0000" when x"15DA",
			x"0000" when x"15DB",
			x"0000" when x"15DC",
			x"0000" when x"15DD",
			x"0000" when x"15DE",
			x"0000" when x"15DF",
			x"0000" when x"15E0",
			x"0000" when x"15E1",
			x"0000" when x"15E2",
			x"0000" when x"15E3",
			x"0000" when x"15E4",
			x"0000" when x"15E5",
			x"0000" when x"15E6",
			x"0000" when x"15E7",
			x"0000" when x"15E8",
			x"0000" when x"15E9",
			x"0000" when x"15EA",
			x"0000" when x"15EB",
			x"0000" when x"15EC",
			x"0000" when x"15ED",
			x"0000" when x"15EE",
			x"0000" when x"15EF",
			x"0000" when x"15F0",
			x"0000" when x"15F1",
			x"0000" when x"15F2",
			x"0000" when x"15F3",
			x"0000" when x"15F4",
			x"0000" when x"15F5",
			x"0000" when x"15F6",
			x"0000" when x"15F7",
			x"0000" when x"15F8",
			x"0000" when x"15F9",
			x"0000" when x"15FA",
			x"0000" when x"15FB",
			x"0000" when x"15FC",
			x"0000" when x"15FD",
			x"0000" when x"15FE",
			x"0000" when x"15FF",
			x"0000" when x"1600",
			x"0000" when x"1601",
			x"0000" when x"1602",
			x"0000" when x"1603",
			x"0000" when x"1604",
			x"0000" when x"1605",
			x"0000" when x"1606",
			x"0000" when x"1607",
			x"0000" when x"1608",
			x"0000" when x"1609",
			x"0000" when x"160A",
			x"0000" when x"160B",
			x"0000" when x"160C",
			x"0000" when x"160D",
			x"0000" when x"160E",
			x"0000" when x"160F",
			x"0000" when x"1610",
			x"0000" when x"1611",
			x"0000" when x"1612",
			x"0000" when x"1613",
			x"0000" when x"1614",
			x"0000" when x"1615",
			x"0000" when x"1616",
			x"0000" when x"1617",
			x"0000" when x"1618",
			x"0000" when x"1619",
			x"0000" when x"161A",
			x"0000" when x"161B",
			x"0000" when x"161C",
			x"0000" when x"161D",
			x"0000" when x"161E",
			x"0000" when x"161F",
			x"0000" when x"1620",
			x"0000" when x"1621",
			x"0000" when x"1622",
			x"0000" when x"1623",
			x"0000" when x"1624",
			x"0000" when x"1625",
			x"0000" when x"1626",
			x"0000" when x"1627",
			x"0000" when x"1628",
			x"0000" when x"1629",
			x"0000" when x"162A",
			x"0000" when x"162B",
			x"0000" when x"162C",
			x"0000" when x"162D",
			x"0000" when x"162E",
			x"0000" when x"162F",
			x"0000" when x"1630",
			x"0000" when x"1631",
			x"0000" when x"1632",
			x"0000" when x"1633",
			x"0000" when x"1634",
			x"0000" when x"1635",
			x"0000" when x"1636",
			x"0000" when x"1637",
			x"0000" when x"1638",
			x"0000" when x"1639",
			x"0000" when x"163A",
			x"0000" when x"163B",
			x"0000" when x"163C",
			x"0000" when x"163D",
			x"0000" when x"163E",
			x"0000" when x"163F",
			x"0000" when x"1640",
			x"0000" when x"1641",
			x"0000" when x"1642",
			x"0000" when x"1643",
			x"0000" when x"1644",
			x"0000" when x"1645",
			x"0000" when x"1646",
			x"0000" when x"1647",
			x"0000" when x"1648",
			x"0000" when x"1649",
			x"0000" when x"164A",
			x"0000" when x"164B",
			x"0000" when x"164C",
			x"0000" when x"164D",
			x"0000" when x"164E",
			x"0000" when x"164F",
			x"0000" when x"1650",
			x"0000" when x"1651",
			x"0000" when x"1652",
			x"0000" when x"1653",
			x"0000" when x"1654",
			x"0000" when x"1655",
			x"0000" when x"1656",
			x"0000" when x"1657",
			x"0000" when x"1658",
			x"0000" when x"1659",
			x"0000" when x"165A",
			x"0000" when x"165B",
			x"0000" when x"165C",
			x"0000" when x"165D",
			x"0000" when x"165E",
			x"0000" when x"165F",
			x"0000" when x"1660",
			x"0000" when x"1661",
			x"0000" when x"1662",
			x"0000" when x"1663",
			x"0000" when x"1664",
			x"0000" when x"1665",
			x"0000" when x"1666",
			x"0000" when x"1667",
			x"0000" when x"1668",
			x"0000" when x"1669",
			x"0000" when x"166A",
			x"0000" when x"166B",
			x"0000" when x"166C",
			x"0000" when x"166D",
			x"0000" when x"166E",
			x"0000" when x"166F",
			x"0000" when x"1670",
			x"0000" when x"1671",
			x"0000" when x"1672",
			x"0000" when x"1673",
			x"0000" when x"1674",
			x"0000" when x"1675",
			x"0000" when x"1676",
			x"0000" when x"1677",
			x"0000" when x"1678",
			x"0000" when x"1679",
			x"0000" when x"167A",
			x"0000" when x"167B",
			x"0000" when x"167C",
			x"0000" when x"167D",
			x"0000" when x"167E",
			x"0000" when x"167F",
			x"0000" when x"1680",
			x"0000" when x"1681",
			x"0000" when x"1682",
			x"0000" when x"1683",
			x"0000" when x"1684",
			x"0000" when x"1685",
			x"0000" when x"1686",
			x"0000" when x"1687",
			x"0000" when x"1688",
			x"0000" when x"1689",
			x"0000" when x"168A",
			x"0000" when x"168B",
			x"0000" when x"168C",
			x"0000" when x"168D",
			x"0000" when x"168E",
			x"0000" when x"168F",
			x"0000" when x"1690",
			x"0000" when x"1691",
			x"0000" when x"1692",
			x"0000" when x"1693",
			x"0000" when x"1694",
			x"0000" when x"1695",
			x"0000" when x"1696",
			x"0000" when x"1697",
			x"0000" when x"1698",
			x"0000" when x"1699",
			x"0000" when x"169A",
			x"0000" when x"169B",
			x"0000" when x"169C",
			x"0000" when x"169D",
			x"0000" when x"169E",
			x"0000" when x"169F",
			x"0000" when x"16A0",
			x"0000" when x"16A1",
			x"0000" when x"16A2",
			x"0000" when x"16A3",
			x"0000" when x"16A4",
			x"0000" when x"16A5",
			x"0000" when x"16A6",
			x"0000" when x"16A7",
			x"0000" when x"16A8",
			x"0000" when x"16A9",
			x"0000" when x"16AA",
			x"0000" when x"16AB",
			x"0000" when x"16AC",
			x"0000" when x"16AD",
			x"0000" when x"16AE",
			x"0000" when x"16AF",
			x"0000" when x"16B0",
			x"0000" when x"16B1",
			x"0000" when x"16B2",
			x"0000" when x"16B3",
			x"0000" when x"16B4",
			x"0000" when x"16B5",
			x"0000" when x"16B6",
			x"0000" when x"16B7",
			x"0000" when x"16B8",
			x"0000" when x"16B9",
			x"0000" when x"16BA",
			x"0000" when x"16BB",
			x"0000" when x"16BC",
			x"0000" when x"16BD",
			x"0000" when x"16BE",
			x"0000" when x"16BF",
			x"0000" when x"16C0",
			x"0000" when x"16C1",
			x"0000" when x"16C2",
			x"0000" when x"16C3",
			x"0000" when x"16C4",
			x"0000" when x"16C5",
			x"0000" when x"16C6",
			x"0000" when x"16C7",
			x"0000" when x"16C8",
			x"0000" when x"16C9",
			x"0000" when x"16CA",
			x"0000" when x"16CB",
			x"0000" when x"16CC",
			x"0000" when x"16CD",
			x"0000" when x"16CE",
			x"0000" when x"16CF",
			x"0000" when x"16D0",
			x"0000" when x"16D1",
			x"0000" when x"16D2",
			x"0000" when x"16D3",
			x"0000" when x"16D4",
			x"0000" when x"16D5",
			x"0000" when x"16D6",
			x"0000" when x"16D7",
			x"0000" when x"16D8",
			x"0000" when x"16D9",
			x"0000" when x"16DA",
			x"0000" when x"16DB",
			x"0000" when x"16DC",
			x"0000" when x"16DD",
			x"0000" when x"16DE",
			x"0000" when x"16DF",
			x"0000" when x"16E0",
			x"0000" when x"16E1",
			x"0000" when x"16E2",
			x"0000" when x"16E3",
			x"0000" when x"16E4",
			x"0000" when x"16E5",
			x"0000" when x"16E6",
			x"0000" when x"16E7",
			x"0000" when x"16E8",
			x"0000" when x"16E9",
			x"0000" when x"16EA",
			x"0000" when x"16EB",
			x"0000" when x"16EC",
			x"0000" when x"16ED",
			x"0000" when x"16EE",
			x"0000" when x"16EF",
			x"0000" when x"16F0",
			x"0000" when x"16F1",
			x"0000" when x"16F2",
			x"0000" when x"16F3",
			x"0000" when x"16F4",
			x"0000" when x"16F5",
			x"0000" when x"16F6",
			x"0000" when x"16F7",
			x"0000" when x"16F8",
			x"0000" when x"16F9",
			x"0000" when x"16FA",
			x"0000" when x"16FB",
			x"0000" when x"16FC",
			x"0000" when x"16FD",
			x"0000" when x"16FE",
			x"0000" when x"16FF",
			x"0000" when x"1700",
			x"0000" when x"1701",
			x"0000" when x"1702",
			x"0000" when x"1703",
			x"0000" when x"1704",
			x"0000" when x"1705",
			x"0000" when x"1706",
			x"0000" when x"1707",
			x"0000" when x"1708",
			x"0000" when x"1709",
			x"0000" when x"170A",
			x"0000" when x"170B",
			x"0000" when x"170C",
			x"0000" when x"170D",
			x"0000" when x"170E",
			x"0000" when x"170F",
			x"0000" when x"1710",
			x"0000" when x"1711",
			x"0000" when x"1712",
			x"0000" when x"1713",
			x"0000" when x"1714",
			x"0000" when x"1715",
			x"0000" when x"1716",
			x"0000" when x"1717",
			x"0000" when x"1718",
			x"0000" when x"1719",
			x"0000" when x"171A",
			x"0000" when x"171B",
			x"0000" when x"171C",
			x"0000" when x"171D",
			x"0000" when x"171E",
			x"0000" when x"171F",
			x"0000" when x"1720",
			x"0000" when x"1721",
			x"0000" when x"1722",
			x"0000" when x"1723",
			x"0000" when x"1724",
			x"0000" when x"1725",
			x"0000" when x"1726",
			x"0000" when x"1727",
			x"0000" when x"1728",
			x"0000" when x"1729",
			x"0000" when x"172A",
			x"0000" when x"172B",
			x"0000" when x"172C",
			x"0000" when x"172D",
			x"0000" when x"172E",
			x"0000" when x"172F",
			x"0000" when x"1730",
			x"0000" when x"1731",
			x"0000" when x"1732",
			x"0000" when x"1733",
			x"0000" when x"1734",
			x"0000" when x"1735",
			x"0000" when x"1736",
			x"0000" when x"1737",
			x"0000" when x"1738",
			x"0000" when x"1739",
			x"0000" when x"173A",
			x"0000" when x"173B",
			x"0000" when x"173C",
			x"0000" when x"173D",
			x"0000" when x"173E",
			x"0000" when x"173F",
			x"0000" when x"1740",
			x"0000" when x"1741",
			x"0000" when x"1742",
			x"0000" when x"1743",
			x"0000" when x"1744",
			x"0000" when x"1745",
			x"0000" when x"1746",
			x"0000" when x"1747",
			x"0000" when x"1748",
			x"0000" when x"1749",
			x"0000" when x"174A",
			x"0000" when x"174B",
			x"0000" when x"174C",
			x"0000" when x"174D",
			x"0000" when x"174E",
			x"0000" when x"174F",
			x"0000" when x"1750",
			x"0000" when x"1751",
			x"0000" when x"1752",
			x"0000" when x"1753",
			x"0000" when x"1754",
			x"0000" when x"1755",
			x"0000" when x"1756",
			x"0000" when x"1757",
			x"0000" when x"1758",
			x"0000" when x"1759",
			x"0000" when x"175A",
			x"0000" when x"175B",
			x"0000" when x"175C",
			x"0000" when x"175D",
			x"0000" when x"175E",
			x"0000" when x"175F",
			x"0000" when x"1760",
			x"0000" when x"1761",
			x"0000" when x"1762",
			x"0000" when x"1763",
			x"0000" when x"1764",
			x"0000" when x"1765",
			x"0000" when x"1766",
			x"0000" when x"1767",
			x"0000" when x"1768",
			x"0000" when x"1769",
			x"0000" when x"176A",
			x"0000" when x"176B",
			x"0000" when x"176C",
			x"0000" when x"176D",
			x"0000" when x"176E",
			x"0000" when x"176F",
			x"0000" when x"1770",
			x"0000" when x"1771",
			x"0000" when x"1772",
			x"0000" when x"1773",
			x"0000" when x"1774",
			x"0000" when x"1775",
			x"0000" when x"1776",
			x"0000" when x"1777",
			x"0000" when x"1778",
			x"0000" when x"1779",
			x"0000" when x"177A",
			x"0000" when x"177B",
			x"0000" when x"177C",
			x"0000" when x"177D",
			x"0000" when x"177E",
			x"0000" when x"177F",
			x"0000" when x"1780",
			x"0000" when x"1781",
			x"0000" when x"1782",
			x"0000" when x"1783",
			x"0000" when x"1784",
			x"0000" when x"1785",
			x"0000" when x"1786",
			x"0000" when x"1787",
			x"0000" when x"1788",
			x"0000" when x"1789",
			x"0000" when x"178A",
			x"0000" when x"178B",
			x"0000" when x"178C",
			x"0000" when x"178D",
			x"0000" when x"178E",
			x"0000" when x"178F",
			x"0000" when x"1790",
			x"0000" when x"1791",
			x"0000" when x"1792",
			x"0000" when x"1793",
			x"0000" when x"1794",
			x"0000" when x"1795",
			x"0000" when x"1796",
			x"0000" when x"1797",
			x"0000" when x"1798",
			x"0000" when x"1799",
			x"0000" when x"179A",
			x"0000" when x"179B",
			x"0000" when x"179C",
			x"0000" when x"179D",
			x"0000" when x"179E",
			x"0000" when x"179F",
			x"0000" when x"17A0",
			x"0000" when x"17A1",
			x"0000" when x"17A2",
			x"0000" when x"17A3",
			x"0000" when x"17A4",
			x"0000" when x"17A5",
			x"0000" when x"17A6",
			x"0000" when x"17A7",
			x"0000" when x"17A8",
			x"0000" when x"17A9",
			x"0000" when x"17AA",
			x"0000" when x"17AB",
			x"0000" when x"17AC",
			x"0000" when x"17AD",
			x"0000" when x"17AE",
			x"0000" when x"17AF",
			x"0000" when x"17B0",
			x"0000" when x"17B1",
			x"0000" when x"17B2",
			x"0000" when x"17B3",
			x"0000" when x"17B4",
			x"0000" when x"17B5",
			x"0000" when x"17B6",
			x"0000" when x"17B7",
			x"0000" when x"17B8",
			x"0000" when x"17B9",
			x"0000" when x"17BA",
			x"0000" when x"17BB",
			x"0000" when x"17BC",
			x"0000" when x"17BD",
			x"0000" when x"17BE",
			x"0000" when x"17BF",
			x"0000" when x"17C0",
			x"0000" when x"17C1",
			x"0000" when x"17C2",
			x"0000" when x"17C3",
			x"0000" when x"17C4",
			x"0000" when x"17C5",
			x"0000" when x"17C6",
			x"0000" when x"17C7",
			x"0000" when x"17C8",
			x"0000" when x"17C9",
			x"0000" when x"17CA",
			x"0000" when x"17CB",
			x"0000" when x"17CC",
			x"0000" when x"17CD",
			x"0000" when x"17CE",
			x"0000" when x"17CF",
			x"0000" when x"17D0",
			x"0000" when x"17D1",
			x"0000" when x"17D2",
			x"0000" when x"17D3",
			x"0000" when x"17D4",
			x"0000" when x"17D5",
			x"0000" when x"17D6",
			x"0000" when x"17D7",
			x"0000" when x"17D8",
			x"0000" when x"17D9",
			x"0000" when x"17DA",
			x"0000" when x"17DB",
			x"0000" when x"17DC",
			x"0000" when x"17DD",
			x"0000" when x"17DE",
			x"0000" when x"17DF",
			x"0000" when x"17E0",
			x"0000" when x"17E1",
			x"0000" when x"17E2",
			x"0000" when x"17E3",
			x"0000" when x"17E4",
			x"0000" when x"17E5",
			x"0000" when x"17E6",
			x"0000" when x"17E7",
			x"0000" when x"17E8",
			x"0000" when x"17E9",
			x"0000" when x"17EA",
			x"0000" when x"17EB",
			x"0000" when x"17EC",
			x"0000" when x"17ED",
			x"0000" when x"17EE",
			x"0000" when x"17EF",
			x"0000" when x"17F0",
			x"0000" when x"17F1",
			x"0000" when x"17F2",
			x"0000" when x"17F3",
			x"0000" when x"17F4",
			x"0000" when x"17F5",
			x"0000" when x"17F6",
			x"0000" when x"17F7",
			x"0000" when x"17F8",
			x"0000" when x"17F9",
			x"0000" when x"17FA",
			x"0000" when x"17FB",
			x"0000" when x"17FC",
			x"0000" when x"17FD",
			x"0000" when x"17FE",
			x"0000" when x"17FF",
			x"0000" when x"1800",
			x"0000" when x"1801",
			x"0000" when x"1802",
			x"0000" when x"1803",
			x"0000" when x"1804",
			x"0000" when x"1805",
			x"0000" when x"1806",
			x"0000" when x"1807",
			x"0000" when x"1808",
			x"0000" when x"1809",
			x"0000" when x"180A",
			x"0000" when x"180B",
			x"0000" when x"180C",
			x"0000" when x"180D",
			x"0000" when x"180E",
			x"0000" when x"180F",
			x"0000" when x"1810",
			x"0000" when x"1811",
			x"0000" when x"1812",
			x"0000" when x"1813",
			x"0000" when x"1814",
			x"0000" when x"1815",
			x"0000" when x"1816",
			x"0000" when x"1817",
			x"0000" when x"1818",
			x"0000" when x"1819",
			x"0000" when x"181A",
			x"0000" when x"181B",
			x"0000" when x"181C",
			x"0000" when x"181D",
			x"0000" when x"181E",
			x"0000" when x"181F",
			x"0000" when x"1820",
			x"0000" when x"1821",
			x"0000" when x"1822",
			x"0000" when x"1823",
			x"0000" when x"1824",
			x"0000" when x"1825",
			x"0000" when x"1826",
			x"0000" when x"1827",
			x"0000" when x"1828",
			x"0000" when x"1829",
			x"0000" when x"182A",
			x"0000" when x"182B",
			x"0000" when x"182C",
			x"0000" when x"182D",
			x"0000" when x"182E",
			x"0000" when x"182F",
			x"0000" when x"1830",
			x"0000" when x"1831",
			x"0000" when x"1832",
			x"0000" when x"1833",
			x"0000" when x"1834",
			x"0000" when x"1835",
			x"0000" when x"1836",
			x"0000" when x"1837",
			x"0000" when x"1838",
			x"0000" when x"1839",
			x"0000" when x"183A",
			x"0000" when x"183B",
			x"0000" when x"183C",
			x"0000" when x"183D",
			x"0000" when x"183E",
			x"0000" when x"183F",
			x"0000" when x"1840",
			x"0000" when x"1841",
			x"0000" when x"1842",
			x"0000" when x"1843",
			x"0000" when x"1844",
			x"0000" when x"1845",
			x"0000" when x"1846",
			x"0000" when x"1847",
			x"0000" when x"1848",
			x"0000" when x"1849",
			x"0000" when x"184A",
			x"0000" when x"184B",
			x"0000" when x"184C",
			x"0000" when x"184D",
			x"0000" when x"184E",
			x"0000" when x"184F",
			x"0000" when x"1850",
			x"0000" when x"1851",
			x"0000" when x"1852",
			x"0000" when x"1853",
			x"0000" when x"1854",
			x"0000" when x"1855",
			x"0000" when x"1856",
			x"0000" when x"1857",
			x"0000" when x"1858",
			x"0000" when x"1859",
			x"0000" when x"185A",
			x"0000" when x"185B",
			x"0000" when x"185C",
			x"0000" when x"185D",
			x"0000" when x"185E",
			x"0000" when x"185F",
			x"0000" when x"1860",
			x"0000" when x"1861",
			x"0000" when x"1862",
			x"0000" when x"1863",
			x"0000" when x"1864",
			x"0000" when x"1865",
			x"0000" when x"1866",
			x"0000" when x"1867",
			x"0000" when x"1868",
			x"0000" when x"1869",
			x"0000" when x"186A",
			x"0000" when x"186B",
			x"0000" when x"186C",
			x"0000" when x"186D",
			x"0000" when x"186E",
			x"0000" when x"186F",
			x"0000" when x"1870",
			x"0000" when x"1871",
			x"0000" when x"1872",
			x"0000" when x"1873",
			x"0000" when x"1874",
			x"0000" when x"1875",
			x"0000" when x"1876",
			x"0000" when x"1877",
			x"0000" when x"1878",
			x"0000" when x"1879",
			x"0000" when x"187A",
			x"0000" when x"187B",
			x"0000" when x"187C",
			x"0000" when x"187D",
			x"0000" when x"187E",
			x"0000" when x"187F",
			x"0000" when x"1880",
			x"0000" when x"1881",
			x"0000" when x"1882",
			x"0000" when x"1883",
			x"0000" when x"1884",
			x"0000" when x"1885",
			x"0000" when x"1886",
			x"0000" when x"1887",
			x"0000" when x"1888",
			x"0000" when x"1889",
			x"0000" when x"188A",
			x"0000" when x"188B",
			x"0000" when x"188C",
			x"0000" when x"188D",
			x"0000" when x"188E",
			x"0000" when x"188F",
			x"0000" when x"1890",
			x"0000" when x"1891",
			x"0000" when x"1892",
			x"0000" when x"1893",
			x"0000" when x"1894",
			x"0000" when x"1895",
			x"0000" when x"1896",
			x"0000" when x"1897",
			x"0000" when x"1898",
			x"0000" when x"1899",
			x"0000" when x"189A",
			x"0000" when x"189B",
			x"0000" when x"189C",
			x"0000" when x"189D",
			x"0000" when x"189E",
			x"0000" when x"189F",
			x"0000" when x"18A0",
			x"0000" when x"18A1",
			x"0000" when x"18A2",
			x"0000" when x"18A3",
			x"0000" when x"18A4",
			x"0000" when x"18A5",
			x"0000" when x"18A6",
			x"0000" when x"18A7",
			x"0000" when x"18A8",
			x"0000" when x"18A9",
			x"0000" when x"18AA",
			x"0000" when x"18AB",
			x"0000" when x"18AC",
			x"0000" when x"18AD",
			x"0000" when x"18AE",
			x"0000" when x"18AF",
			x"0000" when x"18B0",
			x"0000" when x"18B1",
			x"0000" when x"18B2",
			x"0000" when x"18B3",
			x"0000" when x"18B4",
			x"0000" when x"18B5",
			x"0000" when x"18B6",
			x"0000" when x"18B7",
			x"0000" when x"18B8",
			x"0000" when x"18B9",
			x"0000" when x"18BA",
			x"0000" when x"18BB",
			x"0000" when x"18BC",
			x"0000" when x"18BD",
			x"0000" when x"18BE",
			x"0000" when x"18BF",
			x"0000" when x"18C0",
			x"0000" when x"18C1",
			x"0000" when x"18C2",
			x"0000" when x"18C3",
			x"0000" when x"18C4",
			x"0000" when x"18C5",
			x"0000" when x"18C6",
			x"0000" when x"18C7",
			x"0000" when x"18C8",
			x"0000" when x"18C9",
			x"0000" when x"18CA",
			x"0000" when x"18CB",
			x"0000" when x"18CC",
			x"0000" when x"18CD",
			x"0000" when x"18CE",
			x"0000" when x"18CF",
			x"0000" when x"18D0",
			x"0000" when x"18D1",
			x"0000" when x"18D2",
			x"0000" when x"18D3",
			x"0000" when x"18D4",
			x"0000" when x"18D5",
			x"0000" when x"18D6",
			x"0000" when x"18D7",
			x"0000" when x"18D8",
			x"0000" when x"18D9",
			x"0000" when x"18DA",
			x"0000" when x"18DB",
			x"0000" when x"18DC",
			x"0000" when x"18DD",
			x"0000" when x"18DE",
			x"0000" when x"18DF",
			x"0000" when x"18E0",
			x"0000" when x"18E1",
			x"0000" when x"18E2",
			x"0000" when x"18E3",
			x"0000" when x"18E4",
			x"0000" when x"18E5",
			x"0000" when x"18E6",
			x"0000" when x"18E7",
			x"0000" when x"18E8",
			x"0000" when x"18E9",
			x"0000" when x"18EA",
			x"0000" when x"18EB",
			x"0000" when x"18EC",
			x"0000" when x"18ED",
			x"0000" when x"18EE",
			x"0000" when x"18EF",
			x"0000" when x"18F0",
			x"0000" when x"18F1",
			x"0000" when x"18F2",
			x"0000" when x"18F3",
			x"0000" when x"18F4",
			x"0000" when x"18F5",
			x"0000" when x"18F6",
			x"0000" when x"18F7",
			x"0000" when x"18F8",
			x"0000" when x"18F9",
			x"0000" when x"18FA",
			x"0000" when x"18FB",
			x"0000" when x"18FC",
			x"0000" when x"18FD",
			x"0000" when x"18FE",
			x"0000" when x"18FF",
			x"0000" when x"1900",
			x"0000" when x"1901",
			x"0000" when x"1902",
			x"0000" when x"1903",
			x"0000" when x"1904",
			x"0000" when x"1905",
			x"0000" when x"1906",
			x"0000" when x"1907",
			x"0000" when x"1908",
			x"0000" when x"1909",
			x"0000" when x"190A",
			x"0000" when x"190B",
			x"0000" when x"190C",
			x"0000" when x"190D",
			x"0000" when x"190E",
			x"0000" when x"190F",
			x"0000" when x"1910",
			x"0000" when x"1911",
			x"0000" when x"1912",
			x"0000" when x"1913",
			x"0000" when x"1914",
			x"0000" when x"1915",
			x"0000" when x"1916",
			x"0000" when x"1917",
			x"0000" when x"1918",
			x"0000" when x"1919",
			x"0000" when x"191A",
			x"0000" when x"191B",
			x"0000" when x"191C",
			x"0000" when x"191D",
			x"0000" when x"191E",
			x"0000" when x"191F",
			x"0000" when x"1920",
			x"0000" when x"1921",
			x"0000" when x"1922",
			x"0000" when x"1923",
			x"0000" when x"1924",
			x"0000" when x"1925",
			x"0000" when x"1926",
			x"0000" when x"1927",
			x"0000" when x"1928",
			x"0000" when x"1929",
			x"0000" when x"192A",
			x"0000" when x"192B",
			x"0000" when x"192C",
			x"0000" when x"192D",
			x"0000" when x"192E",
			x"0000" when x"192F",
			x"0000" when x"1930",
			x"0000" when x"1931",
			x"0000" when x"1932",
			x"0000" when x"1933",
			x"0000" when x"1934",
			x"0000" when x"1935",
			x"0000" when x"1936",
			x"0000" when x"1937",
			x"0000" when x"1938",
			x"0000" when x"1939",
			x"0000" when x"193A",
			x"0000" when x"193B",
			x"0000" when x"193C",
			x"0000" when x"193D",
			x"0000" when x"193E",
			x"0000" when x"193F",
			x"0000" when x"1940",
			x"0000" when x"1941",
			x"0000" when x"1942",
			x"0000" when x"1943",
			x"0000" when x"1944",
			x"0000" when x"1945",
			x"0000" when x"1946",
			x"0000" when x"1947",
			x"0000" when x"1948",
			x"0000" when x"1949",
			x"0000" when x"194A",
			x"0000" when x"194B",
			x"0000" when x"194C",
			x"0000" when x"194D",
			x"0000" when x"194E",
			x"0000" when x"194F",
			x"0000" when x"1950",
			x"0000" when x"1951",
			x"0000" when x"1952",
			x"0000" when x"1953",
			x"0000" when x"1954",
			x"0000" when x"1955",
			x"0000" when x"1956",
			x"0000" when x"1957",
			x"0000" when x"1958",
			x"0000" when x"1959",
			x"0000" when x"195A",
			x"0000" when x"195B",
			x"0000" when x"195C",
			x"0000" when x"195D",
			x"0000" when x"195E",
			x"0000" when x"195F",
			x"0000" when x"1960",
			x"0000" when x"1961",
			x"0000" when x"1962",
			x"0000" when x"1963",
			x"0000" when x"1964",
			x"0000" when x"1965",
			x"0000" when x"1966",
			x"0000" when x"1967",
			x"0000" when x"1968",
			x"0000" when x"1969",
			x"0000" when x"196A",
			x"0000" when x"196B",
			x"0000" when x"196C",
			x"0000" when x"196D",
			x"0000" when x"196E",
			x"0000" when x"196F",
			x"0000" when x"1970",
			x"0000" when x"1971",
			x"0000" when x"1972",
			x"0000" when x"1973",
			x"0000" when x"1974",
			x"0000" when x"1975",
			x"0000" when x"1976",
			x"0000" when x"1977",
			x"0000" when x"1978",
			x"0000" when x"1979",
			x"0000" when x"197A",
			x"0000" when x"197B",
			x"0000" when x"197C",
			x"0000" when x"197D",
			x"0000" when x"197E",
			x"0000" when x"197F",
			x"0000" when x"1980",
			x"0000" when x"1981",
			x"0000" when x"1982",
			x"0000" when x"1983",
			x"0000" when x"1984",
			x"0000" when x"1985",
			x"0000" when x"1986",
			x"0000" when x"1987",
			x"0000" when x"1988",
			x"0000" when x"1989",
			x"0000" when x"198A",
			x"0000" when x"198B",
			x"0000" when x"198C",
			x"0000" when x"198D",
			x"0000" when x"198E",
			x"0000" when x"198F",
			x"0000" when x"1990",
			x"0000" when x"1991",
			x"0000" when x"1992",
			x"0000" when x"1993",
			x"0000" when x"1994",
			x"0000" when x"1995",
			x"0000" when x"1996",
			x"0000" when x"1997",
			x"0000" when x"1998",
			x"0000" when x"1999",
			x"0000" when x"199A",
			x"0000" when x"199B",
			x"0000" when x"199C",
			x"0000" when x"199D",
			x"0000" when x"199E",
			x"0000" when x"199F",
			x"0000" when x"19A0",
			x"0000" when x"19A1",
			x"0000" when x"19A2",
			x"0000" when x"19A3",
			x"0000" when x"19A4",
			x"0000" when x"19A5",
			x"0000" when x"19A6",
			x"0000" when x"19A7",
			x"0000" when x"19A8",
			x"0000" when x"19A9",
			x"0000" when x"19AA",
			x"0000" when x"19AB",
			x"0000" when x"19AC",
			x"0000" when x"19AD",
			x"0000" when x"19AE",
			x"0000" when x"19AF",
			x"0000" when x"19B0",
			x"0000" when x"19B1",
			x"0000" when x"19B2",
			x"0000" when x"19B3",
			x"0000" when x"19B4",
			x"0000" when x"19B5",
			x"0000" when x"19B6",
			x"0000" when x"19B7",
			x"0000" when x"19B8",
			x"0000" when x"19B9",
			x"0000" when x"19BA",
			x"0000" when x"19BB",
			x"0000" when x"19BC",
			x"0000" when x"19BD",
			x"0000" when x"19BE",
			x"0000" when x"19BF",
			x"0000" when x"19C0",
			x"0000" when x"19C1",
			x"0000" when x"19C2",
			x"0000" when x"19C3",
			x"0000" when x"19C4",
			x"0000" when x"19C5",
			x"0000" when x"19C6",
			x"0000" when x"19C7",
			x"0000" when x"19C8",
			x"0000" when x"19C9",
			x"0000" when x"19CA",
			x"0000" when x"19CB",
			x"0000" when x"19CC",
			x"0000" when x"19CD",
			x"0000" when x"19CE",
			x"0000" when x"19CF",
			x"0000" when x"19D0",
			x"0000" when x"19D1",
			x"0000" when x"19D2",
			x"0000" when x"19D3",
			x"0000" when x"19D4",
			x"0000" when x"19D5",
			x"0000" when x"19D6",
			x"0000" when x"19D7",
			x"0000" when x"19D8",
			x"0000" when x"19D9",
			x"0000" when x"19DA",
			x"0000" when x"19DB",
			x"0000" when x"19DC",
			x"0000" when x"19DD",
			x"0000" when x"19DE",
			x"0000" when x"19DF",
			x"0000" when x"19E0",
			x"0000" when x"19E1",
			x"0000" when x"19E2",
			x"0000" when x"19E3",
			x"0000" when x"19E4",
			x"0000" when x"19E5",
			x"0000" when x"19E6",
			x"0000" when x"19E7",
			x"0000" when x"19E8",
			x"0000" when x"19E9",
			x"0000" when x"19EA",
			x"0000" when x"19EB",
			x"0000" when x"19EC",
			x"0000" when x"19ED",
			x"0000" when x"19EE",
			x"0000" when x"19EF",
			x"0000" when x"19F0",
			x"0000" when x"19F1",
			x"0000" when x"19F2",
			x"0000" when x"19F3",
			x"0000" when x"19F4",
			x"0000" when x"19F5",
			x"0000" when x"19F6",
			x"0000" when x"19F7",
			x"0000" when x"19F8",
			x"0000" when x"19F9",
			x"0000" when x"19FA",
			x"0000" when x"19FB",
			x"0000" when x"19FC",
			x"0000" when x"19FD",
			x"0000" when x"19FE",
			x"0000" when x"19FF",
			x"0000" when x"1A00",
			x"0000" when x"1A01",
			x"0000" when x"1A02",
			x"0000" when x"1A03",
			x"0000" when x"1A04",
			x"0000" when x"1A05",
			x"0000" when x"1A06",
			x"0000" when x"1A07",
			x"0000" when x"1A08",
			x"0000" when x"1A09",
			x"0000" when x"1A0A",
			x"0000" when x"1A0B",
			x"0000" when x"1A0C",
			x"0000" when x"1A0D",
			x"0000" when x"1A0E",
			x"0000" when x"1A0F",
			x"0000" when x"1A10",
			x"0000" when x"1A11",
			x"0000" when x"1A12",
			x"0000" when x"1A13",
			x"0000" when x"1A14",
			x"0000" when x"1A15",
			x"0000" when x"1A16",
			x"0000" when x"1A17",
			x"0000" when x"1A18",
			x"0000" when x"1A19",
			x"0000" when x"1A1A",
			x"0000" when x"1A1B",
			x"0000" when x"1A1C",
			x"0000" when x"1A1D",
			x"0000" when x"1A1E",
			x"0000" when x"1A1F",
			x"0000" when x"1A20",
			x"0000" when x"1A21",
			x"0000" when x"1A22",
			x"0000" when x"1A23",
			x"0000" when x"1A24",
			x"0000" when x"1A25",
			x"0000" when x"1A26",
			x"0000" when x"1A27",
			x"0000" when x"1A28",
			x"0000" when x"1A29",
			x"0000" when x"1A2A",
			x"0000" when x"1A2B",
			x"0000" when x"1A2C",
			x"0000" when x"1A2D",
			x"0000" when x"1A2E",
			x"0000" when x"1A2F",
			x"0000" when x"1A30",
			x"0000" when x"1A31",
			x"0000" when x"1A32",
			x"0000" when x"1A33",
			x"0000" when x"1A34",
			x"0000" when x"1A35",
			x"0000" when x"1A36",
			x"0000" when x"1A37",
			x"0000" when x"1A38",
			x"0000" when x"1A39",
			x"0000" when x"1A3A",
			x"0000" when x"1A3B",
			x"0000" when x"1A3C",
			x"0000" when x"1A3D",
			x"0000" when x"1A3E",
			x"0000" when x"1A3F",
			x"0000" when x"1A40",
			x"0000" when x"1A41",
			x"0000" when x"1A42",
			x"0000" when x"1A43",
			x"0000" when x"1A44",
			x"0000" when x"1A45",
			x"0000" when x"1A46",
			x"0000" when x"1A47",
			x"0000" when x"1A48",
			x"0000" when x"1A49",
			x"0000" when x"1A4A",
			x"0000" when x"1A4B",
			x"0000" when x"1A4C",
			x"0000" when x"1A4D",
			x"0000" when x"1A4E",
			x"0000" when x"1A4F",
			x"0000" when x"1A50",
			x"0000" when x"1A51",
			x"0000" when x"1A52",
			x"0000" when x"1A53",
			x"0000" when x"1A54",
			x"0000" when x"1A55",
			x"0000" when x"1A56",
			x"0000" when x"1A57",
			x"0000" when x"1A58",
			x"0000" when x"1A59",
			x"0000" when x"1A5A",
			x"0000" when x"1A5B",
			x"0000" when x"1A5C",
			x"0000" when x"1A5D",
			x"0000" when x"1A5E",
			x"0000" when x"1A5F",
			x"0000" when x"1A60",
			x"0000" when x"1A61",
			x"0000" when x"1A62",
			x"0000" when x"1A63",
			x"0000" when x"1A64",
			x"0000" when x"1A65",
			x"0000" when x"1A66",
			x"0000" when x"1A67",
			x"0000" when x"1A68",
			x"0000" when x"1A69",
			x"0000" when x"1A6A",
			x"0000" when x"1A6B",
			x"0000" when x"1A6C",
			x"0000" when x"1A6D",
			x"0000" when x"1A6E",
			x"0000" when x"1A6F",
			x"0000" when x"1A70",
			x"0000" when x"1A71",
			x"0000" when x"1A72",
			x"0000" when x"1A73",
			x"0000" when x"1A74",
			x"0000" when x"1A75",
			x"0000" when x"1A76",
			x"0000" when x"1A77",
			x"0000" when x"1A78",
			x"0000" when x"1A79",
			x"0000" when x"1A7A",
			x"0000" when x"1A7B",
			x"0000" when x"1A7C",
			x"0000" when x"1A7D",
			x"0000" when x"1A7E",
			x"0000" when x"1A7F",
			x"0000" when x"1A80",
			x"0000" when x"1A81",
			x"0000" when x"1A82",
			x"0000" when x"1A83",
			x"0000" when x"1A84",
			x"0000" when x"1A85",
			x"0000" when x"1A86",
			x"0000" when x"1A87",
			x"0000" when x"1A88",
			x"0000" when x"1A89",
			x"0000" when x"1A8A",
			x"0000" when x"1A8B",
			x"0000" when x"1A8C",
			x"0000" when x"1A8D",
			x"0000" when x"1A8E",
			x"0000" when x"1A8F",
			x"0000" when x"1A90",
			x"0000" when x"1A91",
			x"0000" when x"1A92",
			x"0000" when x"1A93",
			x"0000" when x"1A94",
			x"0000" when x"1A95",
			x"0000" when x"1A96",
			x"0000" when x"1A97",
			x"0000" when x"1A98",
			x"0000" when x"1A99",
			x"0000" when x"1A9A",
			x"0000" when x"1A9B",
			x"0000" when x"1A9C",
			x"0000" when x"1A9D",
			x"0000" when x"1A9E",
			x"0000" when x"1A9F",
			x"0000" when x"1AA0",
			x"0000" when x"1AA1",
			x"0000" when x"1AA2",
			x"0000" when x"1AA3",
			x"0000" when x"1AA4",
			x"0000" when x"1AA5",
			x"0000" when x"1AA6",
			x"0000" when x"1AA7",
			x"0000" when x"1AA8",
			x"0000" when x"1AA9",
			x"0000" when x"1AAA",
			x"0000" when x"1AAB",
			x"0000" when x"1AAC",
			x"0000" when x"1AAD",
			x"0000" when x"1AAE",
			x"0000" when x"1AAF",
			x"0000" when x"1AB0",
			x"0000" when x"1AB1",
			x"0000" when x"1AB2",
			x"0000" when x"1AB3",
			x"0000" when x"1AB4",
			x"0000" when x"1AB5",
			x"0000" when x"1AB6",
			x"0000" when x"1AB7",
			x"0000" when x"1AB8",
			x"0000" when x"1AB9",
			x"0000" when x"1ABA",
			x"0000" when x"1ABB",
			x"0000" when x"1ABC",
			x"0000" when x"1ABD",
			x"0000" when x"1ABE",
			x"0000" when x"1ABF",
			x"0000" when x"1AC0",
			x"0000" when x"1AC1",
			x"0000" when x"1AC2",
			x"0000" when x"1AC3",
			x"0000" when x"1AC4",
			x"0000" when x"1AC5",
			x"0000" when x"1AC6",
			x"0000" when x"1AC7",
			x"0000" when x"1AC8",
			x"0000" when x"1AC9",
			x"0000" when x"1ACA",
			x"0000" when x"1ACB",
			x"0000" when x"1ACC",
			x"0000" when x"1ACD",
			x"0000" when x"1ACE",
			x"0000" when x"1ACF",
			x"0000" when x"1AD0",
			x"0000" when x"1AD1",
			x"0000" when x"1AD2",
			x"0000" when x"1AD3",
			x"0000" when x"1AD4",
			x"0000" when x"1AD5",
			x"0000" when x"1AD6",
			x"0000" when x"1AD7",
			x"0000" when x"1AD8",
			x"0000" when x"1AD9",
			x"0000" when x"1ADA",
			x"0000" when x"1ADB",
			x"0000" when x"1ADC",
			x"0000" when x"1ADD",
			x"0000" when x"1ADE",
			x"0000" when x"1ADF",
			x"0000" when x"1AE0",
			x"0000" when x"1AE1",
			x"0000" when x"1AE2",
			x"0000" when x"1AE3",
			x"0000" when x"1AE4",
			x"0000" when x"1AE5",
			x"0000" when x"1AE6",
			x"0000" when x"1AE7",
			x"0000" when x"1AE8",
			x"0000" when x"1AE9",
			x"0000" when x"1AEA",
			x"0000" when x"1AEB",
			x"0000" when x"1AEC",
			x"0000" when x"1AED",
			x"0000" when x"1AEE",
			x"0000" when x"1AEF",
			x"0000" when x"1AF0",
			x"0000" when x"1AF1",
			x"0000" when x"1AF2",
			x"0000" when x"1AF3",
			x"0000" when x"1AF4",
			x"0000" when x"1AF5",
			x"0000" when x"1AF6",
			x"0000" when x"1AF7",
			x"0000" when x"1AF8",
			x"0000" when x"1AF9",
			x"0000" when x"1AFA",
			x"0000" when x"1AFB",
			x"0000" when x"1AFC",
			x"0000" when x"1AFD",
			x"0000" when x"1AFE",
			x"0000" when x"1AFF",
			x"0000" when x"1B00",
			x"0000" when x"1B01",
			x"0000" when x"1B02",
			x"0000" when x"1B03",
			x"0000" when x"1B04",
			x"0000" when x"1B05",
			x"0000" when x"1B06",
			x"0000" when x"1B07",
			x"0000" when x"1B08",
			x"0000" when x"1B09",
			x"0000" when x"1B0A",
			x"0000" when x"1B0B",
			x"0000" when x"1B0C",
			x"0000" when x"1B0D",
			x"0000" when x"1B0E",
			x"0000" when x"1B0F",
			x"0000" when x"1B10",
			x"0000" when x"1B11",
			x"0000" when x"1B12",
			x"0000" when x"1B13",
			x"0000" when x"1B14",
			x"0000" when x"1B15",
			x"0000" when x"1B16",
			x"0000" when x"1B17",
			x"0000" when x"1B18",
			x"0000" when x"1B19",
			x"0000" when x"1B1A",
			x"0000" when x"1B1B",
			x"0000" when x"1B1C",
			x"0000" when x"1B1D",
			x"0000" when x"1B1E",
			x"0000" when x"1B1F",
			x"0000" when x"1B20",
			x"0000" when x"1B21",
			x"0000" when x"1B22",
			x"0000" when x"1B23",
			x"0000" when x"1B24",
			x"0000" when x"1B25",
			x"0000" when x"1B26",
			x"0000" when x"1B27",
			x"0000" when x"1B28",
			x"0000" when x"1B29",
			x"0000" when x"1B2A",
			x"0000" when x"1B2B",
			x"0000" when x"1B2C",
			x"0000" when x"1B2D",
			x"0000" when x"1B2E",
			x"0000" when x"1B2F",
			x"0000" when x"1B30",
			x"0000" when x"1B31",
			x"0000" when x"1B32",
			x"0000" when x"1B33",
			x"0000" when x"1B34",
			x"0000" when x"1B35",
			x"0000" when x"1B36",
			x"0000" when x"1B37",
			x"0000" when x"1B38",
			x"0000" when x"1B39",
			x"0000" when x"1B3A",
			x"0000" when x"1B3B",
			x"0000" when x"1B3C",
			x"0000" when x"1B3D",
			x"0000" when x"1B3E",
			x"0000" when x"1B3F",
			x"0000" when x"1B40",
			x"0000" when x"1B41",
			x"0000" when x"1B42",
			x"0000" when x"1B43",
			x"0000" when x"1B44",
			x"0000" when x"1B45",
			x"0000" when x"1B46",
			x"0000" when x"1B47",
			x"0000" when x"1B48",
			x"0000" when x"1B49",
			x"0000" when x"1B4A",
			x"0000" when x"1B4B",
			x"0000" when x"1B4C",
			x"0000" when x"1B4D",
			x"0000" when x"1B4E",
			x"0000" when x"1B4F",
			x"0000" when x"1B50",
			x"0000" when x"1B51",
			x"0000" when x"1B52",
			x"0000" when x"1B53",
			x"0000" when x"1B54",
			x"0000" when x"1B55",
			x"0000" when x"1B56",
			x"0000" when x"1B57",
			x"0000" when x"1B58",
			x"0000" when x"1B59",
			x"0000" when x"1B5A",
			x"0000" when x"1B5B",
			x"0000" when x"1B5C",
			x"0000" when x"1B5D",
			x"0000" when x"1B5E",
			x"0000" when x"1B5F",
			x"0000" when x"1B60",
			x"0000" when x"1B61",
			x"0000" when x"1B62",
			x"0000" when x"1B63",
			x"0000" when x"1B64",
			x"0000" when x"1B65",
			x"0000" when x"1B66",
			x"0000" when x"1B67",
			x"0000" when x"1B68",
			x"0000" when x"1B69",
			x"0000" when x"1B6A",
			x"0000" when x"1B6B",
			x"0000" when x"1B6C",
			x"0000" when x"1B6D",
			x"0000" when x"1B6E",
			x"0000" when x"1B6F",
			x"0000" when x"1B70",
			x"0000" when x"1B71",
			x"0000" when x"1B72",
			x"0000" when x"1B73",
			x"0000" when x"1B74",
			x"0000" when x"1B75",
			x"0000" when x"1B76",
			x"0000" when x"1B77",
			x"0000" when x"1B78",
			x"0000" when x"1B79",
			x"0000" when x"1B7A",
			x"0000" when x"1B7B",
			x"0000" when x"1B7C",
			x"0000" when x"1B7D",
			x"0000" when x"1B7E",
			x"0000" when x"1B7F",
			x"0000" when x"1B80",
			x"0000" when x"1B81",
			x"0000" when x"1B82",
			x"0000" when x"1B83",
			x"0000" when x"1B84",
			x"0000" when x"1B85",
			x"0000" when x"1B86",
			x"0000" when x"1B87",
			x"0000" when x"1B88",
			x"0000" when x"1B89",
			x"0000" when x"1B8A",
			x"0000" when x"1B8B",
			x"0000" when x"1B8C",
			x"0000" when x"1B8D",
			x"0000" when x"1B8E",
			x"0000" when x"1B8F",
			x"0000" when x"1B90",
			x"0000" when x"1B91",
			x"0000" when x"1B92",
			x"0000" when x"1B93",
			x"0000" when x"1B94",
			x"0000" when x"1B95",
			x"0000" when x"1B96",
			x"0000" when x"1B97",
			x"0000" when x"1B98",
			x"0000" when x"1B99",
			x"0000" when x"1B9A",
			x"0000" when x"1B9B",
			x"0000" when x"1B9C",
			x"0000" when x"1B9D",
			x"0000" when x"1B9E",
			x"0000" when x"1B9F",
			x"0000" when x"1BA0",
			x"0000" when x"1BA1",
			x"0000" when x"1BA2",
			x"0000" when x"1BA3",
			x"0000" when x"1BA4",
			x"0000" when x"1BA5",
			x"0000" when x"1BA6",
			x"0000" when x"1BA7",
			x"0000" when x"1BA8",
			x"0000" when x"1BA9",
			x"0000" when x"1BAA",
			x"0000" when x"1BAB",
			x"0000" when x"1BAC",
			x"0000" when x"1BAD",
			x"0000" when x"1BAE",
			x"0000" when x"1BAF",
			x"0000" when x"1BB0",
			x"0000" when x"1BB1",
			x"0000" when x"1BB2",
			x"0000" when x"1BB3",
			x"0000" when x"1BB4",
			x"0000" when x"1BB5",
			x"0000" when x"1BB6",
			x"0000" when x"1BB7",
			x"0000" when x"1BB8",
			x"0000" when x"1BB9",
			x"0000" when x"1BBA",
			x"0000" when x"1BBB",
			x"0000" when x"1BBC",
			x"0000" when x"1BBD",
			x"0000" when x"1BBE",
			x"0000" when x"1BBF",
			x"0000" when x"1BC0",
			x"0000" when x"1BC1",
			x"0000" when x"1BC2",
			x"0000" when x"1BC3",
			x"0000" when x"1BC4",
			x"0000" when x"1BC5",
			x"0000" when x"1BC6",
			x"0000" when x"1BC7",
			x"0000" when x"1BC8",
			x"0000" when x"1BC9",
			x"0000" when x"1BCA",
			x"0000" when x"1BCB",
			x"0000" when x"1BCC",
			x"0000" when x"1BCD",
			x"0000" when x"1BCE",
			x"0000" when x"1BCF",
			x"0000" when x"1BD0",
			x"0000" when x"1BD1",
			x"0000" when x"1BD2",
			x"0000" when x"1BD3",
			x"0000" when x"1BD4",
			x"0000" when x"1BD5",
			x"0000" when x"1BD6",
			x"0000" when x"1BD7",
			x"0000" when x"1BD8",
			x"0000" when x"1BD9",
			x"0000" when x"1BDA",
			x"0000" when x"1BDB",
			x"0000" when x"1BDC",
			x"0000" when x"1BDD",
			x"0000" when x"1BDE",
			x"0000" when x"1BDF",
			x"0000" when x"1BE0",
			x"0000" when x"1BE1",
			x"0000" when x"1BE2",
			x"0000" when x"1BE3",
			x"0000" when x"1BE4",
			x"0000" when x"1BE5",
			x"0000" when x"1BE6",
			x"0000" when x"1BE7",
			x"0000" when x"1BE8",
			x"0000" when x"1BE9",
			x"0000" when x"1BEA",
			x"0000" when x"1BEB",
			x"0000" when x"1BEC",
			x"0000" when x"1BED",
			x"0000" when x"1BEE",
			x"0000" when x"1BEF",
			x"0000" when x"1BF0",
			x"0000" when x"1BF1",
			x"0000" when x"1BF2",
			x"0000" when x"1BF3",
			x"0000" when x"1BF4",
			x"0000" when x"1BF5",
			x"0000" when x"1BF6",
			x"0000" when x"1BF7",
			x"0000" when x"1BF8",
			x"0000" when x"1BF9",
			x"0000" when x"1BFA",
			x"0000" when x"1BFB",
			x"0000" when x"1BFC",
			x"0000" when x"1BFD",
			x"0000" when x"1BFE",
			x"0000" when x"1BFF",
			x"0000" when x"1C00",
			x"0000" when x"1C01",
			x"0000" when x"1C02",
			x"0000" when x"1C03",
			x"0000" when x"1C04",
			x"0000" when x"1C05",
			x"0000" when x"1C06",
			x"0000" when x"1C07",
			x"0000" when x"1C08",
			x"0000" when x"1C09",
			x"0000" when x"1C0A",
			x"0000" when x"1C0B",
			x"0000" when x"1C0C",
			x"0000" when x"1C0D",
			x"0000" when x"1C0E",
			x"0000" when x"1C0F",
			x"0000" when x"1C10",
			x"0000" when x"1C11",
			x"0000" when x"1C12",
			x"0000" when x"1C13",
			x"0000" when x"1C14",
			x"0000" when x"1C15",
			x"0000" when x"1C16",
			x"0000" when x"1C17",
			x"0000" when x"1C18",
			x"0000" when x"1C19",
			x"0000" when x"1C1A",
			x"0000" when x"1C1B",
			x"0000" when x"1C1C",
			x"0000" when x"1C1D",
			x"0000" when x"1C1E",
			x"0000" when x"1C1F",
			x"0000" when x"1C20",
			x"0000" when x"1C21",
			x"0000" when x"1C22",
			x"0000" when x"1C23",
			x"0000" when x"1C24",
			x"0000" when x"1C25",
			x"0000" when x"1C26",
			x"0000" when x"1C27",
			x"0000" when x"1C28",
			x"0000" when x"1C29",
			x"0000" when x"1C2A",
			x"0000" when x"1C2B",
			x"0000" when x"1C2C",
			x"0000" when x"1C2D",
			x"0000" when x"1C2E",
			x"0000" when x"1C2F",
			x"0000" when x"1C30",
			x"0000" when x"1C31",
			x"0000" when x"1C32",
			x"0000" when x"1C33",
			x"0000" when x"1C34",
			x"0000" when x"1C35",
			x"0000" when x"1C36",
			x"0000" when x"1C37",
			x"0000" when x"1C38",
			x"0000" when x"1C39",
			x"0000" when x"1C3A",
			x"0000" when x"1C3B",
			x"0000" when x"1C3C",
			x"0000" when x"1C3D",
			x"0000" when x"1C3E",
			x"0000" when x"1C3F",
			x"0000" when x"1C40",
			x"0000" when x"1C41",
			x"0000" when x"1C42",
			x"0000" when x"1C43",
			x"0000" when x"1C44",
			x"0000" when x"1C45",
			x"0000" when x"1C46",
			x"0000" when x"1C47",
			x"0000" when x"1C48",
			x"0000" when x"1C49",
			x"0000" when x"1C4A",
			x"0000" when x"1C4B",
			x"0000" when x"1C4C",
			x"0000" when x"1C4D",
			x"0000" when x"1C4E",
			x"0000" when x"1C4F",
			x"0000" when x"1C50",
			x"0000" when x"1C51",
			x"0000" when x"1C52",
			x"0000" when x"1C53",
			x"0000" when x"1C54",
			x"0000" when x"1C55",
			x"0000" when x"1C56",
			x"0000" when x"1C57",
			x"0000" when x"1C58",
			x"0000" when x"1C59",
			x"0000" when x"1C5A",
			x"0000" when x"1C5B",
			x"0000" when x"1C5C",
			x"0000" when x"1C5D",
			x"0000" when x"1C5E",
			x"0000" when x"1C5F",
			x"0000" when x"1C60",
			x"0000" when x"1C61",
			x"0000" when x"1C62",
			x"0000" when x"1C63",
			x"0000" when x"1C64",
			x"0000" when x"1C65",
			x"0000" when x"1C66",
			x"0000" when x"1C67",
			x"0000" when x"1C68",
			x"0000" when x"1C69",
			x"0000" when x"1C6A",
			x"0000" when x"1C6B",
			x"0000" when x"1C6C",
			x"0000" when x"1C6D",
			x"0000" when x"1C6E",
			x"0000" when x"1C6F",
			x"0000" when x"1C70",
			x"0000" when x"1C71",
			x"0000" when x"1C72",
			x"0000" when x"1C73",
			x"0000" when x"1C74",
			x"0000" when x"1C75",
			x"0000" when x"1C76",
			x"0000" when x"1C77",
			x"0000" when x"1C78",
			x"0000" when x"1C79",
			x"0000" when x"1C7A",
			x"0000" when x"1C7B",
			x"0000" when x"1C7C",
			x"0000" when x"1C7D",
			x"0000" when x"1C7E",
			x"0000" when x"1C7F",
			x"0000" when x"1C80",
			x"0000" when x"1C81",
			x"0000" when x"1C82",
			x"0000" when x"1C83",
			x"0000" when x"1C84",
			x"0000" when x"1C85",
			x"0000" when x"1C86",
			x"0000" when x"1C87",
			x"0000" when x"1C88",
			x"0000" when x"1C89",
			x"0000" when x"1C8A",
			x"0000" when x"1C8B",
			x"0000" when x"1C8C",
			x"0000" when x"1C8D",
			x"0000" when x"1C8E",
			x"0000" when x"1C8F",
			x"0000" when x"1C90",
			x"0000" when x"1C91",
			x"0000" when x"1C92",
			x"0000" when x"1C93",
			x"0000" when x"1C94",
			x"0000" when x"1C95",
			x"0000" when x"1C96",
			x"0000" when x"1C97",
			x"0000" when x"1C98",
			x"0000" when x"1C99",
			x"0000" when x"1C9A",
			x"0000" when x"1C9B",
			x"0000" when x"1C9C",
			x"0000" when x"1C9D",
			x"0000" when x"1C9E",
			x"0000" when x"1C9F",
			x"0000" when x"1CA0",
			x"0000" when x"1CA1",
			x"0000" when x"1CA2",
			x"0000" when x"1CA3",
			x"0000" when x"1CA4",
			x"0000" when x"1CA5",
			x"0000" when x"1CA6",
			x"0000" when x"1CA7",
			x"0000" when x"1CA8",
			x"0000" when x"1CA9",
			x"0000" when x"1CAA",
			x"0000" when x"1CAB",
			x"0000" when x"1CAC",
			x"0000" when x"1CAD",
			x"0000" when x"1CAE",
			x"0000" when x"1CAF",
			x"0000" when x"1CB0",
			x"0000" when x"1CB1",
			x"0000" when x"1CB2",
			x"0000" when x"1CB3",
			x"0000" when x"1CB4",
			x"0000" when x"1CB5",
			x"0000" when x"1CB6",
			x"0000" when x"1CB7",
			x"0000" when x"1CB8",
			x"0000" when x"1CB9",
			x"0000" when x"1CBA",
			x"0000" when x"1CBB",
			x"0000" when x"1CBC",
			x"0000" when x"1CBD",
			x"0000" when x"1CBE",
			x"0000" when x"1CBF",
			x"0000" when x"1CC0",
			x"0000" when x"1CC1",
			x"0000" when x"1CC2",
			x"0000" when x"1CC3",
			x"0000" when x"1CC4",
			x"0000" when x"1CC5",
			x"0000" when x"1CC6",
			x"0000" when x"1CC7",
			x"0000" when x"1CC8",
			x"0000" when x"1CC9",
			x"0000" when x"1CCA",
			x"0000" when x"1CCB",
			x"0000" when x"1CCC",
			x"0000" when x"1CCD",
			x"0000" when x"1CCE",
			x"0000" when x"1CCF",
			x"0000" when x"1CD0",
			x"0000" when x"1CD1",
			x"0000" when x"1CD2",
			x"0000" when x"1CD3",
			x"0000" when x"1CD4",
			x"0000" when x"1CD5",
			x"0000" when x"1CD6",
			x"0000" when x"1CD7",
			x"0000" when x"1CD8",
			x"0000" when x"1CD9",
			x"0000" when x"1CDA",
			x"0000" when x"1CDB",
			x"0000" when x"1CDC",
			x"0000" when x"1CDD",
			x"0000" when x"1CDE",
			x"0000" when x"1CDF",
			x"0000" when x"1CE0",
			x"0000" when x"1CE1",
			x"0000" when x"1CE2",
			x"0000" when x"1CE3",
			x"0000" when x"1CE4",
			x"0000" when x"1CE5",
			x"0000" when x"1CE6",
			x"0000" when x"1CE7",
			x"0000" when x"1CE8",
			x"0000" when x"1CE9",
			x"0000" when x"1CEA",
			x"0000" when x"1CEB",
			x"0000" when x"1CEC",
			x"0000" when x"1CED",
			x"0000" when x"1CEE",
			x"0000" when x"1CEF",
			x"0000" when x"1CF0",
			x"0000" when x"1CF1",
			x"0000" when x"1CF2",
			x"0000" when x"1CF3",
			x"0000" when x"1CF4",
			x"0000" when x"1CF5",
			x"0000" when x"1CF6",
			x"0000" when x"1CF7",
			x"0000" when x"1CF8",
			x"0000" when x"1CF9",
			x"0000" when x"1CFA",
			x"0000" when x"1CFB",
			x"0000" when x"1CFC",
			x"0000" when x"1CFD",
			x"0000" when x"1CFE",
			x"0000" when x"1CFF",
			x"0000" when x"1D00",
			x"0000" when x"1D01",
			x"0000" when x"1D02",
			x"0000" when x"1D03",
			x"0000" when x"1D04",
			x"0000" when x"1D05",
			x"0000" when x"1D06",
			x"0000" when x"1D07",
			x"0000" when x"1D08",
			x"0000" when x"1D09",
			x"0000" when x"1D0A",
			x"0000" when x"1D0B",
			x"0000" when x"1D0C",
			x"0000" when x"1D0D",
			x"0000" when x"1D0E",
			x"0000" when x"1D0F",
			x"0000" when x"1D10",
			x"0000" when x"1D11",
			x"0000" when x"1D12",
			x"0000" when x"1D13",
			x"0000" when x"1D14",
			x"0000" when x"1D15",
			x"0000" when x"1D16",
			x"0000" when x"1D17",
			x"0000" when x"1D18",
			x"0000" when x"1D19",
			x"0000" when x"1D1A",
			x"0000" when x"1D1B",
			x"0000" when x"1D1C",
			x"0000" when x"1D1D",
			x"0000" when x"1D1E",
			x"0000" when x"1D1F",
			x"0000" when x"1D20",
			x"0000" when x"1D21",
			x"0000" when x"1D22",
			x"0000" when x"1D23",
			x"0000" when x"1D24",
			x"0000" when x"1D25",
			x"0000" when x"1D26",
			x"0000" when x"1D27",
			x"0000" when x"1D28",
			x"0000" when x"1D29",
			x"0000" when x"1D2A",
			x"0000" when x"1D2B",
			x"0000" when x"1D2C",
			x"0000" when x"1D2D",
			x"0000" when x"1D2E",
			x"0000" when x"1D2F",
			x"0000" when x"1D30",
			x"0000" when x"1D31",
			x"0000" when x"1D32",
			x"0000" when x"1D33",
			x"0000" when x"1D34",
			x"0000" when x"1D35",
			x"0000" when x"1D36",
			x"0000" when x"1D37",
			x"0000" when x"1D38",
			x"0000" when x"1D39",
			x"0000" when x"1D3A",
			x"0000" when x"1D3B",
			x"0000" when x"1D3C",
			x"0000" when x"1D3D",
			x"0000" when x"1D3E",
			x"0000" when x"1D3F",
			x"0000" when x"1D40",
			x"0000" when x"1D41",
			x"0000" when x"1D42",
			x"0000" when x"1D43",
			x"0000" when x"1D44",
			x"0000" when x"1D45",
			x"0000" when x"1D46",
			x"0000" when x"1D47",
			x"0000" when x"1D48",
			x"0000" when x"1D49",
			x"0000" when x"1D4A",
			x"0000" when x"1D4B",
			x"0000" when x"1D4C",
			x"0000" when x"1D4D",
			x"0000" when x"1D4E",
			x"0000" when x"1D4F",
			x"0000" when x"1D50",
			x"0000" when x"1D51",
			x"0000" when x"1D52",
			x"0000" when x"1D53",
			x"0000" when x"1D54",
			x"0000" when x"1D55",
			x"0000" when x"1D56",
			x"0000" when x"1D57",
			x"0000" when x"1D58",
			x"0000" when x"1D59",
			x"0000" when x"1D5A",
			x"0000" when x"1D5B",
			x"0000" when x"1D5C",
			x"0000" when x"1D5D",
			x"0000" when x"1D5E",
			x"0000" when x"1D5F",
			x"0000" when x"1D60",
			x"0000" when x"1D61",
			x"0000" when x"1D62",
			x"0000" when x"1D63",
			x"0000" when x"1D64",
			x"0000" when x"1D65",
			x"0000" when x"1D66",
			x"0000" when x"1D67",
			x"0000" when x"1D68",
			x"0000" when x"1D69",
			x"0000" when x"1D6A",
			x"0000" when x"1D6B",
			x"0000" when x"1D6C",
			x"0000" when x"1D6D",
			x"0000" when x"1D6E",
			x"0000" when x"1D6F",
			x"0000" when x"1D70",
			x"0000" when x"1D71",
			x"0000" when x"1D72",
			x"0000" when x"1D73",
			x"0000" when x"1D74",
			x"0000" when x"1D75",
			x"0000" when x"1D76",
			x"0000" when x"1D77",
			x"0000" when x"1D78",
			x"0000" when x"1D79",
			x"0000" when x"1D7A",
			x"0000" when x"1D7B",
			x"0000" when x"1D7C",
			x"0000" when x"1D7D",
			x"0000" when x"1D7E",
			x"0000" when x"1D7F",
			x"0000" when x"1D80",
			x"0000" when x"1D81",
			x"0000" when x"1D82",
			x"0000" when x"1D83",
			x"0000" when x"1D84",
			x"0000" when x"1D85",
			x"0000" when x"1D86",
			x"0000" when x"1D87",
			x"0000" when x"1D88",
			x"0000" when x"1D89",
			x"0000" when x"1D8A",
			x"0000" when x"1D8B",
			x"0000" when x"1D8C",
			x"0000" when x"1D8D",
			x"0000" when x"1D8E",
			x"0000" when x"1D8F",
			x"0000" when x"1D90",
			x"0000" when x"1D91",
			x"0000" when x"1D92",
			x"0000" when x"1D93",
			x"0000" when x"1D94",
			x"0000" when x"1D95",
			x"0000" when x"1D96",
			x"0000" when x"1D97",
			x"0000" when x"1D98",
			x"0000" when x"1D99",
			x"0000" when x"1D9A",
			x"0000" when x"1D9B",
			x"0000" when x"1D9C",
			x"0000" when x"1D9D",
			x"0000" when x"1D9E",
			x"0000" when x"1D9F",
			x"0000" when x"1DA0",
			x"0000" when x"1DA1",
			x"0000" when x"1DA2",
			x"0000" when x"1DA3",
			x"0000" when x"1DA4",
			x"0000" when x"1DA5",
			x"0000" when x"1DA6",
			x"0000" when x"1DA7",
			x"0000" when x"1DA8",
			x"0000" when x"1DA9",
			x"0000" when x"1DAA",
			x"0000" when x"1DAB",
			x"0000" when x"1DAC",
			x"0000" when x"1DAD",
			x"0000" when x"1DAE",
			x"0000" when x"1DAF",
			x"0000" when x"1DB0",
			x"0000" when x"1DB1",
			x"0000" when x"1DB2",
			x"0000" when x"1DB3",
			x"0000" when x"1DB4",
			x"0000" when x"1DB5",
			x"0000" when x"1DB6",
			x"0000" when x"1DB7",
			x"0000" when x"1DB8",
			x"0000" when x"1DB9",
			x"0000" when x"1DBA",
			x"0000" when x"1DBB",
			x"0000" when x"1DBC",
			x"0000" when x"1DBD",
			x"0000" when x"1DBE",
			x"0000" when x"1DBF",
			x"0000" when x"1DC0",
			x"0000" when x"1DC1",
			x"0000" when x"1DC2",
			x"0000" when x"1DC3",
			x"0000" when x"1DC4",
			x"0000" when x"1DC5",
			x"0000" when x"1DC6",
			x"0000" when x"1DC7",
			x"0000" when x"1DC8",
			x"0000" when x"1DC9",
			x"0000" when x"1DCA",
			x"0000" when x"1DCB",
			x"0000" when x"1DCC",
			x"0000" when x"1DCD",
			x"0000" when x"1DCE",
			x"0000" when x"1DCF",
			x"0000" when x"1DD0",
			x"0000" when x"1DD1",
			x"0000" when x"1DD2",
			x"0000" when x"1DD3",
			x"0000" when x"1DD4",
			x"0000" when x"1DD5",
			x"0000" when x"1DD6",
			x"0000" when x"1DD7",
			x"0000" when x"1DD8",
			x"0000" when x"1DD9",
			x"0000" when x"1DDA",
			x"0000" when x"1DDB",
			x"0000" when x"1DDC",
			x"0000" when x"1DDD",
			x"0000" when x"1DDE",
			x"0000" when x"1DDF",
			x"0000" when x"1DE0",
			x"0000" when x"1DE1",
			x"0000" when x"1DE2",
			x"0000" when x"1DE3",
			x"0000" when x"1DE4",
			x"0000" when x"1DE5",
			x"0000" when x"1DE6",
			x"0000" when x"1DE7",
			x"0000" when x"1DE8",
			x"0000" when x"1DE9",
			x"0000" when x"1DEA",
			x"0000" when x"1DEB",
			x"0000" when x"1DEC",
			x"0000" when x"1DED",
			x"0000" when x"1DEE",
			x"0000" when x"1DEF",
			x"0000" when x"1DF0",
			x"0000" when x"1DF1",
			x"0000" when x"1DF2",
			x"0000" when x"1DF3",
			x"0000" when x"1DF4",
			x"0000" when x"1DF5",
			x"0000" when x"1DF6",
			x"0000" when x"1DF7",
			x"0000" when x"1DF8",
			x"0000" when x"1DF9",
			x"0000" when x"1DFA",
			x"0000" when x"1DFB",
			x"0000" when x"1DFC",
			x"0000" when x"1DFD",
			x"0000" when x"1DFE",
			x"0000" when x"1DFF",
			x"0000" when x"1E00",
			x"0000" when x"1E01",
			x"0000" when x"1E02",
			x"0000" when x"1E03",
			x"0000" when x"1E04",
			x"0000" when x"1E05",
			x"0000" when x"1E06",
			x"0000" when x"1E07",
			x"0000" when x"1E08",
			x"0000" when x"1E09",
			x"0000" when x"1E0A",
			x"0000" when x"1E0B",
			x"0000" when x"1E0C",
			x"0000" when x"1E0D",
			x"0000" when x"1E0E",
			x"0000" when x"1E0F",
			x"0000" when x"1E10",
			x"0000" when x"1E11",
			x"0000" when x"1E12",
			x"0000" when x"1E13",
			x"0000" when x"1E14",
			x"0000" when x"1E15",
			x"0000" when x"1E16",
			x"0000" when x"1E17",
			x"0000" when x"1E18",
			x"0000" when x"1E19",
			x"0000" when x"1E1A",
			x"0000" when x"1E1B",
			x"0000" when x"1E1C",
			x"0000" when x"1E1D",
			x"0000" when x"1E1E",
			x"0000" when x"1E1F",
			x"0000" when x"1E20",
			x"0000" when x"1E21",
			x"0000" when x"1E22",
			x"0000" when x"1E23",
			x"0000" when x"1E24",
			x"0000" when x"1E25",
			x"0000" when x"1E26",
			x"0000" when x"1E27",
			x"0000" when x"1E28",
			x"0000" when x"1E29",
			x"0000" when x"1E2A",
			x"0000" when x"1E2B",
			x"0000" when x"1E2C",
			x"0000" when x"1E2D",
			x"0000" when x"1E2E",
			x"0000" when x"1E2F",
			x"0000" when x"1E30",
			x"0000" when x"1E31",
			x"0000" when x"1E32",
			x"0000" when x"1E33",
			x"0000" when x"1E34",
			x"0000" when x"1E35",
			x"0000" when x"1E36",
			x"0000" when x"1E37",
			x"0000" when x"1E38",
			x"0000" when x"1E39",
			x"0000" when x"1E3A",
			x"0000" when x"1E3B",
			x"0000" when x"1E3C",
			x"0000" when x"1E3D",
			x"0000" when x"1E3E",
			x"0000" when x"1E3F",
			x"0000" when x"1E40",
			x"0000" when x"1E41",
			x"0000" when x"1E42",
			x"0000" when x"1E43",
			x"0000" when x"1E44",
			x"0000" when x"1E45",
			x"0000" when x"1E46",
			x"0000" when x"1E47",
			x"0000" when x"1E48",
			x"0000" when x"1E49",
			x"0000" when x"1E4A",
			x"0000" when x"1E4B",
			x"0000" when x"1E4C",
			x"0000" when x"1E4D",
			x"0000" when x"1E4E",
			x"0000" when x"1E4F",
			x"0000" when x"1E50",
			x"0000" when x"1E51",
			x"0000" when x"1E52",
			x"0000" when x"1E53",
			x"0000" when x"1E54",
			x"0000" when x"1E55",
			x"0000" when x"1E56",
			x"0000" when x"1E57",
			x"0000" when x"1E58",
			x"0000" when x"1E59",
			x"0000" when x"1E5A",
			x"0000" when x"1E5B",
			x"0000" when x"1E5C",
			x"0000" when x"1E5D",
			x"0000" when x"1E5E",
			x"0000" when x"1E5F",
			x"0000" when x"1E60",
			x"0000" when x"1E61",
			x"0000" when x"1E62",
			x"0000" when x"1E63",
			x"0000" when x"1E64",
			x"0000" when x"1E65",
			x"0000" when x"1E66",
			x"0000" when x"1E67",
			x"0000" when x"1E68",
			x"0000" when x"1E69",
			x"0000" when x"1E6A",
			x"0000" when x"1E6B",
			x"0000" when x"1E6C",
			x"0000" when x"1E6D",
			x"0000" when x"1E6E",
			x"0000" when x"1E6F",
			x"0000" when x"1E70",
			x"0000" when x"1E71",
			x"0000" when x"1E72",
			x"0000" when x"1E73",
			x"0000" when x"1E74",
			x"0000" when x"1E75",
			x"0000" when x"1E76",
			x"0000" when x"1E77",
			x"0000" when x"1E78",
			x"0000" when x"1E79",
			x"0000" when x"1E7A",
			x"0000" when x"1E7B",
			x"0000" when x"1E7C",
			x"0000" when x"1E7D",
			x"0000" when x"1E7E",
			x"0000" when x"1E7F",
			x"0000" when x"1E80",
			x"0000" when x"1E81",
			x"0000" when x"1E82",
			x"0000" when x"1E83",
			x"0000" when x"1E84",
			x"0000" when x"1E85",
			x"0000" when x"1E86",
			x"0000" when x"1E87",
			x"0000" when x"1E88",
			x"0000" when x"1E89",
			x"0000" when x"1E8A",
			x"0000" when x"1E8B",
			x"0000" when x"1E8C",
			x"0000" when x"1E8D",
			x"0000" when x"1E8E",
			x"0000" when x"1E8F",
			x"0000" when x"1E90",
			x"0000" when x"1E91",
			x"0000" when x"1E92",
			x"0000" when x"1E93",
			x"0000" when x"1E94",
			x"0000" when x"1E95",
			x"0000" when x"1E96",
			x"0000" when x"1E97",
			x"0000" when x"1E98",
			x"0000" when x"1E99",
			x"0000" when x"1E9A",
			x"0000" when x"1E9B",
			x"0000" when x"1E9C",
			x"0000" when x"1E9D",
			x"0000" when x"1E9E",
			x"0000" when x"1E9F",
			x"0000" when x"1EA0",
			x"0000" when x"1EA1",
			x"0000" when x"1EA2",
			x"0000" when x"1EA3",
			x"0000" when x"1EA4",
			x"0000" when x"1EA5",
			x"0000" when x"1EA6",
			x"0000" when x"1EA7",
			x"0000" when x"1EA8",
			x"0000" when x"1EA9",
			x"0000" when x"1EAA",
			x"0000" when x"1EAB",
			x"0000" when x"1EAC",
			x"0000" when x"1EAD",
			x"0000" when x"1EAE",
			x"0000" when x"1EAF",
			x"0000" when x"1EB0",
			x"0000" when x"1EB1",
			x"0000" when x"1EB2",
			x"0000" when x"1EB3",
			x"0000" when x"1EB4",
			x"0000" when x"1EB5",
			x"0000" when x"1EB6",
			x"0000" when x"1EB7",
			x"0000" when x"1EB8",
			x"0000" when x"1EB9",
			x"0000" when x"1EBA",
			x"0000" when x"1EBB",
			x"0000" when x"1EBC",
			x"0000" when x"1EBD",
			x"0000" when x"1EBE",
			x"0000" when x"1EBF",
			x"0000" when x"1EC0",
			x"0000" when x"1EC1",
			x"0000" when x"1EC2",
			x"0000" when x"1EC3",
			x"0000" when x"1EC4",
			x"0000" when x"1EC5",
			x"0000" when x"1EC6",
			x"0000" when x"1EC7",
			x"0000" when x"1EC8",
			x"0000" when x"1EC9",
			x"0000" when x"1ECA",
			x"0000" when x"1ECB",
			x"0000" when x"1ECC",
			x"0000" when x"1ECD",
			x"0000" when x"1ECE",
			x"0000" when x"1ECF",
			x"0000" when x"1ED0",
			x"0000" when x"1ED1",
			x"0000" when x"1ED2",
			x"0000" when x"1ED3",
			x"0000" when x"1ED4",
			x"0000" when x"1ED5",
			x"0000" when x"1ED6",
			x"0000" when x"1ED7",
			x"0000" when x"1ED8",
			x"0000" when x"1ED9",
			x"0000" when x"1EDA",
			x"0000" when x"1EDB",
			x"0000" when x"1EDC",
			x"0000" when x"1EDD",
			x"0000" when x"1EDE",
			x"0000" when x"1EDF",
			x"0000" when x"1EE0",
			x"0000" when x"1EE1",
			x"0000" when x"1EE2",
			x"0000" when x"1EE3",
			x"0000" when x"1EE4",
			x"0000" when x"1EE5",
			x"0000" when x"1EE6",
			x"0000" when x"1EE7",
			x"0000" when x"1EE8",
			x"0000" when x"1EE9",
			x"0000" when x"1EEA",
			x"0000" when x"1EEB",
			x"0000" when x"1EEC",
			x"0000" when x"1EED",
			x"0000" when x"1EEE",
			x"0000" when x"1EEF",
			x"0000" when x"1EF0",
			x"0000" when x"1EF1",
			x"0000" when x"1EF2",
			x"0000" when x"1EF3",
			x"0000" when x"1EF4",
			x"0000" when x"1EF5",
			x"0000" when x"1EF6",
			x"0000" when x"1EF7",
			x"0000" when x"1EF8",
			x"0000" when x"1EF9",
			x"0000" when x"1EFA",
			x"0000" when x"1EFB",
			x"0000" when x"1EFC",
			x"0000" when x"1EFD",
			x"0000" when x"1EFE",
			x"0000" when x"1EFF",
			x"0000" when x"1F00",
			x"0000" when x"1F01",
			x"0000" when x"1F02",
			x"0000" when x"1F03",
			x"0000" when x"1F04",
			x"0000" when x"1F05",
			x"0000" when x"1F06",
			x"0000" when x"1F07",
			x"0000" when x"1F08",
			x"0000" when x"1F09",
			x"0000" when x"1F0A",
			x"0000" when x"1F0B",
			x"0000" when x"1F0C",
			x"0000" when x"1F0D",
			x"0000" when x"1F0E",
			x"0000" when x"1F0F",
			x"0000" when x"1F10",
			x"0000" when x"1F11",
			x"0000" when x"1F12",
			x"0000" when x"1F13",
			x"0000" when x"1F14",
			x"0000" when x"1F15",
			x"0000" when x"1F16",
			x"0000" when x"1F17",
			x"0000" when x"1F18",
			x"0000" when x"1F19",
			x"0000" when x"1F1A",
			x"0000" when x"1F1B",
			x"0000" when x"1F1C",
			x"0000" when x"1F1D",
			x"0000" when x"1F1E",
			x"0000" when x"1F1F",
			x"0000" when x"1F20",
			x"0000" when x"1F21",
			x"0000" when x"1F22",
			x"0000" when x"1F23",
			x"0000" when x"1F24",
			x"0000" when x"1F25",
			x"0000" when x"1F26",
			x"0000" when x"1F27",
			x"0000" when x"1F28",
			x"0000" when x"1F29",
			x"0000" when x"1F2A",
			x"0000" when x"1F2B",
			x"0000" when x"1F2C",
			x"0000" when x"1F2D",
			x"0000" when x"1F2E",
			x"0000" when x"1F2F",
			x"0000" when x"1F30",
			x"0000" when x"1F31",
			x"0000" when x"1F32",
			x"0000" when x"1F33",
			x"0000" when x"1F34",
			x"0000" when x"1F35",
			x"0000" when x"1F36",
			x"0000" when x"1F37",
			x"0000" when x"1F38",
			x"0000" when x"1F39",
			x"0000" when x"1F3A",
			x"0000" when x"1F3B",
			x"0000" when x"1F3C",
			x"0000" when x"1F3D",
			x"0000" when x"1F3E",
			x"0000" when x"1F3F",
			x"0000" when x"1F40",
			x"0000" when x"1F41",
			x"0000" when x"1F42",
			x"0000" when x"1F43",
			x"0000" when x"1F44",
			x"0000" when x"1F45",
			x"0000" when x"1F46",
			x"0000" when x"1F47",
			x"0000" when x"1F48",
			x"0000" when x"1F49",
			x"0000" when x"1F4A",
			x"0000" when x"1F4B",
			x"0000" when x"1F4C",
			x"0000" when x"1F4D",
			x"0000" when x"1F4E",
			x"0000" when x"1F4F",
			x"0000" when x"1F50",
			x"0000" when x"1F51",
			x"0000" when x"1F52",
			x"0000" when x"1F53",
			x"0000" when x"1F54",
			x"0000" when x"1F55",
			x"0000" when x"1F56",
			x"0000" when x"1F57",
			x"0000" when x"1F58",
			x"0000" when x"1F59",
			x"0000" when x"1F5A",
			x"0000" when x"1F5B",
			x"0000" when x"1F5C",
			x"0000" when x"1F5D",
			x"0000" when x"1F5E",
			x"0000" when x"1F5F",
			x"0000" when x"1F60",
			x"0000" when x"1F61",
			x"0000" when x"1F62",
			x"0000" when x"1F63",
			x"0000" when x"1F64",
			x"0000" when x"1F65",
			x"0000" when x"1F66",
			x"0000" when x"1F67",
			x"0000" when x"1F68",
			x"0000" when x"1F69",
			x"0000" when x"1F6A",
			x"0000" when x"1F6B",
			x"0000" when x"1F6C",
			x"0000" when x"1F6D",
			x"0000" when x"1F6E",
			x"0000" when x"1F6F",
			x"0000" when x"1F70",
			x"0000" when x"1F71",
			x"0000" when x"1F72",
			x"0000" when x"1F73",
			x"0000" when x"1F74",
			x"0000" when x"1F75",
			x"0000" when x"1F76",
			x"0000" when x"1F77",
			x"0000" when x"1F78",
			x"0000" when x"1F79",
			x"0000" when x"1F7A",
			x"0000" when x"1F7B",
			x"0000" when x"1F7C",
			x"0000" when x"1F7D",
			x"0000" when x"1F7E",
			x"0000" when x"1F7F",
			x"0000" when x"1F80",
			x"0000" when x"1F81",
			x"0000" when x"1F82",
			x"0000" when x"1F83",
			x"0000" when x"1F84",
			x"0000" when x"1F85",
			x"0000" when x"1F86",
			x"0000" when x"1F87",
			x"0000" when x"1F88",
			x"0000" when x"1F89",
			x"0000" when x"1F8A",
			x"0000" when x"1F8B",
			x"0000" when x"1F8C",
			x"0000" when x"1F8D",
			x"0000" when x"1F8E",
			x"0000" when x"1F8F",
			x"0000" when x"1F90",
			x"0000" when x"1F91",
			x"0000" when x"1F92",
			x"0000" when x"1F93",
			x"0000" when x"1F94",
			x"0000" when x"1F95",
			x"0000" when x"1F96",
			x"0000" when x"1F97",
			x"0000" when x"1F98",
			x"0000" when x"1F99",
			x"0000" when x"1F9A",
			x"0000" when x"1F9B",
			x"0000" when x"1F9C",
			x"0000" when x"1F9D",
			x"0000" when x"1F9E",
			x"0000" when x"1F9F",
			x"0000" when x"1FA0",
			x"0000" when x"1FA1",
			x"0000" when x"1FA2",
			x"0000" when x"1FA3",
			x"0000" when x"1FA4",
			x"0000" when x"1FA5",
			x"0000" when x"1FA6",
			x"0000" when x"1FA7",
			x"0000" when x"1FA8",
			x"0000" when x"1FA9",
			x"0000" when x"1FAA",
			x"0000" when x"1FAB",
			x"0000" when x"1FAC",
			x"0000" when x"1FAD",
			x"0000" when x"1FAE",
			x"0000" when x"1FAF",
			x"0000" when x"1FB0",
			x"0000" when x"1FB1",
			x"0000" when x"1FB2",
			x"0000" when x"1FB3",
			x"0000" when x"1FB4",
			x"0000" when x"1FB5",
			x"0000" when x"1FB6",
			x"0000" when x"1FB7",
			x"0000" when x"1FB8",
			x"0000" when x"1FB9",
			x"0000" when x"1FBA",
			x"0000" when x"1FBB",
			x"0000" when x"1FBC",
			x"0000" when x"1FBD",
			x"0000" when x"1FBE",
			x"0000" when x"1FBF",
			x"0000" when x"1FC0",
			x"0000" when x"1FC1",
			x"0000" when x"1FC2",
			x"0000" when x"1FC3",
			x"0000" when x"1FC4",
			x"0000" when x"1FC5",
			x"0000" when x"1FC6",
			x"0000" when x"1FC7",
			x"0000" when x"1FC8",
			x"0000" when x"1FC9",
			x"0000" when x"1FCA",
			x"0000" when x"1FCB",
			x"0000" when x"1FCC",
			x"0000" when x"1FCD",
			x"0000" when x"1FCE",
			x"0000" when x"1FCF",
			x"0000" when x"1FD0",
			x"0000" when x"1FD1",
			x"0000" when x"1FD2",
			x"0000" when x"1FD3",
			x"0000" when x"1FD4",
			x"0000" when x"1FD5",
			x"0000" when x"1FD6",
			x"0000" when x"1FD7",
			x"0000" when x"1FD8",
			x"0000" when x"1FD9",
			x"0000" when x"1FDA",
			x"0000" when x"1FDB",
			x"0000" when x"1FDC",
			x"0000" when x"1FDD",
			x"0000" when x"1FDE",
			x"0000" when x"1FDF",
			x"0000" when x"1FE0",
			x"0000" when x"1FE1",
			x"0000" when x"1FE2",
			x"0000" when x"1FE3",
			x"0000" when x"1FE4",
			x"0000" when x"1FE5",
			x"0000" when x"1FE6",
			x"0000" when x"1FE7",
			x"0000" when x"1FE8",
			x"0000" when x"1FE9",
			x"0000" when x"1FEA",
			x"0000" when x"1FEB",
			x"0000" when x"1FEC",
			x"0000" when x"1FED",
			x"0000" when x"1FEE",
			x"0000" when x"1FEF",
			x"0000" when x"1FF0",
			x"0000" when x"1FF1",
			x"0000" when x"1FF2",
			x"0000" when x"1FF3",
			x"0000" when x"1FF4",
			x"0000" when x"1FF5",
			x"0000" when x"1FF6",
			x"0000" when x"1FF7",
			x"0000" when x"1FF8",
			x"0000" when x"1FF9",
			x"0000" when x"1FFA",
			x"0000" when x"1FFB",
			x"0000" when x"1FFC",
			x"0000" when x"1FFD",
			x"0000" when x"1FFE",
			x"0000" when x"1FFF",
			x"0000" when x"2000",
			x"0000" when x"2001",
			x"0000" when x"2002",
			x"0000" when x"2003",
			x"0000" when x"2004",
			x"0000" when x"2005",
			x"0000" when x"2006",
			x"0000" when x"2007",
			x"0000" when x"2008",
			x"0000" when x"2009",
			x"0000" when x"200A",
			x"0000" when x"200B",
			x"0000" when x"200C",
			x"0000" when x"200D",
			x"0000" when x"200E",
			x"0000" when x"200F",
			x"0000" when x"2010",
			x"0000" when x"2011",
			x"0000" when x"2012",
			x"0000" when x"2013",
			x"0000" when x"2014",
			x"0000" when x"2015",
			x"0000" when x"2016",
			x"0000" when x"2017",
			x"0000" when x"2018",
			x"0000" when x"2019",
			x"0000" when x"201A",
			x"0000" when x"201B",
			x"0000" when x"201C",
			x"0000" when x"201D",
			x"0000" when x"201E",
			x"0000" when x"201F",
			x"0000" when x"2020",
			x"0000" when x"2021",
			x"0000" when x"2022",
			x"0000" when x"2023",
			x"0000" when x"2024",
			x"0000" when x"2025",
			x"0000" when x"2026",
			x"0000" when x"2027",
			x"0000" when x"2028",
			x"0000" when x"2029",
			x"0000" when x"202A",
			x"0000" when x"202B",
			x"0000" when x"202C",
			x"0000" when x"202D",
			x"0000" when x"202E",
			x"0000" when x"202F",
			x"0000" when x"2030",
			x"0000" when x"2031",
			x"0000" when x"2032",
			x"0000" when x"2033",
			x"0000" when x"2034",
			x"0000" when x"2035",
			x"0000" when x"2036",
			x"0000" when x"2037",
			x"0000" when x"2038",
			x"0000" when x"2039",
			x"0000" when x"203A",
			x"0000" when x"203B",
			x"0000" when x"203C",
			x"0000" when x"203D",
			x"0000" when x"203E",
			x"0000" when x"203F",
			x"0000" when x"2040",
			x"0000" when x"2041",
			x"0000" when x"2042",
			x"0000" when x"2043",
			x"0000" when x"2044",
			x"0000" when x"2045",
			x"0000" when x"2046",
			x"0000" when x"2047",
			x"0000" when x"2048",
			x"0000" when x"2049",
			x"0000" when x"204A",
			x"0000" when x"204B",
			x"0000" when x"204C",
			x"0000" when x"204D",
			x"0000" when x"204E",
			x"0000" when x"204F",
			x"0000" when x"2050",
			x"0000" when x"2051",
			x"0000" when x"2052",
			x"0000" when x"2053",
			x"0000" when x"2054",
			x"0000" when x"2055",
			x"0000" when x"2056",
			x"0000" when x"2057",
			x"0000" when x"2058",
			x"0000" when x"2059",
			x"0000" when x"205A",
			x"0000" when x"205B",
			x"0000" when x"205C",
			x"0000" when x"205D",
			x"0000" when x"205E",
			x"0000" when x"205F",
			x"0000" when x"2060",
			x"0000" when x"2061",
			x"0000" when x"2062",
			x"0000" when x"2063",
			x"0000" when x"2064",
			x"0000" when x"2065",
			x"0000" when x"2066",
			x"0000" when x"2067",
			x"0000" when x"2068",
			x"0000" when x"2069",
			x"0000" when x"206A",
			x"0000" when x"206B",
			x"0000" when x"206C",
			x"0000" when x"206D",
			x"0000" when x"206E",
			x"0000" when x"206F",
			x"0000" when x"2070",
			x"0000" when x"2071",
			x"0000" when x"2072",
			x"0000" when x"2073",
			x"0000" when x"2074",
			x"0000" when x"2075",
			x"0000" when x"2076",
			x"0000" when x"2077",
			x"0000" when x"2078",
			x"0000" when x"2079",
			x"0000" when x"207A",
			x"0000" when x"207B",
			x"0000" when x"207C",
			x"0000" when x"207D",
			x"0000" when x"207E",
			x"0000" when x"207F",
			x"0000" when x"2080",
			x"0000" when x"2081",
			x"0000" when x"2082",
			x"0000" when x"2083",
			x"0000" when x"2084",
			x"0000" when x"2085",
			x"0000" when x"2086",
			x"0000" when x"2087",
			x"0000" when x"2088",
			x"0000" when x"2089",
			x"0000" when x"208A",
			x"0000" when x"208B",
			x"0000" when x"208C",
			x"0000" when x"208D",
			x"0000" when x"208E",
			x"0000" when x"208F",
			x"0000" when x"2090",
			x"0000" when x"2091",
			x"0000" when x"2092",
			x"0000" when x"2093",
			x"0000" when x"2094",
			x"0000" when x"2095",
			x"0000" when x"2096",
			x"0000" when x"2097",
			x"0000" when x"2098",
			x"0000" when x"2099",
			x"0000" when x"209A",
			x"0000" when x"209B",
			x"0000" when x"209C",
			x"0000" when x"209D",
			x"0000" when x"209E",
			x"0000" when x"209F",
			x"0000" when x"20A0",
			x"0000" when x"20A1",
			x"0000" when x"20A2",
			x"0000" when x"20A3",
			x"0000" when x"20A4",
			x"0000" when x"20A5",
			x"0000" when x"20A6",
			x"0000" when x"20A7",
			x"0000" when x"20A8",
			x"0000" when x"20A9",
			x"0000" when x"20AA",
			x"0000" when x"20AB",
			x"0000" when x"20AC",
			x"0000" when x"20AD",
			x"0000" when x"20AE",
			x"0000" when x"20AF",
			x"0000" when x"20B0",
			x"0000" when x"20B1",
			x"0000" when x"20B2",
			x"0000" when x"20B3",
			x"0000" when x"20B4",
			x"0000" when x"20B5",
			x"0000" when x"20B6",
			x"0000" when x"20B7",
			x"0000" when x"20B8",
			x"0000" when x"20B9",
			x"0000" when x"20BA",
			x"0000" when x"20BB",
			x"0000" when x"20BC",
			x"0000" when x"20BD",
			x"0000" when x"20BE",
			x"0000" when x"20BF",
			x"0000" when x"20C0",
			x"0000" when x"20C1",
			x"0000" when x"20C2",
			x"0000" when x"20C3",
			x"0000" when x"20C4",
			x"0000" when x"20C5",
			x"0000" when x"20C6",
			x"0000" when x"20C7",
			x"0000" when x"20C8",
			x"0000" when x"20C9",
			x"0000" when x"20CA",
			x"0000" when x"20CB",
			x"0000" when x"20CC",
			x"0000" when x"20CD",
			x"0000" when x"20CE",
			x"0000" when x"20CF",
			x"0000" when x"20D0",
			x"0000" when x"20D1",
			x"0000" when x"20D2",
			x"0000" when x"20D3",
			x"0000" when x"20D4",
			x"0000" when x"20D5",
			x"0000" when x"20D6",
			x"0000" when x"20D7",
			x"0000" when x"20D8",
			x"0000" when x"20D9",
			x"0000" when x"20DA",
			x"0000" when x"20DB",
			x"0000" when x"20DC",
			x"0000" when x"20DD",
			x"0000" when x"20DE",
			x"0000" when x"20DF",
			x"0000" when x"20E0",
			x"0000" when x"20E1",
			x"0000" when x"20E2",
			x"0000" when x"20E3",
			x"0000" when x"20E4",
			x"0000" when x"20E5",
			x"0000" when x"20E6",
			x"0000" when x"20E7",
			x"0000" when x"20E8",
			x"0000" when x"20E9",
			x"0000" when x"20EA",
			x"0000" when x"20EB",
			x"0000" when x"20EC",
			x"0000" when x"20ED",
			x"0000" when x"20EE",
			x"0000" when x"20EF",
			x"0000" when x"20F0",
			x"0000" when x"20F1",
			x"0000" when x"20F2",
			x"0000" when x"20F3",
			x"0000" when x"20F4",
			x"0000" when x"20F5",
			x"0000" when x"20F6",
			x"0000" when x"20F7",
			x"0000" when x"20F8",
			x"0000" when x"20F9",
			x"0000" when x"20FA",
			x"0000" when x"20FB",
			x"0000" when x"20FC",
			x"0000" when x"20FD",
			x"0000" when x"20FE",
			x"0000" when x"20FF",
			x"0000" when x"2100",
			x"0000" when x"2101",
			x"0000" when x"2102",
			x"0000" when x"2103",
			x"0000" when x"2104",
			x"0000" when x"2105",
			x"0000" when x"2106",
			x"0000" when x"2107",
			x"0000" when x"2108",
			x"0000" when x"2109",
			x"0000" when x"210A",
			x"0000" when x"210B",
			x"0000" when x"210C",
			x"0000" when x"210D",
			x"0000" when x"210E",
			x"0000" when x"210F",
			x"0000" when x"2110",
			x"0000" when x"2111",
			x"0000" when x"2112",
			x"0000" when x"2113",
			x"0000" when x"2114",
			x"0000" when x"2115",
			x"0000" when x"2116",
			x"0000" when x"2117",
			x"0000" when x"2118",
			x"0000" when x"2119",
			x"0000" when x"211A",
			x"0000" when x"211B",
			x"0000" when x"211C",
			x"0000" when x"211D",
			x"0000" when x"211E",
			x"0000" when x"211F",
			x"0000" when x"2120",
			x"0000" when x"2121",
			x"0000" when x"2122",
			x"0000" when x"2123",
			x"0000" when x"2124",
			x"0000" when x"2125",
			x"0000" when x"2126",
			x"0000" when x"2127",
			x"0000" when x"2128",
			x"0000" when x"2129",
			x"0000" when x"212A",
			x"0000" when x"212B",
			x"0000" when x"212C",
			x"0000" when x"212D",
			x"0000" when x"212E",
			x"0000" when x"212F",
			x"0000" when x"2130",
			x"0000" when x"2131",
			x"0000" when x"2132",
			x"0000" when x"2133",
			x"0000" when x"2134",
			x"0000" when x"2135",
			x"0000" when x"2136",
			x"0000" when x"2137",
			x"0000" when x"2138",
			x"0000" when x"2139",
			x"0000" when x"213A",
			x"0000" when x"213B",
			x"0000" when x"213C",
			x"0000" when x"213D",
			x"0000" when x"213E",
			x"0000" when x"213F",
			x"0000" when x"2140",
			x"0000" when x"2141",
			x"0000" when x"2142",
			x"0000" when x"2143",
			x"0000" when x"2144",
			x"0000" when x"2145",
			x"0000" when x"2146",
			x"0000" when x"2147",
			x"0000" when x"2148",
			x"0000" when x"2149",
			x"0000" when x"214A",
			x"0000" when x"214B",
			x"0000" when x"214C",
			x"0000" when x"214D",
			x"0000" when x"214E",
			x"0000" when x"214F",
			x"0000" when x"2150",
			x"0000" when x"2151",
			x"0000" when x"2152",
			x"0000" when x"2153",
			x"0000" when x"2154",
			x"0000" when x"2155",
			x"0000" when x"2156",
			x"0000" when x"2157",
			x"0000" when x"2158",
			x"0000" when x"2159",
			x"0000" when x"215A",
			x"0000" when x"215B",
			x"0000" when x"215C",
			x"0000" when x"215D",
			x"0000" when x"215E",
			x"0000" when x"215F",
			x"0000" when x"2160",
			x"0000" when x"2161",
			x"0000" when x"2162",
			x"0000" when x"2163",
			x"0000" when x"2164",
			x"0000" when x"2165",
			x"0000" when x"2166",
			x"0000" when x"2167",
			x"0000" when x"2168",
			x"0000" when x"2169",
			x"0000" when x"216A",
			x"0000" when x"216B",
			x"0000" when x"216C",
			x"0000" when x"216D",
			x"0000" when x"216E",
			x"0000" when x"216F",
			x"0000" when x"2170",
			x"0000" when x"2171",
			x"0000" when x"2172",
			x"0000" when x"2173",
			x"0000" when x"2174",
			x"0000" when x"2175",
			x"0000" when x"2176",
			x"0000" when x"2177",
			x"0000" when x"2178",
			x"0000" when x"2179",
			x"0000" when x"217A",
			x"0000" when x"217B",
			x"0000" when x"217C",
			x"0000" when x"217D",
			x"0000" when x"217E",
			x"0000" when x"217F",
			x"0000" when x"2180",
			x"0000" when x"2181",
			x"0000" when x"2182",
			x"0000" when x"2183",
			x"0000" when x"2184",
			x"0000" when x"2185",
			x"0000" when x"2186",
			x"0000" when x"2187",
			x"0000" when x"2188",
			x"0000" when x"2189",
			x"0000" when x"218A",
			x"0000" when x"218B",
			x"0000" when x"218C",
			x"0000" when x"218D",
			x"0000" when x"218E",
			x"0000" when x"218F",
			x"0000" when x"2190",
			x"0000" when x"2191",
			x"0000" when x"2192",
			x"0000" when x"2193",
			x"0000" when x"2194",
			x"0000" when x"2195",
			x"0000" when x"2196",
			x"0000" when x"2197",
			x"0000" when x"2198",
			x"0000" when x"2199",
			x"0000" when x"219A",
			x"0000" when x"219B",
			x"0000" when x"219C",
			x"0000" when x"219D",
			x"0000" when x"219E",
			x"0000" when x"219F",
			x"0000" when x"21A0",
			x"0000" when x"21A1",
			x"0000" when x"21A2",
			x"0000" when x"21A3",
			x"0000" when x"21A4",
			x"0000" when x"21A5",
			x"0000" when x"21A6",
			x"0000" when x"21A7",
			x"0000" when x"21A8",
			x"0000" when x"21A9",
			x"0000" when x"21AA",
			x"0000" when x"21AB",
			x"0000" when x"21AC",
			x"0000" when x"21AD",
			x"0000" when x"21AE",
			x"0000" when x"21AF",
			x"0000" when x"21B0",
			x"0000" when x"21B1",
			x"0000" when x"21B2",
			x"0000" when x"21B3",
			x"0000" when x"21B4",
			x"0000" when x"21B5",
			x"0000" when x"21B6",
			x"0000" when x"21B7",
			x"0000" when x"21B8",
			x"0000" when x"21B9",
			x"0000" when x"21BA",
			x"0000" when x"21BB",
			x"0000" when x"21BC",
			x"0000" when x"21BD",
			x"0000" when x"21BE",
			x"0000" when x"21BF",
			x"0000" when x"21C0",
			x"0000" when x"21C1",
			x"0000" when x"21C2",
			x"0000" when x"21C3",
			x"0000" when x"21C4",
			x"0000" when x"21C5",
			x"0000" when x"21C6",
			x"0000" when x"21C7",
			x"0000" when x"21C8",
			x"0000" when x"21C9",
			x"0000" when x"21CA",
			x"0000" when x"21CB",
			x"0000" when x"21CC",
			x"0000" when x"21CD",
			x"0000" when x"21CE",
			x"0000" when x"21CF",
			x"0000" when x"21D0",
			x"0000" when x"21D1",
			x"0000" when x"21D2",
			x"0000" when x"21D3",
			x"0000" when x"21D4",
			x"0000" when x"21D5",
			x"0000" when x"21D6",
			x"0000" when x"21D7",
			x"0000" when x"21D8",
			x"0000" when x"21D9",
			x"0000" when x"21DA",
			x"0000" when x"21DB",
			x"0000" when x"21DC",
			x"0000" when x"21DD",
			x"0000" when x"21DE",
			x"0000" when x"21DF",
			x"0000" when x"21E0",
			x"0000" when x"21E1",
			x"0000" when x"21E2",
			x"0000" when x"21E3",
			x"0000" when x"21E4",
			x"0000" when x"21E5",
			x"0000" when x"21E6",
			x"0000" when x"21E7",
			x"0000" when x"21E8",
			x"0000" when x"21E9",
			x"0000" when x"21EA",
			x"0000" when x"21EB",
			x"0000" when x"21EC",
			x"0000" when x"21ED",
			x"0000" when x"21EE",
			x"0000" when x"21EF",
			x"0000" when x"21F0",
			x"0000" when x"21F1",
			x"0000" when x"21F2",
			x"0000" when x"21F3",
			x"0000" when x"21F4",
			x"0000" when x"21F5",
			x"0000" when x"21F6",
			x"0000" when x"21F7",
			x"0000" when x"21F8",
			x"0000" when x"21F9",
			x"0000" when x"21FA",
			x"0000" when x"21FB",
			x"0000" when x"21FC",
			x"0000" when x"21FD",
			x"0000" when x"21FE",
			x"0000" when x"21FF",
			x"0000" when x"2200",
			x"0000" when x"2201",
			x"0000" when x"2202",
			x"0000" when x"2203",
			x"0000" when x"2204",
			x"0000" when x"2205",
			x"0000" when x"2206",
			x"0000" when x"2207",
			x"0000" when x"2208",
			x"0000" when x"2209",
			x"0000" when x"220A",
			x"0000" when x"220B",
			x"0000" when x"220C",
			x"0000" when x"220D",
			x"0000" when x"220E",
			x"0000" when x"220F",
			x"0000" when x"2210",
			x"0000" when x"2211",
			x"0000" when x"2212",
			x"0000" when x"2213",
			x"0000" when x"2214",
			x"0000" when x"2215",
			x"0000" when x"2216",
			x"0000" when x"2217",
			x"0000" when x"2218",
			x"0000" when x"2219",
			x"0000" when x"221A",
			x"0000" when x"221B",
			x"0000" when x"221C",
			x"0000" when x"221D",
			x"0000" when x"221E",
			x"0000" when x"221F",
			x"0000" when x"2220",
			x"0000" when x"2221",
			x"0000" when x"2222",
			x"0000" when x"2223",
			x"0000" when x"2224",
			x"0000" when x"2225",
			x"0000" when x"2226",
			x"0000" when x"2227",
			x"0000" when x"2228",
			x"0000" when x"2229",
			x"0000" when x"222A",
			x"0000" when x"222B",
			x"0000" when x"222C",
			x"0000" when x"222D",
			x"0000" when x"222E",
			x"0000" when x"222F",
			x"0000" when x"2230",
			x"0000" when x"2231",
			x"0000" when x"2232",
			x"0000" when x"2233",
			x"0000" when x"2234",
			x"0000" when x"2235",
			x"0000" when x"2236",
			x"0000" when x"2237",
			x"0000" when x"2238",
			x"0000" when x"2239",
			x"0000" when x"223A",
			x"0000" when x"223B",
			x"0000" when x"223C",
			x"0000" when x"223D",
			x"0000" when x"223E",
			x"0000" when x"223F",
			x"0000" when x"2240",
			x"0000" when x"2241",
			x"0000" when x"2242",
			x"0000" when x"2243",
			x"0000" when x"2244",
			x"0000" when x"2245",
			x"0000" when x"2246",
			x"0000" when x"2247",
			x"0000" when x"2248",
			x"0000" when x"2249",
			x"0000" when x"224A",
			x"0000" when x"224B",
			x"0000" when x"224C",
			x"0000" when x"224D",
			x"0000" when x"224E",
			x"0000" when x"224F",
			x"0000" when x"2250",
			x"0000" when x"2251",
			x"0000" when x"2252",
			x"0000" when x"2253",
			x"0000" when x"2254",
			x"0000" when x"2255",
			x"0000" when x"2256",
			x"0000" when x"2257",
			x"0000" when x"2258",
			x"0000" when x"2259",
			x"0000" when x"225A",
			x"0000" when x"225B",
			x"0000" when x"225C",
			x"0000" when x"225D",
			x"0000" when x"225E",
			x"0000" when x"225F",
			x"0000" when x"2260",
			x"0000" when x"2261",
			x"0000" when x"2262",
			x"0000" when x"2263",
			x"0000" when x"2264",
			x"0000" when x"2265",
			x"0000" when x"2266",
			x"0000" when x"2267",
			x"0000" when x"2268",
			x"0000" when x"2269",
			x"0000" when x"226A",
			x"0000" when x"226B",
			x"0000" when x"226C",
			x"0000" when x"226D",
			x"0000" when x"226E",
			x"0000" when x"226F",
			x"0000" when x"2270",
			x"0000" when x"2271",
			x"0000" when x"2272",
			x"0000" when x"2273",
			x"0000" when x"2274",
			x"0000" when x"2275",
			x"0000" when x"2276",
			x"0000" when x"2277",
			x"0000" when x"2278",
			x"0000" when x"2279",
			x"0000" when x"227A",
			x"0000" when x"227B",
			x"0000" when x"227C",
			x"0000" when x"227D",
			x"0000" when x"227E",
			x"0000" when x"227F",
			x"0000" when x"2280",
			x"0000" when x"2281",
			x"0000" when x"2282",
			x"0000" when x"2283",
			x"0000" when x"2284",
			x"0000" when x"2285",
			x"0000" when x"2286",
			x"0000" when x"2287",
			x"0000" when x"2288",
			x"0000" when x"2289",
			x"0000" when x"228A",
			x"0000" when x"228B",
			x"0000" when x"228C",
			x"0000" when x"228D",
			x"0000" when x"228E",
			x"0000" when x"228F",
			x"0000" when x"2290",
			x"0000" when x"2291",
			x"0000" when x"2292",
			x"0000" when x"2293",
			x"0000" when x"2294",
			x"0000" when x"2295",
			x"0000" when x"2296",
			x"0000" when x"2297",
			x"0000" when x"2298",
			x"0000" when x"2299",
			x"0000" when x"229A",
			x"0000" when x"229B",
			x"0000" when x"229C",
			x"0000" when x"229D",
			x"0000" when x"229E",
			x"0000" when x"229F",
			x"0000" when x"22A0",
			x"0000" when x"22A1",
			x"0000" when x"22A2",
			x"0000" when x"22A3",
			x"0000" when x"22A4",
			x"0000" when x"22A5",
			x"0000" when x"22A6",
			x"0000" when x"22A7",
			x"0000" when x"22A8",
			x"0000" when x"22A9",
			x"0000" when x"22AA",
			x"0000" when x"22AB",
			x"0000" when x"22AC",
			x"0000" when x"22AD",
			x"0000" when x"22AE",
			x"0000" when x"22AF",
			x"0000" when x"22B0",
			x"0000" when x"22B1",
			x"0000" when x"22B2",
			x"0000" when x"22B3",
			x"0000" when x"22B4",
			x"0000" when x"22B5",
			x"0000" when x"22B6",
			x"0000" when x"22B7",
			x"0000" when x"22B8",
			x"0000" when x"22B9",
			x"0000" when x"22BA",
			x"0000" when x"22BB",
			x"0000" when x"22BC",
			x"0000" when x"22BD",
			x"0000" when x"22BE",
			x"0000" when x"22BF",
			x"0000" when x"22C0",
			x"0000" when x"22C1",
			x"0000" when x"22C2",
			x"0000" when x"22C3",
			x"0000" when x"22C4",
			x"0000" when x"22C5",
			x"0000" when x"22C6",
			x"0000" when x"22C7",
			x"0000" when x"22C8",
			x"0000" when x"22C9",
			x"0000" when x"22CA",
			x"0000" when x"22CB",
			x"0000" when x"22CC",
			x"0000" when x"22CD",
			x"0000" when x"22CE",
			x"0000" when x"22CF",
			x"0000" when x"22D0",
			x"0000" when x"22D1",
			x"0000" when x"22D2",
			x"0000" when x"22D3",
			x"0000" when x"22D4",
			x"0000" when x"22D5",
			x"0000" when x"22D6",
			x"0000" when x"22D7",
			x"0000" when x"22D8",
			x"0000" when x"22D9",
			x"0000" when x"22DA",
			x"0000" when x"22DB",
			x"0000" when x"22DC",
			x"0000" when x"22DD",
			x"0000" when x"22DE",
			x"0000" when x"22DF",
			x"0000" when x"22E0",
			x"0000" when x"22E1",
			x"0000" when x"22E2",
			x"0000" when x"22E3",
			x"0000" when x"22E4",
			x"0000" when x"22E5",
			x"0000" when x"22E6",
			x"0000" when x"22E7",
			x"0000" when x"22E8",
			x"0000" when x"22E9",
			x"0000" when x"22EA",
			x"0000" when x"22EB",
			x"0000" when x"22EC",
			x"0000" when x"22ED",
			x"0000" when x"22EE",
			x"0000" when x"22EF",
			x"0000" when x"22F0",
			x"0000" when x"22F1",
			x"0000" when x"22F2",
			x"0000" when x"22F3",
			x"0000" when x"22F4",
			x"0000" when x"22F5",
			x"0000" when x"22F6",
			x"0000" when x"22F7",
			x"0000" when x"22F8",
			x"0000" when x"22F9",
			x"0000" when x"22FA",
			x"0000" when x"22FB",
			x"0000" when x"22FC",
			x"0000" when x"22FD",
			x"0000" when x"22FE",
			x"0000" when x"22FF",
			x"0000" when x"2300",
			x"0000" when x"2301",
			x"0000" when x"2302",
			x"0000" when x"2303",
			x"0000" when x"2304",
			x"0000" when x"2305",
			x"0000" when x"2306",
			x"0000" when x"2307",
			x"0000" when x"2308",
			x"0000" when x"2309",
			x"0000" when x"230A",
			x"0000" when x"230B",
			x"0000" when x"230C",
			x"0000" when x"230D",
			x"0000" when x"230E",
			x"0000" when x"230F",
			x"0000" when x"2310",
			x"0000" when x"2311",
			x"0000" when x"2312",
			x"0000" when x"2313",
			x"0000" when x"2314",
			x"0000" when x"2315",
			x"0000" when x"2316",
			x"0000" when x"2317",
			x"0000" when x"2318",
			x"0000" when x"2319",
			x"0000" when x"231A",
			x"0000" when x"231B",
			x"0000" when x"231C",
			x"0000" when x"231D",
			x"0000" when x"231E",
			x"0000" when x"231F",
			x"0000" when x"2320",
			x"0000" when x"2321",
			x"0000" when x"2322",
			x"0000" when x"2323",
			x"0000" when x"2324",
			x"0000" when x"2325",
			x"0000" when x"2326",
			x"0000" when x"2327",
			x"0000" when x"2328",
			x"0000" when x"2329",
			x"0000" when x"232A",
			x"0000" when x"232B",
			x"0000" when x"232C",
			x"0000" when x"232D",
			x"0000" when x"232E",
			x"0000" when x"232F",
			x"0000" when x"2330",
			x"0000" when x"2331",
			x"0000" when x"2332",
			x"0000" when x"2333",
			x"0000" when x"2334",
			x"0000" when x"2335",
			x"0000" when x"2336",
			x"0000" when x"2337",
			x"0000" when x"2338",
			x"0000" when x"2339",
			x"0000" when x"233A",
			x"0000" when x"233B",
			x"0000" when x"233C",
			x"0000" when x"233D",
			x"0000" when x"233E",
			x"0000" when x"233F",
			x"0000" when x"2340",
			x"0000" when x"2341",
			x"0000" when x"2342",
			x"0000" when x"2343",
			x"0000" when x"2344",
			x"0000" when x"2345",
			x"0000" when x"2346",
			x"0000" when x"2347",
			x"0000" when x"2348",
			x"0000" when x"2349",
			x"0000" when x"234A",
			x"0000" when x"234B",
			x"0000" when x"234C",
			x"0000" when x"234D",
			x"0000" when x"234E",
			x"0000" when x"234F",
			x"0000" when x"2350",
			x"0000" when x"2351",
			x"0000" when x"2352",
			x"0000" when x"2353",
			x"0000" when x"2354",
			x"0000" when x"2355",
			x"0000" when x"2356",
			x"0000" when x"2357",
			x"0000" when x"2358",
			x"0000" when x"2359",
			x"0000" when x"235A",
			x"0000" when x"235B",
			x"0000" when x"235C",
			x"0000" when x"235D",
			x"0000" when x"235E",
			x"0000" when x"235F",
			x"0000" when x"2360",
			x"0000" when x"2361",
			x"0000" when x"2362",
			x"0000" when x"2363",
			x"0000" when x"2364",
			x"0000" when x"2365",
			x"0000" when x"2366",
			x"0000" when x"2367",
			x"0000" when x"2368",
			x"0000" when x"2369",
			x"0000" when x"236A",
			x"0000" when x"236B",
			x"0000" when x"236C",
			x"0000" when x"236D",
			x"0000" when x"236E",
			x"0000" when x"236F",
			x"0000" when x"2370",
			x"0000" when x"2371",
			x"0000" when x"2372",
			x"0000" when x"2373",
			x"0000" when x"2374",
			x"0000" when x"2375",
			x"0000" when x"2376",
			x"0000" when x"2377",
			x"0000" when x"2378",
			x"0000" when x"2379",
			x"0000" when x"237A",
			x"0000" when x"237B",
			x"0000" when x"237C",
			x"0000" when x"237D",
			x"0000" when x"237E",
			x"0000" when x"237F",
			x"0000" when x"2380",
			x"0000" when x"2381",
			x"0000" when x"2382",
			x"0000" when x"2383",
			x"0000" when x"2384",
			x"0000" when x"2385",
			x"0000" when x"2386",
			x"0000" when x"2387",
			x"0000" when x"2388",
			x"0000" when x"2389",
			x"0000" when x"238A",
			x"0000" when x"238B",
			x"0000" when x"238C",
			x"0000" when x"238D",
			x"0000" when x"238E",
			x"0000" when x"238F",
			x"0000" when x"2390",
			x"0000" when x"2391",
			x"0000" when x"2392",
			x"0000" when x"2393",
			x"0000" when x"2394",
			x"0000" when x"2395",
			x"0000" when x"2396",
			x"0000" when x"2397",
			x"0000" when x"2398",
			x"0000" when x"2399",
			x"0000" when x"239A",
			x"0000" when x"239B",
			x"0000" when x"239C",
			x"0000" when x"239D",
			x"0000" when x"239E",
			x"0000" when x"239F",
			x"0000" when x"23A0",
			x"0000" when x"23A1",
			x"0000" when x"23A2",
			x"0000" when x"23A3",
			x"0000" when x"23A4",
			x"0000" when x"23A5",
			x"0000" when x"23A6",
			x"0000" when x"23A7",
			x"0000" when x"23A8",
			x"0000" when x"23A9",
			x"0000" when x"23AA",
			x"0000" when x"23AB",
			x"0000" when x"23AC",
			x"0000" when x"23AD",
			x"0000" when x"23AE",
			x"0000" when x"23AF",
			x"0000" when x"23B0",
			x"0000" when x"23B1",
			x"0000" when x"23B2",
			x"0000" when x"23B3",
			x"0000" when x"23B4",
			x"0000" when x"23B5",
			x"0000" when x"23B6",
			x"0000" when x"23B7",
			x"0000" when x"23B8",
			x"0000" when x"23B9",
			x"0000" when x"23BA",
			x"0000" when x"23BB",
			x"0000" when x"23BC",
			x"0000" when x"23BD",
			x"0000" when x"23BE",
			x"0000" when x"23BF",
			x"0000" when x"23C0",
			x"0000" when x"23C1",
			x"0000" when x"23C2",
			x"0000" when x"23C3",
			x"0000" when x"23C4",
			x"0000" when x"23C5",
			x"0000" when x"23C6",
			x"0000" when x"23C7",
			x"0000" when x"23C8",
			x"0000" when x"23C9",
			x"0000" when x"23CA",
			x"0000" when x"23CB",
			x"0000" when x"23CC",
			x"0000" when x"23CD",
			x"0000" when x"23CE",
			x"0000" when x"23CF",
			x"0000" when x"23D0",
			x"0000" when x"23D1",
			x"0000" when x"23D2",
			x"0000" when x"23D3",
			x"0000" when x"23D4",
			x"0000" when x"23D5",
			x"0000" when x"23D6",
			x"0000" when x"23D7",
			x"0000" when x"23D8",
			x"0000" when x"23D9",
			x"0000" when x"23DA",
			x"0000" when x"23DB",
			x"0000" when x"23DC",
			x"0000" when x"23DD",
			x"0000" when x"23DE",
			x"0000" when x"23DF",
			x"0000" when x"23E0",
			x"0000" when x"23E1",
			x"0000" when x"23E2",
			x"0000" when x"23E3",
			x"0000" when x"23E4",
			x"0000" when x"23E5",
			x"0000" when x"23E6",
			x"0000" when x"23E7",
			x"0000" when x"23E8",
			x"0000" when x"23E9",
			x"0000" when x"23EA",
			x"0000" when x"23EB",
			x"0000" when x"23EC",
			x"0000" when x"23ED",
			x"0000" when x"23EE",
			x"0000" when x"23EF",
			x"0000" when x"23F0",
			x"0000" when x"23F1",
			x"0000" when x"23F2",
			x"0000" when x"23F3",
			x"0000" when x"23F4",
			x"0000" when x"23F5",
			x"0000" when x"23F6",
			x"0000" when x"23F7",
			x"0000" when x"23F8",
			x"0000" when x"23F9",
			x"0000" when x"23FA",
			x"0000" when x"23FB",
			x"0000" when x"23FC",
			x"0000" when x"23FD",
			x"0000" when x"23FE",
			x"0000" when x"23FF",
			x"0000" when x"2400",
			x"0000" when x"2401",
			x"0000" when x"2402",
			x"0000" when x"2403",
			x"0000" when x"2404",
			x"0000" when x"2405",
			x"0000" when x"2406",
			x"0000" when x"2407",
			x"0000" when x"2408",
			x"0000" when x"2409",
			x"0000" when x"240A",
			x"0000" when x"240B",
			x"0000" when x"240C",
			x"0000" when x"240D",
			x"0000" when x"240E",
			x"0000" when x"240F",
			x"0000" when x"2410",
			x"0000" when x"2411",
			x"0000" when x"2412",
			x"0000" when x"2413",
			x"0000" when x"2414",
			x"0000" when x"2415",
			x"0000" when x"2416",
			x"0000" when x"2417",
			x"0000" when x"2418",
			x"0000" when x"2419",
			x"0000" when x"241A",
			x"0000" when x"241B",
			x"0000" when x"241C",
			x"0000" when x"241D",
			x"0000" when x"241E",
			x"0000" when x"241F",
			x"0000" when x"2420",
			x"0000" when x"2421",
			x"0000" when x"2422",
			x"0000" when x"2423",
			x"0000" when x"2424",
			x"0000" when x"2425",
			x"0000" when x"2426",
			x"0000" when x"2427",
			x"0000" when x"2428",
			x"0000" when x"2429",
			x"0000" when x"242A",
			x"0000" when x"242B",
			x"0000" when x"242C",
			x"0000" when x"242D",
			x"0000" when x"242E",
			x"0000" when x"242F",
			x"0000" when x"2430",
			x"0000" when x"2431",
			x"0000" when x"2432",
			x"0000" when x"2433",
			x"0000" when x"2434",
			x"0000" when x"2435",
			x"0000" when x"2436",
			x"0000" when x"2437",
			x"0000" when x"2438",
			x"0000" when x"2439",
			x"0000" when x"243A",
			x"0000" when x"243B",
			x"0000" when x"243C",
			x"0000" when x"243D",
			x"0000" when x"243E",
			x"0000" when x"243F",
			x"0000" when x"2440",
			x"0000" when x"2441",
			x"0000" when x"2442",
			x"0000" when x"2443",
			x"0000" when x"2444",
			x"0000" when x"2445",
			x"0000" when x"2446",
			x"0000" when x"2447",
			x"0000" when x"2448",
			x"0000" when x"2449",
			x"0000" when x"244A",
			x"0000" when x"244B",
			x"0000" when x"244C",
			x"0000" when x"244D",
			x"0000" when x"244E",
			x"0000" when x"244F",
			x"0000" when x"2450",
			x"0000" when x"2451",
			x"0000" when x"2452",
			x"0000" when x"2453",
			x"0000" when x"2454",
			x"0000" when x"2455",
			x"0000" when x"2456",
			x"0000" when x"2457",
			x"0000" when x"2458",
			x"0000" when x"2459",
			x"0000" when x"245A",
			x"0000" when x"245B",
			x"0000" when x"245C",
			x"0000" when x"245D",
			x"0000" when x"245E",
			x"0000" when x"245F",
			x"0000" when x"2460",
			x"0000" when x"2461",
			x"0000" when x"2462",
			x"0000" when x"2463",
			x"0000" when x"2464",
			x"0000" when x"2465",
			x"0000" when x"2466",
			x"0000" when x"2467",
			x"0000" when x"2468",
			x"0000" when x"2469",
			x"0000" when x"246A",
			x"0000" when x"246B",
			x"0000" when x"246C",
			x"0000" when x"246D",
			x"0000" when x"246E",
			x"0000" when x"246F",
			x"0000" when x"2470",
			x"0000" when x"2471",
			x"0000" when x"2472",
			x"0000" when x"2473",
			x"0000" when x"2474",
			x"0000" when x"2475",
			x"0000" when x"2476",
			x"0000" when x"2477",
			x"0000" when x"2478",
			x"0000" when x"2479",
			x"0000" when x"247A",
			x"0000" when x"247B",
			x"0000" when x"247C",
			x"0000" when x"247D",
			x"0000" when x"247E",
			x"0000" when x"247F",
			x"0000" when x"2480",
			x"0000" when x"2481",
			x"0000" when x"2482",
			x"0000" when x"2483",
			x"0000" when x"2484",
			x"0000" when x"2485",
			x"0000" when x"2486",
			x"0000" when x"2487",
			x"0000" when x"2488",
			x"0000" when x"2489",
			x"0000" when x"248A",
			x"0000" when x"248B",
			x"0000" when x"248C",
			x"0000" when x"248D",
			x"0000" when x"248E",
			x"0000" when x"248F",
			x"0000" when x"2490",
			x"0000" when x"2491",
			x"0000" when x"2492",
			x"0000" when x"2493",
			x"0000" when x"2494",
			x"0000" when x"2495",
			x"0000" when x"2496",
			x"0000" when x"2497",
			x"0000" when x"2498",
			x"0000" when x"2499",
			x"0000" when x"249A",
			x"0000" when x"249B",
			x"0000" when x"249C",
			x"0000" when x"249D",
			x"0000" when x"249E",
			x"0000" when x"249F",
			x"0000" when x"24A0",
			x"0000" when x"24A1",
			x"0000" when x"24A2",
			x"0000" when x"24A3",
			x"0000" when x"24A4",
			x"0000" when x"24A5",
			x"0000" when x"24A6",
			x"0000" when x"24A7",
			x"0000" when x"24A8",
			x"0000" when x"24A9",
			x"0000" when x"24AA",
			x"0000" when x"24AB",
			x"0000" when x"24AC",
			x"0000" when x"24AD",
			x"0000" when x"24AE",
			x"0000" when x"24AF",
			x"0000" when x"24B0",
			x"0000" when x"24B1",
			x"0000" when x"24B2",
			x"0000" when x"24B3",
			x"0000" when x"24B4",
			x"0000" when x"24B5",
			x"0000" when x"24B6",
			x"0000" when x"24B7",
			x"0000" when x"24B8",
			x"0000" when x"24B9",
			x"0000" when x"24BA",
			x"0000" when x"24BB",
			x"0000" when x"24BC",
			x"0000" when x"24BD",
			x"0000" when x"24BE",
			x"0000" when x"24BF",
			x"0000" when x"24C0",
			x"0000" when x"24C1",
			x"0000" when x"24C2",
			x"0000" when x"24C3",
			x"0000" when x"24C4",
			x"0000" when x"24C5",
			x"0000" when x"24C6",
			x"0000" when x"24C7",
			x"0000" when x"24C8",
			x"0000" when x"24C9",
			x"0000" when x"24CA",
			x"0000" when x"24CB",
			x"0000" when x"24CC",
			x"0000" when x"24CD",
			x"0000" when x"24CE",
			x"0000" when x"24CF",
			x"0000" when x"24D0",
			x"0000" when x"24D1",
			x"0000" when x"24D2",
			x"0000" when x"24D3",
			x"0000" when x"24D4",
			x"0000" when x"24D5",
			x"0000" when x"24D6",
			x"0000" when x"24D7",
			x"0000" when x"24D8",
			x"0000" when x"24D9",
			x"0000" when x"24DA",
			x"0000" when x"24DB",
			x"0000" when x"24DC",
			x"0000" when x"24DD",
			x"0000" when x"24DE",
			x"0000" when x"24DF",
			x"0000" when x"24E0",
			x"0000" when x"24E1",
			x"0000" when x"24E2",
			x"0000" when x"24E3",
			x"0000" when x"24E4",
			x"0000" when x"24E5",
			x"0000" when x"24E6",
			x"0000" when x"24E7",
			x"0000" when x"24E8",
			x"0000" when x"24E9",
			x"0000" when x"24EA",
			x"0000" when x"24EB",
			x"0000" when x"24EC",
			x"0000" when x"24ED",
			x"0000" when x"24EE",
			x"0000" when x"24EF",
			x"0000" when x"24F0",
			x"0000" when x"24F1",
			x"0000" when x"24F2",
			x"0000" when x"24F3",
			x"0000" when x"24F4",
			x"0000" when x"24F5",
			x"0000" when x"24F6",
			x"0000" when x"24F7",
			x"0000" when x"24F8",
			x"0000" when x"24F9",
			x"0000" when x"24FA",
			x"0000" when x"24FB",
			x"0000" when x"24FC",
			x"0000" when x"24FD",
			x"0000" when x"24FE",
			x"0000" when x"24FF",
			x"0000" when x"2500",
			x"0000" when x"2501",
			x"0000" when x"2502",
			x"0000" when x"2503",
			x"0000" when x"2504",
			x"0000" when x"2505",
			x"0000" when x"2506",
			x"0000" when x"2507",
			x"0000" when x"2508",
			x"0000" when x"2509",
			x"0000" when x"250A",
			x"0000" when x"250B",
			x"0000" when x"250C",
			x"0000" when x"250D",
			x"0000" when x"250E",
			x"0000" when x"250F",
			x"0000" when x"2510",
			x"0000" when x"2511",
			x"0000" when x"2512",
			x"0000" when x"2513",
			x"0000" when x"2514",
			x"0000" when x"2515",
			x"0000" when x"2516",
			x"0000" when x"2517",
			x"0000" when x"2518",
			x"0000" when x"2519",
			x"0000" when x"251A",
			x"0000" when x"251B",
			x"0000" when x"251C",
			x"0000" when x"251D",
			x"0000" when x"251E",
			x"0000" when x"251F",
			x"0000" when x"2520",
			x"0000" when x"2521",
			x"0000" when x"2522",
			x"0000" when x"2523",
			x"0000" when x"2524",
			x"0000" when x"2525",
			x"0000" when x"2526",
			x"0000" when x"2527",
			x"0000" when x"2528",
			x"0000" when x"2529",
			x"0000" when x"252A",
			x"0000" when x"252B",
			x"0000" when x"252C",
			x"0000" when x"252D",
			x"0000" when x"252E",
			x"0000" when x"252F",
			x"0000" when x"2530",
			x"0000" when x"2531",
			x"0000" when x"2532",
			x"0000" when x"2533",
			x"0000" when x"2534",
			x"0000" when x"2535",
			x"0000" when x"2536",
			x"0000" when x"2537",
			x"0000" when x"2538",
			x"0000" when x"2539",
			x"0000" when x"253A",
			x"0000" when x"253B",
			x"0000" when x"253C",
			x"0000" when x"253D",
			x"0000" when x"253E",
			x"0000" when x"253F",
			x"0000" when x"2540",
			x"0000" when x"2541",
			x"0000" when x"2542",
			x"0000" when x"2543",
			x"0000" when x"2544",
			x"0000" when x"2545",
			x"0000" when x"2546",
			x"0000" when x"2547",
			x"0000" when x"2548",
			x"0000" when x"2549",
			x"0000" when x"254A",
			x"0000" when x"254B",
			x"0000" when x"254C",
			x"0000" when x"254D",
			x"0000" when x"254E",
			x"0000" when x"254F",
			x"0000" when x"2550",
			x"0000" when x"2551",
			x"0000" when x"2552",
			x"0000" when x"2553",
			x"0000" when x"2554",
			x"0000" when x"2555",
			x"0000" when x"2556",
			x"0000" when x"2557",
			x"0000" when x"2558",
			x"0000" when x"2559",
			x"0000" when x"255A",
			x"0000" when x"255B",
			x"0000" when x"255C",
			x"0000" when x"255D",
			x"0000" when x"255E",
			x"0000" when x"255F",
			x"0000" when x"2560",
			x"0000" when x"2561",
			x"0000" when x"2562",
			x"0000" when x"2563",
			x"0000" when x"2564",
			x"0000" when x"2565",
			x"0000" when x"2566",
			x"0000" when x"2567",
			x"0000" when x"2568",
			x"0000" when x"2569",
			x"0000" when x"256A",
			x"0000" when x"256B",
			x"0000" when x"256C",
			x"0000" when x"256D",
			x"0000" when x"256E",
			x"0000" when x"256F",
			x"0000" when x"2570",
			x"0000" when x"2571",
			x"0000" when x"2572",
			x"0000" when x"2573",
			x"0000" when x"2574",
			x"0000" when x"2575",
			x"0000" when x"2576",
			x"0000" when x"2577",
			x"0000" when x"2578",
			x"0000" when x"2579",
			x"0000" when x"257A",
			x"0000" when x"257B",
			x"0000" when x"257C",
			x"0000" when x"257D",
			x"0000" when x"257E",
			x"0000" when x"257F",
			x"0000" when x"2580",
			x"0000" when x"2581",
			x"0000" when x"2582",
			x"0000" when x"2583",
			x"0000" when x"2584",
			x"0000" when x"2585",
			x"0000" when x"2586",
			x"0000" when x"2587",
			x"0000" when x"2588",
			x"0000" when x"2589",
			x"0000" when x"258A",
			x"0000" when x"258B",
			x"0000" when x"258C",
			x"0000" when x"258D",
			x"0000" when x"258E",
			x"0000" when x"258F",
			x"0000" when x"2590",
			x"0000" when x"2591",
			x"0000" when x"2592",
			x"0000" when x"2593",
			x"0000" when x"2594",
			x"0000" when x"2595",
			x"0000" when x"2596",
			x"0000" when x"2597",
			x"0000" when x"2598",
			x"0000" when x"2599",
			x"0000" when x"259A",
			x"0000" when x"259B",
			x"0000" when x"259C",
			x"0000" when x"259D",
			x"0000" when x"259E",
			x"0000" when x"259F",
			x"0000" when x"25A0",
			x"0000" when x"25A1",
			x"0000" when x"25A2",
			x"0000" when x"25A3",
			x"0000" when x"25A4",
			x"0000" when x"25A5",
			x"0000" when x"25A6",
			x"0000" when x"25A7",
			x"0000" when x"25A8",
			x"0000" when x"25A9",
			x"0000" when x"25AA",
			x"0000" when x"25AB",
			x"0000" when x"25AC",
			x"0000" when x"25AD",
			x"0000" when x"25AE",
			x"0000" when x"25AF",
			x"0000" when x"25B0",
			x"0000" when x"25B1",
			x"0000" when x"25B2",
			x"0000" when x"25B3",
			x"0000" when x"25B4",
			x"0000" when x"25B5",
			x"0000" when x"25B6",
			x"0000" when x"25B7",
			x"0000" when x"25B8",
			x"0000" when x"25B9",
			x"0000" when x"25BA",
			x"0000" when x"25BB",
			x"0000" when x"25BC",
			x"0000" when x"25BD",
			x"0000" when x"25BE",
			x"0000" when x"25BF",
			x"0000" when x"25C0",
			x"0000" when x"25C1",
			x"0000" when x"25C2",
			x"0000" when x"25C3",
			x"0000" when x"25C4",
			x"0000" when x"25C5",
			x"0000" when x"25C6",
			x"0000" when x"25C7",
			x"0000" when x"25C8",
			x"0000" when x"25C9",
			x"0000" when x"25CA",
			x"0000" when x"25CB",
			x"0000" when x"25CC",
			x"0000" when x"25CD",
			x"0000" when x"25CE",
			x"0000" when x"25CF",
			x"0000" when x"25D0",
			x"0000" when x"25D1",
			x"0000" when x"25D2",
			x"0000" when x"25D3",
			x"0000" when x"25D4",
			x"0000" when x"25D5",
			x"0000" when x"25D6",
			x"0000" when x"25D7",
			x"0000" when x"25D8",
			x"0000" when x"25D9",
			x"0000" when x"25DA",
			x"0000" when x"25DB",
			x"0000" when x"25DC",
			x"0000" when x"25DD",
			x"0000" when x"25DE",
			x"0000" when x"25DF",
			x"0000" when x"25E0",
			x"0000" when x"25E1",
			x"0000" when x"25E2",
			x"0000" when x"25E3",
			x"0000" when x"25E4",
			x"0000" when x"25E5",
			x"0000" when x"25E6",
			x"0000" when x"25E7",
			x"0000" when x"25E8",
			x"0000" when x"25E9",
			x"0000" when x"25EA",
			x"0000" when x"25EB",
			x"0000" when x"25EC",
			x"0000" when x"25ED",
			x"0000" when x"25EE",
			x"0000" when x"25EF",
			x"0000" when x"25F0",
			x"0000" when x"25F1",
			x"0000" when x"25F2",
			x"0000" when x"25F3",
			x"0000" when x"25F4",
			x"0000" when x"25F5",
			x"0000" when x"25F6",
			x"0000" when x"25F7",
			x"0000" when x"25F8",
			x"0000" when x"25F9",
			x"0000" when x"25FA",
			x"0000" when x"25FB",
			x"0000" when x"25FC",
			x"0000" when x"25FD",
			x"0000" when x"25FE",
			x"0000" when x"25FF",
			x"0000" when x"2600",
			x"0000" when x"2601",
			x"0000" when x"2602",
			x"0000" when x"2603",
			x"0000" when x"2604",
			x"0000" when x"2605",
			x"0000" when x"2606",
			x"0000" when x"2607",
			x"0000" when x"2608",
			x"0000" when x"2609",
			x"0000" when x"260A",
			x"0000" when x"260B",
			x"0000" when x"260C",
			x"0000" when x"260D",
			x"0000" when x"260E",
			x"0000" when x"260F",
			x"0000" when x"2610",
			x"0000" when x"2611",
			x"0000" when x"2612",
			x"0000" when x"2613",
			x"0000" when x"2614",
			x"0000" when x"2615",
			x"0000" when x"2616",
			x"0000" when x"2617",
			x"0000" when x"2618",
			x"0000" when x"2619",
			x"0000" when x"261A",
			x"0000" when x"261B",
			x"0000" when x"261C",
			x"0000" when x"261D",
			x"0000" when x"261E",
			x"0000" when x"261F",
			x"0000" when x"2620",
			x"0000" when x"2621",
			x"0000" when x"2622",
			x"0000" when x"2623",
			x"0000" when x"2624",
			x"0000" when x"2625",
			x"0000" when x"2626",
			x"0000" when x"2627",
			x"0000" when x"2628",
			x"0000" when x"2629",
			x"0000" when x"262A",
			x"0000" when x"262B",
			x"0000" when x"262C",
			x"0000" when x"262D",
			x"0000" when x"262E",
			x"0000" when x"262F",
			x"0000" when x"2630",
			x"0000" when x"2631",
			x"0000" when x"2632",
			x"0000" when x"2633",
			x"0000" when x"2634",
			x"0000" when x"2635",
			x"0000" when x"2636",
			x"0000" when x"2637",
			x"0000" when x"2638",
			x"0000" when x"2639",
			x"0000" when x"263A",
			x"0000" when x"263B",
			x"0000" when x"263C",
			x"0000" when x"263D",
			x"0000" when x"263E",
			x"0000" when x"263F",
			x"0000" when x"2640",
			x"0000" when x"2641",
			x"0000" when x"2642",
			x"0000" when x"2643",
			x"0000" when x"2644",
			x"0000" when x"2645",
			x"0000" when x"2646",
			x"0000" when x"2647",
			x"0000" when x"2648",
			x"0000" when x"2649",
			x"0000" when x"264A",
			x"0000" when x"264B",
			x"0000" when x"264C",
			x"0000" when x"264D",
			x"0000" when x"264E",
			x"0000" when x"264F",
			x"0000" when x"2650",
			x"0000" when x"2651",
			x"0000" when x"2652",
			x"0000" when x"2653",
			x"0000" when x"2654",
			x"0000" when x"2655",
			x"0000" when x"2656",
			x"0000" when x"2657",
			x"0000" when x"2658",
			x"0000" when x"2659",
			x"0000" when x"265A",
			x"0000" when x"265B",
			x"0000" when x"265C",
			x"0000" when x"265D",
			x"0000" when x"265E",
			x"0000" when x"265F",
			x"0000" when x"2660",
			x"0000" when x"2661",
			x"0000" when x"2662",
			x"0000" when x"2663",
			x"0000" when x"2664",
			x"0000" when x"2665",
			x"0000" when x"2666",
			x"0000" when x"2667",
			x"0000" when x"2668",
			x"0000" when x"2669",
			x"0000" when x"266A",
			x"0000" when x"266B",
			x"0000" when x"266C",
			x"0000" when x"266D",
			x"0000" when x"266E",
			x"0000" when x"266F",
			x"0000" when x"2670",
			x"0000" when x"2671",
			x"0000" when x"2672",
			x"0000" when x"2673",
			x"0000" when x"2674",
			x"0000" when x"2675",
			x"0000" when x"2676",
			x"0000" when x"2677",
			x"0000" when x"2678",
			x"0000" when x"2679",
			x"0000" when x"267A",
			x"0000" when x"267B",
			x"0000" when x"267C",
			x"0000" when x"267D",
			x"0000" when x"267E",
			x"0000" when x"267F",
			x"0000" when x"2680",
			x"0000" when x"2681",
			x"0000" when x"2682",
			x"0000" when x"2683",
			x"0000" when x"2684",
			x"0000" when x"2685",
			x"0000" when x"2686",
			x"0000" when x"2687",
			x"0000" when x"2688",
			x"0000" when x"2689",
			x"0000" when x"268A",
			x"0000" when x"268B",
			x"0000" when x"268C",
			x"0000" when x"268D",
			x"0000" when x"268E",
			x"0000" when x"268F",
			x"0000" when x"2690",
			x"0000" when x"2691",
			x"0000" when x"2692",
			x"0000" when x"2693",
			x"0000" when x"2694",
			x"0000" when x"2695",
			x"0000" when x"2696",
			x"0000" when x"2697",
			x"0000" when x"2698",
			x"0000" when x"2699",
			x"0000" when x"269A",
			x"0000" when x"269B",
			x"0000" when x"269C",
			x"0000" when x"269D",
			x"0000" when x"269E",
			x"0000" when x"269F",
			x"0000" when x"26A0",
			x"0000" when x"26A1",
			x"0000" when x"26A2",
			x"0000" when x"26A3",
			x"0000" when x"26A4",
			x"0000" when x"26A5",
			x"0000" when x"26A6",
			x"0000" when x"26A7",
			x"0000" when x"26A8",
			x"0000" when x"26A9",
			x"0000" when x"26AA",
			x"0000" when x"26AB",
			x"0000" when x"26AC",
			x"0000" when x"26AD",
			x"0000" when x"26AE",
			x"0000" when x"26AF",
			x"0000" when x"26B0",
			x"0000" when x"26B1",
			x"0000" when x"26B2",
			x"0000" when x"26B3",
			x"0000" when x"26B4",
			x"0000" when x"26B5",
			x"0000" when x"26B6",
			x"0000" when x"26B7",
			x"0000" when x"26B8",
			x"0000" when x"26B9",
			x"0000" when x"26BA",
			x"0000" when x"26BB",
			x"0000" when x"26BC",
			x"0000" when x"26BD",
			x"0000" when x"26BE",
			x"0000" when x"26BF",
			x"0000" when x"26C0",
			x"0000" when x"26C1",
			x"0000" when x"26C2",
			x"0000" when x"26C3",
			x"0000" when x"26C4",
			x"0000" when x"26C5",
			x"0000" when x"26C6",
			x"0000" when x"26C7",
			x"0000" when x"26C8",
			x"0000" when x"26C9",
			x"0000" when x"26CA",
			x"0000" when x"26CB",
			x"0000" when x"26CC",
			x"0000" when x"26CD",
			x"0000" when x"26CE",
			x"0000" when x"26CF",
			x"0000" when x"26D0",
			x"0000" when x"26D1",
			x"0000" when x"26D2",
			x"0000" when x"26D3",
			x"0000" when x"26D4",
			x"0000" when x"26D5",
			x"0000" when x"26D6",
			x"0000" when x"26D7",
			x"0000" when x"26D8",
			x"0000" when x"26D9",
			x"0000" when x"26DA",
			x"0000" when x"26DB",
			x"0000" when x"26DC",
			x"0000" when x"26DD",
			x"0000" when x"26DE",
			x"0000" when x"26DF",
			x"0000" when x"26E0",
			x"0000" when x"26E1",
			x"0000" when x"26E2",
			x"0000" when x"26E3",
			x"0000" when x"26E4",
			x"0000" when x"26E5",
			x"0000" when x"26E6",
			x"0000" when x"26E7",
			x"0000" when x"26E8",
			x"0000" when x"26E9",
			x"0000" when x"26EA",
			x"0000" when x"26EB",
			x"0000" when x"26EC",
			x"0000" when x"26ED",
			x"0000" when x"26EE",
			x"0000" when x"26EF",
			x"0000" when x"26F0",
			x"0000" when x"26F1",
			x"0000" when x"26F2",
			x"0000" when x"26F3",
			x"0000" when x"26F4",
			x"0000" when x"26F5",
			x"0000" when x"26F6",
			x"0000" when x"26F7",
			x"0000" when x"26F8",
			x"0000" when x"26F9",
			x"0000" when x"26FA",
			x"0000" when x"26FB",
			x"0000" when x"26FC",
			x"0000" when x"26FD",
			x"0000" when x"26FE",
			x"0000" when x"26FF",
			x"0000" when x"2700",
			x"0000" when x"2701",
			x"0000" when x"2702",
			x"0000" when x"2703",
			x"0000" when x"2704",
			x"0000" when x"2705",
			x"0000" when x"2706",
			x"0000" when x"2707",
			x"0000" when x"2708",
			x"0000" when x"2709",
			x"0000" when x"270A",
			x"0000" when x"270B",
			x"0000" when x"270C",
			x"0000" when x"270D",
			x"0000" when x"270E",
			x"0000" when x"270F",
			x"0000" when x"2710",
			x"0000" when x"2711",
			x"0000" when x"2712",
			x"0000" when x"2713",
			x"0000" when x"2714",
			x"0000" when x"2715",
			x"0000" when x"2716",
			x"0000" when x"2717",
			x"0000" when x"2718",
			x"0000" when x"2719",
			x"0000" when x"271A",
			x"0000" when x"271B",
			x"0000" when x"271C",
			x"0000" when x"271D",
			x"0000" when x"271E",
			x"0000" when x"271F",
			x"0000" when x"2720",
			x"0000" when x"2721",
			x"0000" when x"2722",
			x"0000" when x"2723",
			x"0000" when x"2724",
			x"0000" when x"2725",
			x"0000" when x"2726",
			x"0000" when x"2727",
			x"0000" when x"2728",
			x"0000" when x"2729",
			x"0000" when x"272A",
			x"0000" when x"272B",
			x"0000" when x"272C",
			x"0000" when x"272D",
			x"0000" when x"272E",
			x"0000" when x"272F",
			x"0000" when x"2730",
			x"0000" when x"2731",
			x"0000" when x"2732",
			x"0000" when x"2733",
			x"0000" when x"2734",
			x"0000" when x"2735",
			x"0000" when x"2736",
			x"0000" when x"2737",
			x"0000" when x"2738",
			x"0000" when x"2739",
			x"0000" when x"273A",
			x"0000" when x"273B",
			x"0000" when x"273C",
			x"0000" when x"273D",
			x"0000" when x"273E",
			x"0000" when x"273F",
			x"0000" when x"2740",
			x"0000" when x"2741",
			x"0000" when x"2742",
			x"0000" when x"2743",
			x"0000" when x"2744",
			x"0000" when x"2745",
			x"0000" when x"2746",
			x"0000" when x"2747",
			x"0000" when x"2748",
			x"0000" when x"2749",
			x"0000" when x"274A",
			x"0000" when x"274B",
			x"0000" when x"274C",
			x"0000" when x"274D",
			x"0000" when x"274E",
			x"0000" when x"274F",
			x"0000" when x"2750",
			x"0000" when x"2751",
			x"0000" when x"2752",
			x"0000" when x"2753",
			x"0000" when x"2754",
			x"0000" when x"2755",
			x"0000" when x"2756",
			x"0000" when x"2757",
			x"0000" when x"2758",
			x"0000" when x"2759",
			x"0000" when x"275A",
			x"0000" when x"275B",
			x"0000" when x"275C",
			x"0000" when x"275D",
			x"0000" when x"275E",
			x"0000" when x"275F",
			x"0000" when x"2760",
			x"0000" when x"2761",
			x"0000" when x"2762",
			x"0000" when x"2763",
			x"0000" when x"2764",
			x"0000" when x"2765",
			x"0000" when x"2766",
			x"0000" when x"2767",
			x"0000" when x"2768",
			x"0000" when x"2769",
			x"0000" when x"276A",
			x"0000" when x"276B",
			x"0000" when x"276C",
			x"0000" when x"276D",
			x"0000" when x"276E",
			x"0000" when x"276F",
			x"0000" when x"2770",
			x"0000" when x"2771",
			x"0000" when x"2772",
			x"0000" when x"2773",
			x"0000" when x"2774",
			x"0000" when x"2775",
			x"0000" when x"2776",
			x"0000" when x"2777",
			x"0000" when x"2778",
			x"0000" when x"2779",
			x"0000" when x"277A",
			x"0000" when x"277B",
			x"0000" when x"277C",
			x"0000" when x"277D",
			x"0000" when x"277E",
			x"0000" when x"277F",
			x"0000" when x"2780",
			x"0000" when x"2781",
			x"0000" when x"2782",
			x"0000" when x"2783",
			x"0000" when x"2784",
			x"0000" when x"2785",
			x"0000" when x"2786",
			x"0000" when x"2787",
			x"0000" when x"2788",
			x"0000" when x"2789",
			x"0000" when x"278A",
			x"0000" when x"278B",
			x"0000" when x"278C",
			x"0000" when x"278D",
			x"0000" when x"278E",
			x"0000" when x"278F",
			x"0000" when x"2790",
			x"0000" when x"2791",
			x"0000" when x"2792",
			x"0000" when x"2793",
			x"0000" when x"2794",
			x"0000" when x"2795",
			x"0000" when x"2796",
			x"0000" when x"2797",
			x"0000" when x"2798",
			x"0000" when x"2799",
			x"0000" when x"279A",
			x"0000" when x"279B",
			x"0000" when x"279C",
			x"0000" when x"279D",
			x"0000" when x"279E",
			x"0000" when x"279F",
			x"0000" when x"27A0",
			x"0000" when x"27A1",
			x"0000" when x"27A2",
			x"0000" when x"27A3",
			x"0000" when x"27A4",
			x"0000" when x"27A5",
			x"0000" when x"27A6",
			x"0000" when x"27A7",
			x"0000" when x"27A8",
			x"0000" when x"27A9",
			x"0000" when x"27AA",
			x"0000" when x"27AB",
			x"0000" when x"27AC",
			x"0000" when x"27AD",
			x"0000" when x"27AE",
			x"0000" when x"27AF",
			x"0000" when x"27B0",
			x"0000" when x"27B1",
			x"0000" when x"27B2",
			x"0000" when x"27B3",
			x"0000" when x"27B4",
			x"0000" when x"27B5",
			x"0000" when x"27B6",
			x"0000" when x"27B7",
			x"0000" when x"27B8",
			x"0000" when x"27B9",
			x"0000" when x"27BA",
			x"0000" when x"27BB",
			x"0000" when x"27BC",
			x"0000" when x"27BD",
			x"0000" when x"27BE",
			x"0000" when x"27BF",
			x"0000" when x"27C0",
			x"0000" when x"27C1",
			x"0000" when x"27C2",
			x"0000" when x"27C3",
			x"0000" when x"27C4",
			x"0000" when x"27C5",
			x"0000" when x"27C6",
			x"0000" when x"27C7",
			x"0000" when x"27C8",
			x"0000" when x"27C9",
			x"0000" when x"27CA",
			x"0000" when x"27CB",
			x"0000" when x"27CC",
			x"0000" when x"27CD",
			x"0000" when x"27CE",
			x"0000" when x"27CF",
			x"0000" when x"27D0",
			x"0000" when x"27D1",
			x"0000" when x"27D2",
			x"0000" when x"27D3",
			x"0000" when x"27D4",
			x"0000" when x"27D5",
			x"0000" when x"27D6",
			x"0000" when x"27D7",
			x"0000" when x"27D8",
			x"0000" when x"27D9",
			x"0000" when x"27DA",
			x"0000" when x"27DB",
			x"0000" when x"27DC",
			x"0000" when x"27DD",
			x"0000" when x"27DE",
			x"0000" when x"27DF",
			x"0000" when x"27E0",
			x"0000" when x"27E1",
			x"0000" when x"27E2",
			x"0000" when x"27E3",
			x"0000" when x"27E4",
			x"0000" when x"27E5",
			x"0000" when x"27E6",
			x"0000" when x"27E7",
			x"0000" when x"27E8",
			x"0000" when x"27E9",
			x"0000" when x"27EA",
			x"0000" when x"27EB",
			x"0000" when x"27EC",
			x"0000" when x"27ED",
			x"0000" when x"27EE",
			x"0000" when x"27EF",
			x"0000" when x"27F0",
			x"0000" when x"27F1",
			x"0000" when x"27F2",
			x"0000" when x"27F3",
			x"0000" when x"27F4",
			x"0000" when x"27F5",
			x"0000" when x"27F6",
			x"0000" when x"27F7",
			x"0000" when x"27F8",
			x"0000" when x"27F9",
			x"0000" when x"27FA",
			x"0000" when x"27FB",
			x"0000" when x"27FC",
			x"0000" when x"27FD",
			x"0000" when x"27FE",
			x"0000" when x"27FF",
			x"0000" when x"2800",
			x"0000" when x"2801",
			x"0000" when x"2802",
			x"0000" when x"2803",
			x"0000" when x"2804",
			x"0000" when x"2805",
			x"0000" when x"2806",
			x"0000" when x"2807",
			x"0000" when x"2808",
			x"0000" when x"2809",
			x"0000" when x"280A",
			x"0000" when x"280B",
			x"0000" when x"280C",
			x"0000" when x"280D",
			x"0000" when x"280E",
			x"0000" when x"280F",
			x"0000" when x"2810",
			x"0000" when x"2811",
			x"0000" when x"2812",
			x"0000" when x"2813",
			x"0000" when x"2814",
			x"0000" when x"2815",
			x"0000" when x"2816",
			x"0000" when x"2817",
			x"0000" when x"2818",
			x"0000" when x"2819",
			x"0000" when x"281A",
			x"0000" when x"281B",
			x"0000" when x"281C",
			x"0000" when x"281D",
			x"0000" when x"281E",
			x"0000" when x"281F",
			x"0000" when x"2820",
			x"0000" when x"2821",
			x"0000" when x"2822",
			x"0000" when x"2823",
			x"0000" when x"2824",
			x"0000" when x"2825",
			x"0000" when x"2826",
			x"0000" when x"2827",
			x"0000" when x"2828",
			x"0000" when x"2829",
			x"0000" when x"282A",
			x"0000" when x"282B",
			x"0000" when x"282C",
			x"0000" when x"282D",
			x"0000" when x"282E",
			x"0000" when x"282F",
			x"0000" when x"2830",
			x"0000" when x"2831",
			x"0000" when x"2832",
			x"0000" when x"2833",
			x"0000" when x"2834",
			x"0000" when x"2835",
			x"0000" when x"2836",
			x"0000" when x"2837",
			x"0000" when x"2838",
			x"0000" when x"2839",
			x"0000" when x"283A",
			x"0000" when x"283B",
			x"0000" when x"283C",
			x"0000" when x"283D",
			x"0000" when x"283E",
			x"0000" when x"283F",
			x"0000" when x"2840",
			x"0000" when x"2841",
			x"0000" when x"2842",
			x"0000" when x"2843",
			x"0000" when x"2844",
			x"0000" when x"2845",
			x"0000" when x"2846",
			x"0000" when x"2847",
			x"0000" when x"2848",
			x"0000" when x"2849",
			x"0000" when x"284A",
			x"0000" when x"284B",
			x"0000" when x"284C",
			x"0000" when x"284D",
			x"0000" when x"284E",
			x"0000" when x"284F",
			x"0000" when x"2850",
			x"0000" when x"2851",
			x"0000" when x"2852",
			x"0000" when x"2853",
			x"0000" when x"2854",
			x"0000" when x"2855",
			x"0000" when x"2856",
			x"0000" when x"2857",
			x"0000" when x"2858",
			x"0000" when x"2859",
			x"0000" when x"285A",
			x"0000" when x"285B",
			x"0000" when x"285C",
			x"0000" when x"285D",
			x"0000" when x"285E",
			x"0000" when x"285F",
			x"0000" when x"2860",
			x"0000" when x"2861",
			x"0000" when x"2862",
			x"0000" when x"2863",
			x"0000" when x"2864",
			x"0000" when x"2865",
			x"0000" when x"2866",
			x"0000" when x"2867",
			x"0000" when x"2868",
			x"0000" when x"2869",
			x"0000" when x"286A",
			x"0000" when x"286B",
			x"0000" when x"286C",
			x"0000" when x"286D",
			x"0000" when x"286E",
			x"0000" when x"286F",
			x"0000" when x"2870",
			x"0000" when x"2871",
			x"0000" when x"2872",
			x"0000" when x"2873",
			x"0000" when x"2874",
			x"0000" when x"2875",
			x"0000" when x"2876",
			x"0000" when x"2877",
			x"0000" when x"2878",
			x"0000" when x"2879",
			x"0000" when x"287A",
			x"0000" when x"287B",
			x"0000" when x"287C",
			x"0000" when x"287D",
			x"0000" when x"287E",
			x"0000" when x"287F",
			x"0000" when x"2880",
			x"0000" when x"2881",
			x"0000" when x"2882",
			x"0000" when x"2883",
			x"0000" when x"2884",
			x"0000" when x"2885",
			x"0000" when x"2886",
			x"0000" when x"2887",
			x"0000" when x"2888",
			x"0000" when x"2889",
			x"0000" when x"288A",
			x"0000" when x"288B",
			x"0000" when x"288C",
			x"0000" when x"288D",
			x"0000" when x"288E",
			x"0000" when x"288F",
			x"0000" when x"2890",
			x"0000" when x"2891",
			x"0000" when x"2892",
			x"0000" when x"2893",
			x"0000" when x"2894",
			x"0000" when x"2895",
			x"0000" when x"2896",
			x"0000" when x"2897",
			x"0000" when x"2898",
			x"0000" when x"2899",
			x"0000" when x"289A",
			x"0000" when x"289B",
			x"0000" when x"289C",
			x"0000" when x"289D",
			x"0000" when x"289E",
			x"0000" when x"289F",
			x"0000" when x"28A0",
			x"0000" when x"28A1",
			x"0000" when x"28A2",
			x"0000" when x"28A3",
			x"0000" when x"28A4",
			x"0000" when x"28A5",
			x"0000" when x"28A6",
			x"0000" when x"28A7",
			x"0000" when x"28A8",
			x"0000" when x"28A9",
			x"0000" when x"28AA",
			x"0000" when x"28AB",
			x"0000" when x"28AC",
			x"0000" when x"28AD",
			x"0000" when x"28AE",
			x"0000" when x"28AF",
			x"0000" when x"28B0",
			x"0000" when x"28B1",
			x"0000" when x"28B2",
			x"0000" when x"28B3",
			x"0000" when x"28B4",
			x"0000" when x"28B5",
			x"0000" when x"28B6",
			x"0000" when x"28B7",
			x"0000" when x"28B8",
			x"0000" when x"28B9",
			x"0000" when x"28BA",
			x"0000" when x"28BB",
			x"0000" when x"28BC",
			x"0000" when x"28BD",
			x"0000" when x"28BE",
			x"0000" when x"28BF",
			x"0000" when x"28C0",
			x"0000" when x"28C1",
			x"0000" when x"28C2",
			x"0000" when x"28C3",
			x"0000" when x"28C4",
			x"0000" when x"28C5",
			x"0000" when x"28C6",
			x"0000" when x"28C7",
			x"0000" when x"28C8",
			x"0000" when x"28C9",
			x"0000" when x"28CA",
			x"0000" when x"28CB",
			x"0000" when x"28CC",
			x"0000" when x"28CD",
			x"0000" when x"28CE",
			x"0000" when x"28CF",
			x"0000" when x"28D0",
			x"0000" when x"28D1",
			x"0000" when x"28D2",
			x"0000" when x"28D3",
			x"0000" when x"28D4",
			x"0000" when x"28D5",
			x"0000" when x"28D6",
			x"0000" when x"28D7",
			x"0000" when x"28D8",
			x"0000" when x"28D9",
			x"0000" when x"28DA",
			x"0000" when x"28DB",
			x"0000" when x"28DC",
			x"0000" when x"28DD",
			x"0000" when x"28DE",
			x"0000" when x"28DF",
			x"0000" when x"28E0",
			x"0000" when x"28E1",
			x"0000" when x"28E2",
			x"0000" when x"28E3",
			x"0000" when x"28E4",
			x"0000" when x"28E5",
			x"0000" when x"28E6",
			x"0000" when x"28E7",
			x"0000" when x"28E8",
			x"0000" when x"28E9",
			x"0000" when x"28EA",
			x"0000" when x"28EB",
			x"0000" when x"28EC",
			x"0000" when x"28ED",
			x"0000" when x"28EE",
			x"0000" when x"28EF",
			x"0000" when x"28F0",
			x"0000" when x"28F1",
			x"0000" when x"28F2",
			x"0000" when x"28F3",
			x"0000" when x"28F4",
			x"0000" when x"28F5",
			x"0000" when x"28F6",
			x"0000" when x"28F7",
			x"0000" when x"28F8",
			x"0000" when x"28F9",
			x"0000" when x"28FA",
			x"0000" when x"28FB",
			x"0000" when x"28FC",
			x"0000" when x"28FD",
			x"0000" when x"28FE",
			x"0000" when x"28FF",
			x"0000" when x"2900",
			x"0000" when x"2901",
			x"0000" when x"2902",
			x"0000" when x"2903",
			x"0000" when x"2904",
			x"0000" when x"2905",
			x"0000" when x"2906",
			x"0000" when x"2907",
			x"0000" when x"2908",
			x"0000" when x"2909",
			x"0000" when x"290A",
			x"0000" when x"290B",
			x"0000" when x"290C",
			x"0000" when x"290D",
			x"0000" when x"290E",
			x"0000" when x"290F",
			x"0000" when x"2910",
			x"0000" when x"2911",
			x"0000" when x"2912",
			x"0000" when x"2913",
			x"0000" when x"2914",
			x"0000" when x"2915",
			x"0000" when x"2916",
			x"0000" when x"2917",
			x"0000" when x"2918",
			x"0000" when x"2919",
			x"0000" when x"291A",
			x"0000" when x"291B",
			x"0000" when x"291C",
			x"0000" when x"291D",
			x"0000" when x"291E",
			x"0000" when x"291F",
			x"0000" when x"2920",
			x"0000" when x"2921",
			x"0000" when x"2922",
			x"0000" when x"2923",
			x"0000" when x"2924",
			x"0000" when x"2925",
			x"0000" when x"2926",
			x"0000" when x"2927",
			x"0000" when x"2928",
			x"0000" when x"2929",
			x"0000" when x"292A",
			x"0000" when x"292B",
			x"0000" when x"292C",
			x"0000" when x"292D",
			x"0000" when x"292E",
			x"0000" when x"292F",
			x"0000" when x"2930",
			x"0000" when x"2931",
			x"0000" when x"2932",
			x"0000" when x"2933",
			x"0000" when x"2934",
			x"0000" when x"2935",
			x"0000" when x"2936",
			x"0000" when x"2937",
			x"0000" when x"2938",
			x"0000" when x"2939",
			x"0000" when x"293A",
			x"0000" when x"293B",
			x"0000" when x"293C",
			x"0000" when x"293D",
			x"0000" when x"293E",
			x"0000" when x"293F",
			x"0000" when x"2940",
			x"0000" when x"2941",
			x"0000" when x"2942",
			x"0000" when x"2943",
			x"0000" when x"2944",
			x"0000" when x"2945",
			x"0000" when x"2946",
			x"0000" when x"2947",
			x"0000" when x"2948",
			x"0000" when x"2949",
			x"0000" when x"294A",
			x"0000" when x"294B",
			x"0000" when x"294C",
			x"0000" when x"294D",
			x"0000" when x"294E",
			x"0000" when x"294F",
			x"0000" when x"2950",
			x"0000" when x"2951",
			x"0000" when x"2952",
			x"0000" when x"2953",
			x"0000" when x"2954",
			x"0000" when x"2955",
			x"0000" when x"2956",
			x"0000" when x"2957",
			x"0000" when x"2958",
			x"0000" when x"2959",
			x"0000" when x"295A",
			x"0000" when x"295B",
			x"0000" when x"295C",
			x"0000" when x"295D",
			x"0000" when x"295E",
			x"0000" when x"295F",
			x"0000" when x"2960",
			x"0000" when x"2961",
			x"0000" when x"2962",
			x"0000" when x"2963",
			x"0000" when x"2964",
			x"0000" when x"2965",
			x"0000" when x"2966",
			x"0000" when x"2967",
			x"0000" when x"2968",
			x"0000" when x"2969",
			x"0000" when x"296A",
			x"0000" when x"296B",
			x"0000" when x"296C",
			x"0000" when x"296D",
			x"0000" when x"296E",
			x"0000" when x"296F",
			x"0000" when x"2970",
			x"0000" when x"2971",
			x"0000" when x"2972",
			x"0000" when x"2973",
			x"0000" when x"2974",
			x"0000" when x"2975",
			x"0000" when x"2976",
			x"0000" when x"2977",
			x"0000" when x"2978",
			x"0000" when x"2979",
			x"0000" when x"297A",
			x"0000" when x"297B",
			x"0000" when x"297C",
			x"0000" when x"297D",
			x"0000" when x"297E",
			x"0000" when x"297F",
			x"0000" when x"2980",
			x"0000" when x"2981",
			x"0000" when x"2982",
			x"0000" when x"2983",
			x"0000" when x"2984",
			x"0000" when x"2985",
			x"0000" when x"2986",
			x"0000" when x"2987",
			x"0000" when x"2988",
			x"0000" when x"2989",
			x"0000" when x"298A",
			x"0000" when x"298B",
			x"0000" when x"298C",
			x"0000" when x"298D",
			x"0000" when x"298E",
			x"0000" when x"298F",
			x"0000" when x"2990",
			x"0000" when x"2991",
			x"0000" when x"2992",
			x"0000" when x"2993",
			x"0000" when x"2994",
			x"0000" when x"2995",
			x"0000" when x"2996",
			x"0000" when x"2997",
			x"0000" when x"2998",
			x"0000" when x"2999",
			x"0000" when x"299A",
			x"0000" when x"299B",
			x"0000" when x"299C",
			x"0000" when x"299D",
			x"0000" when x"299E",
			x"0000" when x"299F",
			x"0000" when x"29A0",
			x"0000" when x"29A1",
			x"0000" when x"29A2",
			x"0000" when x"29A3",
			x"0000" when x"29A4",
			x"0000" when x"29A5",
			x"0000" when x"29A6",
			x"0000" when x"29A7",
			x"0000" when x"29A8",
			x"0000" when x"29A9",
			x"0000" when x"29AA",
			x"0000" when x"29AB",
			x"0000" when x"29AC",
			x"0000" when x"29AD",
			x"0000" when x"29AE",
			x"0000" when x"29AF",
			x"0000" when x"29B0",
			x"0000" when x"29B1",
			x"0000" when x"29B2",
			x"0000" when x"29B3",
			x"0000" when x"29B4",
			x"0000" when x"29B5",
			x"0000" when x"29B6",
			x"0000" when x"29B7",
			x"0000" when x"29B8",
			x"0000" when x"29B9",
			x"0000" when x"29BA",
			x"0000" when x"29BB",
			x"0000" when x"29BC",
			x"0000" when x"29BD",
			x"0000" when x"29BE",
			x"0000" when x"29BF",
			x"0000" when x"29C0",
			x"0000" when x"29C1",
			x"0000" when x"29C2",
			x"0000" when x"29C3",
			x"0000" when x"29C4",
			x"0000" when x"29C5",
			x"0000" when x"29C6",
			x"0000" when x"29C7",
			x"0000" when x"29C8",
			x"0000" when x"29C9",
			x"0000" when x"29CA",
			x"0000" when x"29CB",
			x"0000" when x"29CC",
			x"0000" when x"29CD",
			x"0000" when x"29CE",
			x"0000" when x"29CF",
			x"0000" when x"29D0",
			x"0000" when x"29D1",
			x"0000" when x"29D2",
			x"0000" when x"29D3",
			x"0000" when x"29D4",
			x"0000" when x"29D5",
			x"0000" when x"29D6",
			x"0000" when x"29D7",
			x"0000" when x"29D8",
			x"0000" when x"29D9",
			x"0000" when x"29DA",
			x"0000" when x"29DB",
			x"0000" when x"29DC",
			x"0000" when x"29DD",
			x"0000" when x"29DE",
			x"0000" when x"29DF",
			x"0000" when x"29E0",
			x"0000" when x"29E1",
			x"0000" when x"29E2",
			x"0000" when x"29E3",
			x"0000" when x"29E4",
			x"0000" when x"29E5",
			x"0000" when x"29E6",
			x"0000" when x"29E7",
			x"0000" when x"29E8",
			x"0000" when x"29E9",
			x"0000" when x"29EA",
			x"0000" when x"29EB",
			x"0000" when x"29EC",
			x"0000" when x"29ED",
			x"0000" when x"29EE",
			x"0000" when x"29EF",
			x"0000" when x"29F0",
			x"0000" when x"29F1",
			x"0000" when x"29F2",
			x"0000" when x"29F3",
			x"0000" when x"29F4",
			x"0000" when x"29F5",
			x"0000" when x"29F6",
			x"0000" when x"29F7",
			x"0000" when x"29F8",
			x"0000" when x"29F9",
			x"0000" when x"29FA",
			x"0000" when x"29FB",
			x"0000" when x"29FC",
			x"0000" when x"29FD",
			x"0000" when x"29FE",
			x"0000" when x"29FF",
			x"0000" when x"2A00",
			x"0000" when x"2A01",
			x"0000" when x"2A02",
			x"0000" when x"2A03",
			x"0000" when x"2A04",
			x"0000" when x"2A05",
			x"0000" when x"2A06",
			x"0000" when x"2A07",
			x"0000" when x"2A08",
			x"0000" when x"2A09",
			x"0000" when x"2A0A",
			x"0000" when x"2A0B",
			x"0000" when x"2A0C",
			x"0000" when x"2A0D",
			x"0000" when x"2A0E",
			x"0000" when x"2A0F",
			x"0000" when x"2A10",
			x"0000" when x"2A11",
			x"0000" when x"2A12",
			x"0000" when x"2A13",
			x"0000" when x"2A14",
			x"0000" when x"2A15",
			x"0000" when x"2A16",
			x"0000" when x"2A17",
			x"0000" when x"2A18",
			x"0000" when x"2A19",
			x"0000" when x"2A1A",
			x"0000" when x"2A1B",
			x"0000" when x"2A1C",
			x"0000" when x"2A1D",
			x"0000" when x"2A1E",
			x"0000" when x"2A1F",
			x"0000" when x"2A20",
			x"0000" when x"2A21",
			x"0000" when x"2A22",
			x"0000" when x"2A23",
			x"0000" when x"2A24",
			x"0000" when x"2A25",
			x"0000" when x"2A26",
			x"0000" when x"2A27",
			x"0000" when x"2A28",
			x"0000" when x"2A29",
			x"0000" when x"2A2A",
			x"0000" when x"2A2B",
			x"0000" when x"2A2C",
			x"0000" when x"2A2D",
			x"0000" when x"2A2E",
			x"0000" when x"2A2F",
			x"0000" when x"2A30",
			x"0000" when x"2A31",
			x"0000" when x"2A32",
			x"0000" when x"2A33",
			x"0000" when x"2A34",
			x"0000" when x"2A35",
			x"0000" when x"2A36",
			x"0000" when x"2A37",
			x"0000" when x"2A38",
			x"0000" when x"2A39",
			x"0000" when x"2A3A",
			x"0000" when x"2A3B",
			x"0000" when x"2A3C",
			x"0000" when x"2A3D",
			x"0000" when x"2A3E",
			x"0000" when x"2A3F",
			x"0000" when x"2A40",
			x"0000" when x"2A41",
			x"0000" when x"2A42",
			x"0000" when x"2A43",
			x"0000" when x"2A44",
			x"0000" when x"2A45",
			x"0000" when x"2A46",
			x"0000" when x"2A47",
			x"0000" when x"2A48",
			x"0000" when x"2A49",
			x"0000" when x"2A4A",
			x"0000" when x"2A4B",
			x"0000" when x"2A4C",
			x"0000" when x"2A4D",
			x"0000" when x"2A4E",
			x"0000" when x"2A4F",
			x"0000" when x"2A50",
			x"0000" when x"2A51",
			x"0000" when x"2A52",
			x"0000" when x"2A53",
			x"0000" when x"2A54",
			x"0000" when x"2A55",
			x"0000" when x"2A56",
			x"0000" when x"2A57",
			x"0000" when x"2A58",
			x"0000" when x"2A59",
			x"0000" when x"2A5A",
			x"0000" when x"2A5B",
			x"0000" when x"2A5C",
			x"0000" when x"2A5D",
			x"0000" when x"2A5E",
			x"0000" when x"2A5F",
			x"0000" when x"2A60",
			x"0000" when x"2A61",
			x"0000" when x"2A62",
			x"0000" when x"2A63",
			x"0000" when x"2A64",
			x"0000" when x"2A65",
			x"0000" when x"2A66",
			x"0000" when x"2A67",
			x"0000" when x"2A68",
			x"0000" when x"2A69",
			x"0000" when x"2A6A",
			x"0000" when x"2A6B",
			x"0000" when x"2A6C",
			x"0000" when x"2A6D",
			x"0000" when x"2A6E",
			x"0000" when x"2A6F",
			x"0000" when x"2A70",
			x"0000" when x"2A71",
			x"0000" when x"2A72",
			x"0000" when x"2A73",
			x"0000" when x"2A74",
			x"0000" when x"2A75",
			x"0000" when x"2A76",
			x"0000" when x"2A77",
			x"0000" when x"2A78",
			x"0000" when x"2A79",
			x"0000" when x"2A7A",
			x"0000" when x"2A7B",
			x"0000" when x"2A7C",
			x"0000" when x"2A7D",
			x"0000" when x"2A7E",
			x"0000" when x"2A7F",
			x"0000" when x"2A80",
			x"0000" when x"2A81",
			x"0000" when x"2A82",
			x"0000" when x"2A83",
			x"0000" when x"2A84",
			x"0000" when x"2A85",
			x"0000" when x"2A86",
			x"0000" when x"2A87",
			x"0000" when x"2A88",
			x"0000" when x"2A89",
			x"0000" when x"2A8A",
			x"0000" when x"2A8B",
			x"0000" when x"2A8C",
			x"0000" when x"2A8D",
			x"0000" when x"2A8E",
			x"0000" when x"2A8F",
			x"0000" when x"2A90",
			x"0000" when x"2A91",
			x"0000" when x"2A92",
			x"0000" when x"2A93",
			x"0000" when x"2A94",
			x"0000" when x"2A95",
			x"0000" when x"2A96",
			x"0000" when x"2A97",
			x"0000" when x"2A98",
			x"0000" when x"2A99",
			x"0000" when x"2A9A",
			x"0000" when x"2A9B",
			x"0000" when x"2A9C",
			x"0000" when x"2A9D",
			x"0000" when x"2A9E",
			x"0000" when x"2A9F",
			x"0000" when x"2AA0",
			x"0000" when x"2AA1",
			x"0000" when x"2AA2",
			x"0000" when x"2AA3",
			x"0000" when x"2AA4",
			x"0000" when x"2AA5",
			x"0000" when x"2AA6",
			x"0000" when x"2AA7",
			x"0000" when x"2AA8",
			x"0000" when x"2AA9",
			x"0000" when x"2AAA",
			x"0000" when x"2AAB",
			x"0000" when x"2AAC",
			x"0000" when x"2AAD",
			x"0000" when x"2AAE",
			x"0000" when x"2AAF",
			x"0000" when x"2AB0",
			x"0000" when x"2AB1",
			x"0000" when x"2AB2",
			x"0000" when x"2AB3",
			x"0000" when x"2AB4",
			x"0000" when x"2AB5",
			x"0000" when x"2AB6",
			x"0000" when x"2AB7",
			x"0000" when x"2AB8",
			x"0000" when x"2AB9",
			x"0000" when x"2ABA",
			x"0000" when x"2ABB",
			x"0000" when x"2ABC",
			x"0000" when x"2ABD",
			x"0000" when x"2ABE",
			x"0000" when x"2ABF",
			x"0000" when x"2AC0",
			x"0000" when x"2AC1",
			x"0000" when x"2AC2",
			x"0000" when x"2AC3",
			x"0000" when x"2AC4",
			x"0000" when x"2AC5",
			x"0000" when x"2AC6",
			x"0000" when x"2AC7",
			x"0000" when x"2AC8",
			x"0000" when x"2AC9",
			x"0000" when x"2ACA",
			x"0000" when x"2ACB",
			x"0000" when x"2ACC",
			x"0000" when x"2ACD",
			x"0000" when x"2ACE",
			x"0000" when x"2ACF",
			x"0000" when x"2AD0",
			x"0000" when x"2AD1",
			x"0000" when x"2AD2",
			x"0000" when x"2AD3",
			x"0000" when x"2AD4",
			x"0000" when x"2AD5",
			x"0000" when x"2AD6",
			x"0000" when x"2AD7",
			x"0000" when x"2AD8",
			x"0000" when x"2AD9",
			x"0000" when x"2ADA",
			x"0000" when x"2ADB",
			x"0000" when x"2ADC",
			x"0000" when x"2ADD",
			x"0000" when x"2ADE",
			x"0000" when x"2ADF",
			x"0000" when x"2AE0",
			x"0000" when x"2AE1",
			x"0000" when x"2AE2",
			x"0000" when x"2AE3",
			x"0000" when x"2AE4",
			x"0000" when x"2AE5",
			x"0000" when x"2AE6",
			x"0000" when x"2AE7",
			x"0000" when x"2AE8",
			x"0000" when x"2AE9",
			x"0000" when x"2AEA",
			x"0000" when x"2AEB",
			x"0000" when x"2AEC",
			x"0000" when x"2AED",
			x"0000" when x"2AEE",
			x"0000" when x"2AEF",
			x"0000" when x"2AF0",
			x"0000" when x"2AF1",
			x"0000" when x"2AF2",
			x"0000" when x"2AF3",
			x"0000" when x"2AF4",
			x"0000" when x"2AF5",
			x"0000" when x"2AF6",
			x"0000" when x"2AF7",
			x"0000" when x"2AF8",
			x"0000" when x"2AF9",
			x"0000" when x"2AFA",
			x"0000" when x"2AFB",
			x"0000" when x"2AFC",
			x"0000" when x"2AFD",
			x"0000" when x"2AFE",
			x"0000" when x"2AFF",
			x"0000" when x"2B00",
			x"0000" when x"2B01",
			x"0000" when x"2B02",
			x"0000" when x"2B03",
			x"0000" when x"2B04",
			x"0000" when x"2B05",
			x"0000" when x"2B06",
			x"0000" when x"2B07",
			x"0000" when x"2B08",
			x"0000" when x"2B09",
			x"0000" when x"2B0A",
			x"0000" when x"2B0B",
			x"0000" when x"2B0C",
			x"0000" when x"2B0D",
			x"0000" when x"2B0E",
			x"0000" when x"2B0F",
			x"0000" when x"2B10",
			x"0000" when x"2B11",
			x"0000" when x"2B12",
			x"0000" when x"2B13",
			x"0000" when x"2B14",
			x"0000" when x"2B15",
			x"0000" when x"2B16",
			x"0000" when x"2B17",
			x"0000" when x"2B18",
			x"0000" when x"2B19",
			x"0000" when x"2B1A",
			x"0000" when x"2B1B",
			x"0000" when x"2B1C",
			x"0000" when x"2B1D",
			x"0000" when x"2B1E",
			x"0000" when x"2B1F",
			x"0000" when x"2B20",
			x"0000" when x"2B21",
			x"0000" when x"2B22",
			x"0000" when x"2B23",
			x"0000" when x"2B24",
			x"0000" when x"2B25",
			x"0000" when x"2B26",
			x"0000" when x"2B27",
			x"0000" when x"2B28",
			x"0000" when x"2B29",
			x"0000" when x"2B2A",
			x"0000" when x"2B2B",
			x"0000" when x"2B2C",
			x"0000" when x"2B2D",
			x"0000" when x"2B2E",
			x"0000" when x"2B2F",
			x"0000" when x"2B30",
			x"0000" when x"2B31",
			x"0000" when x"2B32",
			x"0000" when x"2B33",
			x"0000" when x"2B34",
			x"0000" when x"2B35",
			x"0000" when x"2B36",
			x"0000" when x"2B37",
			x"0000" when x"2B38",
			x"0000" when x"2B39",
			x"0000" when x"2B3A",
			x"0000" when x"2B3B",
			x"0000" when x"2B3C",
			x"0000" when x"2B3D",
			x"0000" when x"2B3E",
			x"0000" when x"2B3F",
			x"0000" when x"2B40",
			x"0000" when x"2B41",
			x"0000" when x"2B42",
			x"0000" when x"2B43",
			x"0000" when x"2B44",
			x"0000" when x"2B45",
			x"0000" when x"2B46",
			x"0000" when x"2B47",
			x"0000" when x"2B48",
			x"0000" when x"2B49",
			x"0000" when x"2B4A",
			x"0000" when x"2B4B",
			x"0000" when x"2B4C",
			x"0000" when x"2B4D",
			x"0000" when x"2B4E",
			x"0000" when x"2B4F",
			x"0000" when x"2B50",
			x"0000" when x"2B51",
			x"0000" when x"2B52",
			x"0000" when x"2B53",
			x"0000" when x"2B54",
			x"0000" when x"2B55",
			x"0000" when x"2B56",
			x"0000" when x"2B57",
			x"0000" when x"2B58",
			x"0000" when x"2B59",
			x"0000" when x"2B5A",
			x"0000" when x"2B5B",
			x"0000" when x"2B5C",
			x"0000" when x"2B5D",
			x"0000" when x"2B5E",
			x"0000" when x"2B5F",
			x"0000" when x"2B60",
			x"0000" when x"2B61",
			x"0000" when x"2B62",
			x"0000" when x"2B63",
			x"0000" when x"2B64",
			x"0000" when x"2B65",
			x"0000" when x"2B66",
			x"0000" when x"2B67",
			x"0000" when x"2B68",
			x"0000" when x"2B69",
			x"0000" when x"2B6A",
			x"0000" when x"2B6B",
			x"0000" when x"2B6C",
			x"0000" when x"2B6D",
			x"0000" when x"2B6E",
			x"0000" when x"2B6F",
			x"0000" when x"2B70",
			x"0000" when x"2B71",
			x"0000" when x"2B72",
			x"0000" when x"2B73",
			x"0000" when x"2B74",
			x"0000" when x"2B75",
			x"0000" when x"2B76",
			x"0000" when x"2B77",
			x"0000" when x"2B78",
			x"0000" when x"2B79",
			x"0000" when x"2B7A",
			x"0000" when x"2B7B",
			x"0000" when x"2B7C",
			x"0000" when x"2B7D",
			x"0000" when x"2B7E",
			x"0000" when x"2B7F",
			x"0000" when x"2B80",
			x"0000" when x"2B81",
			x"0000" when x"2B82",
			x"0000" when x"2B83",
			x"0000" when x"2B84",
			x"0000" when x"2B85",
			x"0000" when x"2B86",
			x"0000" when x"2B87",
			x"0000" when x"2B88",
			x"0000" when x"2B89",
			x"0000" when x"2B8A",
			x"0000" when x"2B8B",
			x"0000" when x"2B8C",
			x"0000" when x"2B8D",
			x"0000" when x"2B8E",
			x"0000" when x"2B8F",
			x"0000" when x"2B90",
			x"0000" when x"2B91",
			x"0000" when x"2B92",
			x"0000" when x"2B93",
			x"0000" when x"2B94",
			x"0000" when x"2B95",
			x"0000" when x"2B96",
			x"0000" when x"2B97",
			x"0000" when x"2B98",
			x"0000" when x"2B99",
			x"0000" when x"2B9A",
			x"0000" when x"2B9B",
			x"0000" when x"2B9C",
			x"0000" when x"2B9D",
			x"0000" when x"2B9E",
			x"0000" when x"2B9F",
			x"0000" when x"2BA0",
			x"0000" when x"2BA1",
			x"0000" when x"2BA2",
			x"0000" when x"2BA3",
			x"0000" when x"2BA4",
			x"0000" when x"2BA5",
			x"0000" when x"2BA6",
			x"0000" when x"2BA7",
			x"0000" when x"2BA8",
			x"0000" when x"2BA9",
			x"0000" when x"2BAA",
			x"0000" when x"2BAB",
			x"0000" when x"2BAC",
			x"0000" when x"2BAD",
			x"0000" when x"2BAE",
			x"0000" when x"2BAF",
			x"0000" when x"2BB0",
			x"0000" when x"2BB1",
			x"0000" when x"2BB2",
			x"0000" when x"2BB3",
			x"0000" when x"2BB4",
			x"0000" when x"2BB5",
			x"0000" when x"2BB6",
			x"0000" when x"2BB7",
			x"0000" when x"2BB8",
			x"0000" when x"2BB9",
			x"0000" when x"2BBA",
			x"0000" when x"2BBB",
			x"0000" when x"2BBC",
			x"0000" when x"2BBD",
			x"0000" when x"2BBE",
			x"0000" when x"2BBF",
			x"0000" when x"2BC0",
			x"0000" when x"2BC1",
			x"0000" when x"2BC2",
			x"0000" when x"2BC3",
			x"0000" when x"2BC4",
			x"0000" when x"2BC5",
			x"0000" when x"2BC6",
			x"0000" when x"2BC7",
			x"0000" when x"2BC8",
			x"0000" when x"2BC9",
			x"0000" when x"2BCA",
			x"0000" when x"2BCB",
			x"0000" when x"2BCC",
			x"0000" when x"2BCD",
			x"0000" when x"2BCE",
			x"0000" when x"2BCF",
			x"0000" when x"2BD0",
			x"0000" when x"2BD1",
			x"0000" when x"2BD2",
			x"0000" when x"2BD3",
			x"0000" when x"2BD4",
			x"0000" when x"2BD5",
			x"0000" when x"2BD6",
			x"0000" when x"2BD7",
			x"0000" when x"2BD8",
			x"0000" when x"2BD9",
			x"0000" when x"2BDA",
			x"0000" when x"2BDB",
			x"0000" when x"2BDC",
			x"0000" when x"2BDD",
			x"0000" when x"2BDE",
			x"0000" when x"2BDF",
			x"0000" when x"2BE0",
			x"0000" when x"2BE1",
			x"0000" when x"2BE2",
			x"0000" when x"2BE3",
			x"0000" when x"2BE4",
			x"0000" when x"2BE5",
			x"0000" when x"2BE6",
			x"0000" when x"2BE7",
			x"0000" when x"2BE8",
			x"0000" when x"2BE9",
			x"0000" when x"2BEA",
			x"0000" when x"2BEB",
			x"0000" when x"2BEC",
			x"0000" when x"2BED",
			x"0000" when x"2BEE",
			x"0000" when x"2BEF",
			x"0000" when x"2BF0",
			x"0000" when x"2BF1",
			x"0000" when x"2BF2",
			x"0000" when x"2BF3",
			x"0000" when x"2BF4",
			x"0000" when x"2BF5",
			x"0000" when x"2BF6",
			x"0000" when x"2BF7",
			x"0000" when x"2BF8",
			x"0000" when x"2BF9",
			x"0000" when x"2BFA",
			x"0000" when x"2BFB",
			x"0000" when x"2BFC",
			x"0000" when x"2BFD",
			x"0000" when x"2BFE",
			x"0000" when x"2BFF",
			x"0000" when x"2C00",
			x"0000" when x"2C01",
			x"0000" when x"2C02",
			x"0000" when x"2C03",
			x"0000" when x"2C04",
			x"0000" when x"2C05",
			x"0000" when x"2C06",
			x"0000" when x"2C07",
			x"0000" when x"2C08",
			x"0000" when x"2C09",
			x"0000" when x"2C0A",
			x"0000" when x"2C0B",
			x"0000" when x"2C0C",
			x"0000" when x"2C0D",
			x"0000" when x"2C0E",
			x"0000" when x"2C0F",
			x"0000" when x"2C10",
			x"0000" when x"2C11",
			x"0000" when x"2C12",
			x"0000" when x"2C13",
			x"0000" when x"2C14",
			x"0000" when x"2C15",
			x"0000" when x"2C16",
			x"0000" when x"2C17",
			x"0000" when x"2C18",
			x"0000" when x"2C19",
			x"0000" when x"2C1A",
			x"0000" when x"2C1B",
			x"0000" when x"2C1C",
			x"0000" when x"2C1D",
			x"0000" when x"2C1E",
			x"0000" when x"2C1F",
			x"0000" when x"2C20",
			x"0000" when x"2C21",
			x"0000" when x"2C22",
			x"0000" when x"2C23",
			x"0000" when x"2C24",
			x"0000" when x"2C25",
			x"0000" when x"2C26",
			x"0000" when x"2C27",
			x"0000" when x"2C28",
			x"0000" when x"2C29",
			x"0000" when x"2C2A",
			x"0000" when x"2C2B",
			x"0000" when x"2C2C",
			x"0000" when x"2C2D",
			x"0000" when x"2C2E",
			x"0000" when x"2C2F",
			x"0000" when x"2C30",
			x"0000" when x"2C31",
			x"0000" when x"2C32",
			x"0000" when x"2C33",
			x"0000" when x"2C34",
			x"0000" when x"2C35",
			x"0000" when x"2C36",
			x"0000" when x"2C37",
			x"0000" when x"2C38",
			x"0000" when x"2C39",
			x"0000" when x"2C3A",
			x"0000" when x"2C3B",
			x"0000" when x"2C3C",
			x"0000" when x"2C3D",
			x"0000" when x"2C3E",
			x"0000" when x"2C3F",
			x"0000" when x"2C40",
			x"0000" when x"2C41",
			x"0000" when x"2C42",
			x"0000" when x"2C43",
			x"0000" when x"2C44",
			x"0000" when x"2C45",
			x"0000" when x"2C46",
			x"0000" when x"2C47",
			x"0000" when x"2C48",
			x"0000" when x"2C49",
			x"0000" when x"2C4A",
			x"0000" when x"2C4B",
			x"0000" when x"2C4C",
			x"0000" when x"2C4D",
			x"0000" when x"2C4E",
			x"0000" when x"2C4F",
			x"0000" when x"2C50",
			x"0000" when x"2C51",
			x"0000" when x"2C52",
			x"0000" when x"2C53",
			x"0000" when x"2C54",
			x"0000" when x"2C55",
			x"0000" when x"2C56",
			x"0000" when x"2C57",
			x"0000" when x"2C58",
			x"0000" when x"2C59",
			x"0000" when x"2C5A",
			x"0000" when x"2C5B",
			x"0000" when x"2C5C",
			x"0000" when x"2C5D",
			x"0000" when x"2C5E",
			x"0000" when x"2C5F",
			x"0000" when x"2C60",
			x"0000" when x"2C61",
			x"0000" when x"2C62",
			x"0000" when x"2C63",
			x"0000" when x"2C64",
			x"0000" when x"2C65",
			x"0000" when x"2C66",
			x"0000" when x"2C67",
			x"0000" when x"2C68",
			x"0000" when x"2C69",
			x"0000" when x"2C6A",
			x"0000" when x"2C6B",
			x"0000" when x"2C6C",
			x"0000" when x"2C6D",
			x"0000" when x"2C6E",
			x"0000" when x"2C6F",
			x"0000" when x"2C70",
			x"0000" when x"2C71",
			x"0000" when x"2C72",
			x"0000" when x"2C73",
			x"0000" when x"2C74",
			x"0000" when x"2C75",
			x"0000" when x"2C76",
			x"0000" when x"2C77",
			x"0000" when x"2C78",
			x"0000" when x"2C79",
			x"0000" when x"2C7A",
			x"0000" when x"2C7B",
			x"0000" when x"2C7C",
			x"0000" when x"2C7D",
			x"0000" when x"2C7E",
			x"0000" when x"2C7F",
			x"0000" when x"2C80",
			x"0000" when x"2C81",
			x"0000" when x"2C82",
			x"0000" when x"2C83",
			x"0000" when x"2C84",
			x"0000" when x"2C85",
			x"0000" when x"2C86",
			x"0000" when x"2C87",
			x"0000" when x"2C88",
			x"0000" when x"2C89",
			x"0000" when x"2C8A",
			x"0000" when x"2C8B",
			x"0000" when x"2C8C",
			x"0000" when x"2C8D",
			x"0000" when x"2C8E",
			x"0000" when x"2C8F",
			x"0000" when x"2C90",
			x"0000" when x"2C91",
			x"0000" when x"2C92",
			x"0000" when x"2C93",
			x"0000" when x"2C94",
			x"0000" when x"2C95",
			x"0000" when x"2C96",
			x"0000" when x"2C97",
			x"0000" when x"2C98",
			x"0000" when x"2C99",
			x"0000" when x"2C9A",
			x"0000" when x"2C9B",
			x"0000" when x"2C9C",
			x"0000" when x"2C9D",
			x"0000" when x"2C9E",
			x"0000" when x"2C9F",
			x"0000" when x"2CA0",
			x"0000" when x"2CA1",
			x"0000" when x"2CA2",
			x"0000" when x"2CA3",
			x"0000" when x"2CA4",
			x"0000" when x"2CA5",
			x"0000" when x"2CA6",
			x"0000" when x"2CA7",
			x"0000" when x"2CA8",
			x"0000" when x"2CA9",
			x"0000" when x"2CAA",
			x"0000" when x"2CAB",
			x"0000" when x"2CAC",
			x"0000" when x"2CAD",
			x"0000" when x"2CAE",
			x"0000" when x"2CAF",
			x"0000" when x"2CB0",
			x"0000" when x"2CB1",
			x"0000" when x"2CB2",
			x"0000" when x"2CB3",
			x"0000" when x"2CB4",
			x"0000" when x"2CB5",
			x"0000" when x"2CB6",
			x"0000" when x"2CB7",
			x"0000" when x"2CB8",
			x"0000" when x"2CB9",
			x"0000" when x"2CBA",
			x"0000" when x"2CBB",
			x"0000" when x"2CBC",
			x"0000" when x"2CBD",
			x"0000" when x"2CBE",
			x"0000" when x"2CBF",
			x"0000" when x"2CC0",
			x"0000" when x"2CC1",
			x"0000" when x"2CC2",
			x"0000" when x"2CC3",
			x"0000" when x"2CC4",
			x"0000" when x"2CC5",
			x"0000" when x"2CC6",
			x"0000" when x"2CC7",
			x"0000" when x"2CC8",
			x"0000" when x"2CC9",
			x"0000" when x"2CCA",
			x"0000" when x"2CCB",
			x"0000" when x"2CCC",
			x"0000" when x"2CCD",
			x"0000" when x"2CCE",
			x"0000" when x"2CCF",
			x"0000" when x"2CD0",
			x"0000" when x"2CD1",
			x"0000" when x"2CD2",
			x"0000" when x"2CD3",
			x"0000" when x"2CD4",
			x"0000" when x"2CD5",
			x"0000" when x"2CD6",
			x"0000" when x"2CD7",
			x"0000" when x"2CD8",
			x"0000" when x"2CD9",
			x"0000" when x"2CDA",
			x"0000" when x"2CDB",
			x"0000" when x"2CDC",
			x"0000" when x"2CDD",
			x"0000" when x"2CDE",
			x"0000" when x"2CDF",
			x"0000" when x"2CE0",
			x"0000" when x"2CE1",
			x"0000" when x"2CE2",
			x"0000" when x"2CE3",
			x"0000" when x"2CE4",
			x"0000" when x"2CE5",
			x"0000" when x"2CE6",
			x"0000" when x"2CE7",
			x"0000" when x"2CE8",
			x"0000" when x"2CE9",
			x"0000" when x"2CEA",
			x"0000" when x"2CEB",
			x"0000" when x"2CEC",
			x"0000" when x"2CED",
			x"0000" when x"2CEE",
			x"0000" when x"2CEF",
			x"0000" when x"2CF0",
			x"0000" when x"2CF1",
			x"0000" when x"2CF2",
			x"0000" when x"2CF3",
			x"0000" when x"2CF4",
			x"0000" when x"2CF5",
			x"0000" when x"2CF6",
			x"0000" when x"2CF7",
			x"0000" when x"2CF8",
			x"0000" when x"2CF9",
			x"0000" when x"2CFA",
			x"0000" when x"2CFB",
			x"0000" when x"2CFC",
			x"0000" when x"2CFD",
			x"0000" when x"2CFE",
			x"0000" when x"2CFF",
			x"0000" when x"2D00",
			x"0000" when x"2D01",
			x"0000" when x"2D02",
			x"0000" when x"2D03",
			x"0000" when x"2D04",
			x"0000" when x"2D05",
			x"0000" when x"2D06",
			x"0000" when x"2D07",
			x"0000" when x"2D08",
			x"0000" when x"2D09",
			x"0000" when x"2D0A",
			x"0000" when x"2D0B",
			x"0000" when x"2D0C",
			x"0000" when x"2D0D",
			x"0000" when x"2D0E",
			x"0000" when x"2D0F",
			x"0000" when x"2D10",
			x"0000" when x"2D11",
			x"0000" when x"2D12",
			x"0000" when x"2D13",
			x"0000" when x"2D14",
			x"0000" when x"2D15",
			x"0000" when x"2D16",
			x"0000" when x"2D17",
			x"0000" when x"2D18",
			x"0000" when x"2D19",
			x"0000" when x"2D1A",
			x"0000" when x"2D1B",
			x"0000" when x"2D1C",
			x"0000" when x"2D1D",
			x"0000" when x"2D1E",
			x"0000" when x"2D1F",
			x"0000" when x"2D20",
			x"0000" when x"2D21",
			x"0000" when x"2D22",
			x"0000" when x"2D23",
			x"0000" when x"2D24",
			x"0000" when x"2D25",
			x"0000" when x"2D26",
			x"0000" when x"2D27",
			x"0000" when x"2D28",
			x"0000" when x"2D29",
			x"0000" when x"2D2A",
			x"0000" when x"2D2B",
			x"0000" when x"2D2C",
			x"0000" when x"2D2D",
			x"0000" when x"2D2E",
			x"0000" when x"2D2F",
			x"0000" when x"2D30",
			x"0000" when x"2D31",
			x"0000" when x"2D32",
			x"0000" when x"2D33",
			x"0000" when x"2D34",
			x"0000" when x"2D35",
			x"0000" when x"2D36",
			x"0000" when x"2D37",
			x"0000" when x"2D38",
			x"0000" when x"2D39",
			x"0000" when x"2D3A",
			x"0000" when x"2D3B",
			x"0000" when x"2D3C",
			x"0000" when x"2D3D",
			x"0000" when x"2D3E",
			x"0000" when x"2D3F",
			x"0000" when x"2D40",
			x"0000" when x"2D41",
			x"0000" when x"2D42",
			x"0000" when x"2D43",
			x"0000" when x"2D44",
			x"0000" when x"2D45",
			x"0000" when x"2D46",
			x"0000" when x"2D47",
			x"0000" when x"2D48",
			x"0000" when x"2D49",
			x"0000" when x"2D4A",
			x"0000" when x"2D4B",
			x"0000" when x"2D4C",
			x"0000" when x"2D4D",
			x"0000" when x"2D4E",
			x"0000" when x"2D4F",
			x"0000" when x"2D50",
			x"0000" when x"2D51",
			x"0000" when x"2D52",
			x"0000" when x"2D53",
			x"0000" when x"2D54",
			x"0000" when x"2D55",
			x"0000" when x"2D56",
			x"0000" when x"2D57",
			x"0000" when x"2D58",
			x"0000" when x"2D59",
			x"0000" when x"2D5A",
			x"0000" when x"2D5B",
			x"0000" when x"2D5C",
			x"0000" when x"2D5D",
			x"0000" when x"2D5E",
			x"0000" when x"2D5F",
			x"0000" when x"2D60",
			x"0000" when x"2D61",
			x"0000" when x"2D62",
			x"0000" when x"2D63",
			x"0000" when x"2D64",
			x"0000" when x"2D65",
			x"0000" when x"2D66",
			x"0000" when x"2D67",
			x"0000" when x"2D68",
			x"0000" when x"2D69",
			x"0000" when x"2D6A",
			x"0000" when x"2D6B",
			x"0000" when x"2D6C",
			x"0000" when x"2D6D",
			x"0000" when x"2D6E",
			x"0000" when x"2D6F",
			x"0000" when x"2D70",
			x"0000" when x"2D71",
			x"0000" when x"2D72",
			x"0000" when x"2D73",
			x"0000" when x"2D74",
			x"0000" when x"2D75",
			x"0000" when x"2D76",
			x"0000" when x"2D77",
			x"0000" when x"2D78",
			x"0000" when x"2D79",
			x"0000" when x"2D7A",
			x"0000" when x"2D7B",
			x"0000" when x"2D7C",
			x"0000" when x"2D7D",
			x"0000" when x"2D7E",
			x"0000" when x"2D7F",
			x"0000" when x"2D80",
			x"0000" when x"2D81",
			x"0000" when x"2D82",
			x"0000" when x"2D83",
			x"0000" when x"2D84",
			x"0000" when x"2D85",
			x"0000" when x"2D86",
			x"0000" when x"2D87",
			x"0000" when x"2D88",
			x"0000" when x"2D89",
			x"0000" when x"2D8A",
			x"0000" when x"2D8B",
			x"0000" when x"2D8C",
			x"0000" when x"2D8D",
			x"0000" when x"2D8E",
			x"0000" when x"2D8F",
			x"0000" when x"2D90",
			x"0000" when x"2D91",
			x"0000" when x"2D92",
			x"0000" when x"2D93",
			x"0000" when x"2D94",
			x"0000" when x"2D95",
			x"0000" when x"2D96",
			x"0000" when x"2D97",
			x"0000" when x"2D98",
			x"0000" when x"2D99",
			x"0000" when x"2D9A",
			x"0000" when x"2D9B",
			x"0000" when x"2D9C",
			x"0000" when x"2D9D",
			x"0000" when x"2D9E",
			x"0000" when x"2D9F",
			x"0000" when x"2DA0",
			x"0000" when x"2DA1",
			x"0000" when x"2DA2",
			x"0000" when x"2DA3",
			x"0000" when x"2DA4",
			x"0000" when x"2DA5",
			x"0000" when x"2DA6",
			x"0000" when x"2DA7",
			x"0000" when x"2DA8",
			x"0000" when x"2DA9",
			x"0000" when x"2DAA",
			x"0000" when x"2DAB",
			x"0000" when x"2DAC",
			x"0000" when x"2DAD",
			x"0000" when x"2DAE",
			x"0000" when x"2DAF",
			x"0000" when x"2DB0",
			x"0000" when x"2DB1",
			x"0000" when x"2DB2",
			x"0000" when x"2DB3",
			x"0000" when x"2DB4",
			x"0000" when x"2DB5",
			x"0000" when x"2DB6",
			x"0000" when x"2DB7",
			x"0000" when x"2DB8",
			x"0000" when x"2DB9",
			x"0000" when x"2DBA",
			x"0000" when x"2DBB",
			x"0000" when x"2DBC",
			x"0000" when x"2DBD",
			x"0000" when x"2DBE",
			x"0000" when x"2DBF",
			x"0000" when x"2DC0",
			x"0000" when x"2DC1",
			x"0000" when x"2DC2",
			x"0000" when x"2DC3",
			x"0000" when x"2DC4",
			x"0000" when x"2DC5",
			x"0000" when x"2DC6",
			x"0000" when x"2DC7",
			x"0000" when x"2DC8",
			x"0000" when x"2DC9",
			x"0000" when x"2DCA",
			x"0000" when x"2DCB",
			x"0000" when x"2DCC",
			x"0000" when x"2DCD",
			x"0000" when x"2DCE",
			x"0000" when x"2DCF",
			x"0000" when x"2DD0",
			x"0000" when x"2DD1",
			x"0000" when x"2DD2",
			x"0000" when x"2DD3",
			x"0000" when x"2DD4",
			x"0000" when x"2DD5",
			x"0000" when x"2DD6",
			x"0000" when x"2DD7",
			x"0000" when x"2DD8",
			x"0000" when x"2DD9",
			x"0000" when x"2DDA",
			x"0000" when x"2DDB",
			x"0000" when x"2DDC",
			x"0000" when x"2DDD",
			x"0000" when x"2DDE",
			x"0000" when x"2DDF",
			x"0000" when x"2DE0",
			x"0000" when x"2DE1",
			x"0000" when x"2DE2",
			x"0000" when x"2DE3",
			x"0000" when x"2DE4",
			x"0000" when x"2DE5",
			x"0000" when x"2DE6",
			x"0000" when x"2DE7",
			x"0000" when x"2DE8",
			x"0000" when x"2DE9",
			x"0000" when x"2DEA",
			x"0000" when x"2DEB",
			x"0000" when x"2DEC",
			x"0000" when x"2DED",
			x"0000" when x"2DEE",
			x"0000" when x"2DEF",
			x"0000" when x"2DF0",
			x"0000" when x"2DF1",
			x"0000" when x"2DF2",
			x"0000" when x"2DF3",
			x"0000" when x"2DF4",
			x"0000" when x"2DF5",
			x"0000" when x"2DF6",
			x"0000" when x"2DF7",
			x"0000" when x"2DF8",
			x"0000" when x"2DF9",
			x"0000" when x"2DFA",
			x"0000" when x"2DFB",
			x"0000" when x"2DFC",
			x"0000" when x"2DFD",
			x"0000" when x"2DFE",
			x"0000" when x"2DFF",
			x"0000" when x"2E00",
			x"0000" when x"2E01",
			x"0000" when x"2E02",
			x"0000" when x"2E03",
			x"0000" when x"2E04",
			x"0000" when x"2E05",
			x"0000" when x"2E06",
			x"0000" when x"2E07",
			x"0000" when x"2E08",
			x"0000" when x"2E09",
			x"0000" when x"2E0A",
			x"0000" when x"2E0B",
			x"0000" when x"2E0C",
			x"0000" when x"2E0D",
			x"0000" when x"2E0E",
			x"0000" when x"2E0F",
			x"0000" when x"2E10",
			x"0000" when x"2E11",
			x"0000" when x"2E12",
			x"0000" when x"2E13",
			x"0000" when x"2E14",
			x"0000" when x"2E15",
			x"0000" when x"2E16",
			x"0000" when x"2E17",
			x"0000" when x"2E18",
			x"0000" when x"2E19",
			x"0000" when x"2E1A",
			x"0000" when x"2E1B",
			x"0000" when x"2E1C",
			x"0000" when x"2E1D",
			x"0000" when x"2E1E",
			x"0000" when x"2E1F",
			x"0000" when x"2E20",
			x"0000" when x"2E21",
			x"0000" when x"2E22",
			x"0000" when x"2E23",
			x"0000" when x"2E24",
			x"0000" when x"2E25",
			x"0000" when x"2E26",
			x"0000" when x"2E27",
			x"0000" when x"2E28",
			x"0000" when x"2E29",
			x"0000" when x"2E2A",
			x"0000" when x"2E2B",
			x"0000" when x"2E2C",
			x"0000" when x"2E2D",
			x"0000" when x"2E2E",
			x"0000" when x"2E2F",
			x"0000" when x"2E30",
			x"0000" when x"2E31",
			x"0000" when x"2E32",
			x"0000" when x"2E33",
			x"0000" when x"2E34",
			x"0000" when x"2E35",
			x"0000" when x"2E36",
			x"0000" when x"2E37",
			x"0000" when x"2E38",
			x"0000" when x"2E39",
			x"0000" when x"2E3A",
			x"0000" when x"2E3B",
			x"0000" when x"2E3C",
			x"0000" when x"2E3D",
			x"0000" when x"2E3E",
			x"0000" when x"2E3F",
			x"0000" when x"2E40",
			x"0000" when x"2E41",
			x"0000" when x"2E42",
			x"0000" when x"2E43",
			x"0000" when x"2E44",
			x"0000" when x"2E45",
			x"0000" when x"2E46",
			x"0000" when x"2E47",
			x"0000" when x"2E48",
			x"0000" when x"2E49",
			x"0000" when x"2E4A",
			x"0000" when x"2E4B",
			x"0000" when x"2E4C",
			x"0000" when x"2E4D",
			x"0000" when x"2E4E",
			x"0000" when x"2E4F",
			x"0000" when x"2E50",
			x"0000" when x"2E51",
			x"0000" when x"2E52",
			x"0000" when x"2E53",
			x"0000" when x"2E54",
			x"0000" when x"2E55",
			x"0000" when x"2E56",
			x"0000" when x"2E57",
			x"0000" when x"2E58",
			x"0000" when x"2E59",
			x"0000" when x"2E5A",
			x"0000" when x"2E5B",
			x"0000" when x"2E5C",
			x"0000" when x"2E5D",
			x"0000" when x"2E5E",
			x"0000" when x"2E5F",
			x"0000" when x"2E60",
			x"0000" when x"2E61",
			x"0000" when x"2E62",
			x"0000" when x"2E63",
			x"0000" when x"2E64",
			x"0000" when x"2E65",
			x"0000" when x"2E66",
			x"0000" when x"2E67",
			x"0000" when x"2E68",
			x"0000" when x"2E69",
			x"0000" when x"2E6A",
			x"0000" when x"2E6B",
			x"0000" when x"2E6C",
			x"0000" when x"2E6D",
			x"0000" when x"2E6E",
			x"0000" when x"2E6F",
			x"0000" when x"2E70",
			x"0000" when x"2E71",
			x"0000" when x"2E72",
			x"0000" when x"2E73",
			x"0000" when x"2E74",
			x"0000" when x"2E75",
			x"0000" when x"2E76",
			x"0000" when x"2E77",
			x"0000" when x"2E78",
			x"0000" when x"2E79",
			x"0000" when x"2E7A",
			x"0000" when x"2E7B",
			x"0000" when x"2E7C",
			x"0000" when x"2E7D",
			x"0000" when x"2E7E",
			x"0000" when x"2E7F",
			x"0000" when x"2E80",
			x"0000" when x"2E81",
			x"0000" when x"2E82",
			x"0000" when x"2E83",
			x"0000" when x"2E84",
			x"0000" when x"2E85",
			x"0000" when x"2E86",
			x"0000" when x"2E87",
			x"0000" when x"2E88",
			x"0000" when x"2E89",
			x"0000" when x"2E8A",
			x"0000" when x"2E8B",
			x"0000" when x"2E8C",
			x"0000" when x"2E8D",
			x"0000" when x"2E8E",
			x"0000" when x"2E8F",
			x"0000" when x"2E90",
			x"0000" when x"2E91",
			x"0000" when x"2E92",
			x"0000" when x"2E93",
			x"0000" when x"2E94",
			x"0000" when x"2E95",
			x"0000" when x"2E96",
			x"0000" when x"2E97",
			x"0000" when x"2E98",
			x"0000" when x"2E99",
			x"0000" when x"2E9A",
			x"0000" when x"2E9B",
			x"0000" when x"2E9C",
			x"0000" when x"2E9D",
			x"0000" when x"2E9E",
			x"0000" when x"2E9F",
			x"0000" when x"2EA0",
			x"0000" when x"2EA1",
			x"0000" when x"2EA2",
			x"0000" when x"2EA3",
			x"0000" when x"2EA4",
			x"0000" when x"2EA5",
			x"0000" when x"2EA6",
			x"0000" when x"2EA7",
			x"0000" when x"2EA8",
			x"0000" when x"2EA9",
			x"0000" when x"2EAA",
			x"0000" when x"2EAB",
			x"0000" when x"2EAC",
			x"0000" when x"2EAD",
			x"0000" when x"2EAE",
			x"0000" when x"2EAF",
			x"0000" when x"2EB0",
			x"0000" when x"2EB1",
			x"0000" when x"2EB2",
			x"0000" when x"2EB3",
			x"0000" when x"2EB4",
			x"0000" when x"2EB5",
			x"0000" when x"2EB6",
			x"0000" when x"2EB7",
			x"0000" when x"2EB8",
			x"0000" when x"2EB9",
			x"0000" when x"2EBA",
			x"0000" when x"2EBB",
			x"0000" when x"2EBC",
			x"0000" when x"2EBD",
			x"0000" when x"2EBE",
			x"0000" when x"2EBF",
			x"0000" when x"2EC0",
			x"0000" when x"2EC1",
			x"0000" when x"2EC2",
			x"0000" when x"2EC3",
			x"0000" when x"2EC4",
			x"0000" when x"2EC5",
			x"0000" when x"2EC6",
			x"0000" when x"2EC7",
			x"0000" when x"2EC8",
			x"0000" when x"2EC9",
			x"0000" when x"2ECA",
			x"0000" when x"2ECB",
			x"0000" when x"2ECC",
			x"0000" when x"2ECD",
			x"0000" when x"2ECE",
			x"0000" when x"2ECF",
			x"0000" when x"2ED0",
			x"0000" when x"2ED1",
			x"0000" when x"2ED2",
			x"0000" when x"2ED3",
			x"0000" when x"2ED4",
			x"0000" when x"2ED5",
			x"0000" when x"2ED6",
			x"0000" when x"2ED7",
			x"0000" when x"2ED8",
			x"0000" when x"2ED9",
			x"0000" when x"2EDA",
			x"0000" when x"2EDB",
			x"0000" when x"2EDC",
			x"0000" when x"2EDD",
			x"0000" when x"2EDE",
			x"0000" when x"2EDF",
			x"0000" when x"2EE0",
			x"0000" when x"2EE1",
			x"0000" when x"2EE2",
			x"0000" when x"2EE3",
			x"0000" when x"2EE4",
			x"0000" when x"2EE5",
			x"0000" when x"2EE6",
			x"0000" when x"2EE7",
			x"0000" when x"2EE8",
			x"0000" when x"2EE9",
			x"0000" when x"2EEA",
			x"0000" when x"2EEB",
			x"0000" when x"2EEC",
			x"0000" when x"2EED",
			x"0000" when x"2EEE",
			x"0000" when x"2EEF",
			x"0000" when x"2EF0",
			x"0000" when x"2EF1",
			x"0000" when x"2EF2",
			x"0000" when x"2EF3",
			x"0000" when x"2EF4",
			x"0000" when x"2EF5",
			x"0000" when x"2EF6",
			x"0000" when x"2EF7",
			x"0000" when x"2EF8",
			x"0000" when x"2EF9",
			x"0000" when x"2EFA",
			x"0000" when x"2EFB",
			x"0000" when x"2EFC",
			x"0000" when x"2EFD",
			x"0000" when x"2EFE",
			x"0000" when x"2EFF",
			x"0000" when x"2F00",
			x"0000" when x"2F01",
			x"0000" when x"2F02",
			x"0000" when x"2F03",
			x"0000" when x"2F04",
			x"0000" when x"2F05",
			x"0000" when x"2F06",
			x"0000" when x"2F07",
			x"0000" when x"2F08",
			x"0000" when x"2F09",
			x"0000" when x"2F0A",
			x"0000" when x"2F0B",
			x"0000" when x"2F0C",
			x"0000" when x"2F0D",
			x"0000" when x"2F0E",
			x"0000" when x"2F0F",
			x"0000" when x"2F10",
			x"0000" when x"2F11",
			x"0000" when x"2F12",
			x"0000" when x"2F13",
			x"0000" when x"2F14",
			x"0000" when x"2F15",
			x"0000" when x"2F16",
			x"0000" when x"2F17",
			x"0000" when x"2F18",
			x"0000" when x"2F19",
			x"0000" when x"2F1A",
			x"0000" when x"2F1B",
			x"0000" when x"2F1C",
			x"0000" when x"2F1D",
			x"0000" when x"2F1E",
			x"0000" when x"2F1F",
			x"0000" when x"2F20",
			x"0000" when x"2F21",
			x"0000" when x"2F22",
			x"0000" when x"2F23",
			x"0000" when x"2F24",
			x"0000" when x"2F25",
			x"0000" when x"2F26",
			x"0000" when x"2F27",
			x"0000" when x"2F28",
			x"0000" when x"2F29",
			x"0000" when x"2F2A",
			x"0000" when x"2F2B",
			x"0000" when x"2F2C",
			x"0000" when x"2F2D",
			x"0000" when x"2F2E",
			x"0000" when x"2F2F",
			x"0000" when x"2F30",
			x"0000" when x"2F31",
			x"0000" when x"2F32",
			x"0000" when x"2F33",
			x"0000" when x"2F34",
			x"0000" when x"2F35",
			x"0000" when x"2F36",
			x"0000" when x"2F37",
			x"0000" when x"2F38",
			x"0000" when x"2F39",
			x"0000" when x"2F3A",
			x"0000" when x"2F3B",
			x"0000" when x"2F3C",
			x"0000" when x"2F3D",
			x"0000" when x"2F3E",
			x"0000" when x"2F3F",
			x"0000" when x"2F40",
			x"0000" when x"2F41",
			x"0000" when x"2F42",
			x"0000" when x"2F43",
			x"0000" when x"2F44",
			x"0000" when x"2F45",
			x"0000" when x"2F46",
			x"0000" when x"2F47",
			x"0000" when x"2F48",
			x"0000" when x"2F49",
			x"0000" when x"2F4A",
			x"0000" when x"2F4B",
			x"0000" when x"2F4C",
			x"0000" when x"2F4D",
			x"0000" when x"2F4E",
			x"0000" when x"2F4F",
			x"0000" when x"2F50",
			x"0000" when x"2F51",
			x"0000" when x"2F52",
			x"0000" when x"2F53",
			x"0000" when x"2F54",
			x"0000" when x"2F55",
			x"0000" when x"2F56",
			x"0000" when x"2F57",
			x"0000" when x"2F58",
			x"0000" when x"2F59",
			x"0000" when x"2F5A",
			x"0000" when x"2F5B",
			x"0000" when x"2F5C",
			x"0000" when x"2F5D",
			x"0000" when x"2F5E",
			x"0000" when x"2F5F",
			x"0000" when x"2F60",
			x"0000" when x"2F61",
			x"0000" when x"2F62",
			x"0000" when x"2F63",
			x"0000" when x"2F64",
			x"0000" when x"2F65",
			x"0000" when x"2F66",
			x"0000" when x"2F67",
			x"0000" when x"2F68",
			x"0000" when x"2F69",
			x"0000" when x"2F6A",
			x"0000" when x"2F6B",
			x"0000" when x"2F6C",
			x"0000" when x"2F6D",
			x"0000" when x"2F6E",
			x"0000" when x"2F6F",
			x"0000" when x"2F70",
			x"0000" when x"2F71",
			x"0000" when x"2F72",
			x"0000" when x"2F73",
			x"0000" when x"2F74",
			x"0000" when x"2F75",
			x"0000" when x"2F76",
			x"0000" when x"2F77",
			x"0000" when x"2F78",
			x"0000" when x"2F79",
			x"0000" when x"2F7A",
			x"0000" when x"2F7B",
			x"0000" when x"2F7C",
			x"0000" when x"2F7D",
			x"0000" when x"2F7E",
			x"0000" when x"2F7F",
			x"0000" when x"2F80",
			x"0000" when x"2F81",
			x"0000" when x"2F82",
			x"0000" when x"2F83",
			x"0000" when x"2F84",
			x"0000" when x"2F85",
			x"0000" when x"2F86",
			x"0000" when x"2F87",
			x"0000" when x"2F88",
			x"0000" when x"2F89",
			x"0000" when x"2F8A",
			x"0000" when x"2F8B",
			x"0000" when x"2F8C",
			x"0000" when x"2F8D",
			x"0000" when x"2F8E",
			x"0000" when x"2F8F",
			x"0000" when x"2F90",
			x"0000" when x"2F91",
			x"0000" when x"2F92",
			x"0000" when x"2F93",
			x"0000" when x"2F94",
			x"0000" when x"2F95",
			x"0000" when x"2F96",
			x"0000" when x"2F97",
			x"0000" when x"2F98",
			x"0000" when x"2F99",
			x"0000" when x"2F9A",
			x"0000" when x"2F9B",
			x"0000" when x"2F9C",
			x"0000" when x"2F9D",
			x"0000" when x"2F9E",
			x"0000" when x"2F9F",
			x"0000" when x"2FA0",
			x"0000" when x"2FA1",
			x"0000" when x"2FA2",
			x"0000" when x"2FA3",
			x"0000" when x"2FA4",
			x"0000" when x"2FA5",
			x"0000" when x"2FA6",
			x"0000" when x"2FA7",
			x"0000" when x"2FA8",
			x"0000" when x"2FA9",
			x"0000" when x"2FAA",
			x"0000" when x"2FAB",
			x"0000" when x"2FAC",
			x"0000" when x"2FAD",
			x"0000" when x"2FAE",
			x"0000" when x"2FAF",
			x"0000" when x"2FB0",
			x"0000" when x"2FB1",
			x"0000" when x"2FB2",
			x"0000" when x"2FB3",
			x"0000" when x"2FB4",
			x"0000" when x"2FB5",
			x"0000" when x"2FB6",
			x"0000" when x"2FB7",
			x"0000" when x"2FB8",
			x"0000" when x"2FB9",
			x"0000" when x"2FBA",
			x"0000" when x"2FBB",
			x"0000" when x"2FBC",
			x"0000" when x"2FBD",
			x"0000" when x"2FBE",
			x"0000" when x"2FBF",
			x"0000" when x"2FC0",
			x"0000" when x"2FC1",
			x"0000" when x"2FC2",
			x"0000" when x"2FC3",
			x"0000" when x"2FC4",
			x"0000" when x"2FC5",
			x"0000" when x"2FC6",
			x"0000" when x"2FC7",
			x"0000" when x"2FC8",
			x"0000" when x"2FC9",
			x"0000" when x"2FCA",
			x"0000" when x"2FCB",
			x"0000" when x"2FCC",
			x"0000" when x"2FCD",
			x"0000" when x"2FCE",
			x"0000" when x"2FCF",
			x"0000" when x"2FD0",
			x"0000" when x"2FD1",
			x"0000" when x"2FD2",
			x"0000" when x"2FD3",
			x"0000" when x"2FD4",
			x"0000" when x"2FD5",
			x"0000" when x"2FD6",
			x"0000" when x"2FD7",
			x"0000" when x"2FD8",
			x"0000" when x"2FD9",
			x"0000" when x"2FDA",
			x"0000" when x"2FDB",
			x"0000" when x"2FDC",
			x"0000" when x"2FDD",
			x"0000" when x"2FDE",
			x"0000" when x"2FDF",
			x"0000" when x"2FE0",
			x"0000" when x"2FE1",
			x"0000" when x"2FE2",
			x"0000" when x"2FE3",
			x"0000" when x"2FE4",
			x"0000" when x"2FE5",
			x"0000" when x"2FE6",
			x"0000" when x"2FE7",
			x"0000" when x"2FE8",
			x"0000" when x"2FE9",
			x"0000" when x"2FEA",
			x"0000" when x"2FEB",
			x"0000" when x"2FEC",
			x"0000" when x"2FED",
			x"0000" when x"2FEE",
			x"0000" when x"2FEF",
			x"0000" when x"2FF0",
			x"0000" when x"2FF1",
			x"0000" when x"2FF2",
			x"0000" when x"2FF3",
			x"0000" when x"2FF4",
			x"0000" when x"2FF5",
			x"0000" when x"2FF6",
			x"0000" when x"2FF7",
			x"0000" when x"2FF8",
			x"0000" when x"2FF9",
			x"0000" when x"2FFA",
			x"0000" when x"2FFB",
			x"0000" when x"2FFC",
			x"0000" when x"2FFD",
			x"0000" when x"2FFE",
			x"0000" when x"2FFF",
			x"0000" when x"3000",
			x"0000" when x"3001",
			x"0000" when x"3002",
			x"0000" when x"3003",
			x"0000" when x"3004",
			x"0000" when x"3005",
			x"0000" when x"3006",
			x"0000" when x"3007",
			x"0000" when x"3008",
			x"0000" when x"3009",
			x"0000" when x"300A",
			x"0000" when x"300B",
			x"0000" when x"300C",
			x"0000" when x"300D",
			x"0000" when x"300E",
			x"0000" when x"300F",
			x"0000" when x"3010",
			x"0000" when x"3011",
			x"0000" when x"3012",
			x"0000" when x"3013",
			x"0000" when x"3014",
			x"0000" when x"3015",
			x"0000" when x"3016",
			x"0000" when x"3017",
			x"0000" when x"3018",
			x"0000" when x"3019",
			x"0000" when x"301A",
			x"0000" when x"301B",
			x"0000" when x"301C",
			x"0000" when x"301D",
			x"0000" when x"301E",
			x"0000" when x"301F",
			x"0000" when x"3020",
			x"0000" when x"3021",
			x"0000" when x"3022",
			x"0000" when x"3023",
			x"0000" when x"3024",
			x"0000" when x"3025",
			x"0000" when x"3026",
			x"0000" when x"3027",
			x"0000" when x"3028",
			x"0000" when x"3029",
			x"0000" when x"302A",
			x"0000" when x"302B",
			x"0000" when x"302C",
			x"0000" when x"302D",
			x"0000" when x"302E",
			x"0000" when x"302F",
			x"0000" when x"3030",
			x"0000" when x"3031",
			x"0000" when x"3032",
			x"0000" when x"3033",
			x"0000" when x"3034",
			x"0000" when x"3035",
			x"0000" when x"3036",
			x"0000" when x"3037",
			x"0000" when x"3038",
			x"0000" when x"3039",
			x"0000" when x"303A",
			x"0000" when x"303B",
			x"0000" when x"303C",
			x"0000" when x"303D",
			x"0000" when x"303E",
			x"0000" when x"303F",
			x"0000" when x"3040",
			x"0000" when x"3041",
			x"0000" when x"3042",
			x"0000" when x"3043",
			x"0000" when x"3044",
			x"0000" when x"3045",
			x"0000" when x"3046",
			x"0000" when x"3047",
			x"0000" when x"3048",
			x"0000" when x"3049",
			x"0000" when x"304A",
			x"0000" when x"304B",
			x"0000" when x"304C",
			x"0000" when x"304D",
			x"0000" when x"304E",
			x"0000" when x"304F",
			x"0000" when x"3050",
			x"0000" when x"3051",
			x"0000" when x"3052",
			x"0000" when x"3053",
			x"0000" when x"3054",
			x"0000" when x"3055",
			x"0000" when x"3056",
			x"0000" when x"3057",
			x"0000" when x"3058",
			x"0000" when x"3059",
			x"0000" when x"305A",
			x"0000" when x"305B",
			x"0000" when x"305C",
			x"0000" when x"305D",
			x"0000" when x"305E",
			x"0000" when x"305F",
			x"0000" when x"3060",
			x"0000" when x"3061",
			x"0000" when x"3062",
			x"0000" when x"3063",
			x"0000" when x"3064",
			x"0000" when x"3065",
			x"0000" when x"3066",
			x"0000" when x"3067",
			x"0000" when x"3068",
			x"0000" when x"3069",
			x"0000" when x"306A",
			x"0000" when x"306B",
			x"0000" when x"306C",
			x"0000" when x"306D",
			x"0000" when x"306E",
			x"0000" when x"306F",
			x"0000" when x"3070",
			x"0000" when x"3071",
			x"0000" when x"3072",
			x"0000" when x"3073",
			x"0000" when x"3074",
			x"0000" when x"3075",
			x"0000" when x"3076",
			x"0000" when x"3077",
			x"0000" when x"3078",
			x"0000" when x"3079",
			x"0000" when x"307A",
			x"0000" when x"307B",
			x"0000" when x"307C",
			x"0000" when x"307D",
			x"0000" when x"307E",
			x"0000" when x"307F",
			x"0000" when x"3080",
			x"0000" when x"3081",
			x"0000" when x"3082",
			x"0000" when x"3083",
			x"0000" when x"3084",
			x"0000" when x"3085",
			x"0000" when x"3086",
			x"0000" when x"3087",
			x"0000" when x"3088",
			x"0000" when x"3089",
			x"0000" when x"308A",
			x"0000" when x"308B",
			x"0000" when x"308C",
			x"0000" when x"308D",
			x"0000" when x"308E",
			x"0000" when x"308F",
			x"0000" when x"3090",
			x"0000" when x"3091",
			x"0000" when x"3092",
			x"0000" when x"3093",
			x"0000" when x"3094",
			x"0000" when x"3095",
			x"0000" when x"3096",
			x"0000" when x"3097",
			x"0000" when x"3098",
			x"0000" when x"3099",
			x"0000" when x"309A",
			x"0000" when x"309B",
			x"0000" when x"309C",
			x"0000" when x"309D",
			x"0000" when x"309E",
			x"0000" when x"309F",
			x"0000" when x"30A0",
			x"0000" when x"30A1",
			x"0000" when x"30A2",
			x"0000" when x"30A3",
			x"0000" when x"30A4",
			x"0000" when x"30A5",
			x"0000" when x"30A6",
			x"0000" when x"30A7",
			x"0000" when x"30A8",
			x"0000" when x"30A9",
			x"0000" when x"30AA",
			x"0000" when x"30AB",
			x"0000" when x"30AC",
			x"0000" when x"30AD",
			x"0000" when x"30AE",
			x"0000" when x"30AF",
			x"0000" when x"30B0",
			x"0000" when x"30B1",
			x"0000" when x"30B2",
			x"0000" when x"30B3",
			x"0000" when x"30B4",
			x"0000" when x"30B5",
			x"0000" when x"30B6",
			x"0000" when x"30B7",
			x"0000" when x"30B8",
			x"0000" when x"30B9",
			x"0000" when x"30BA",
			x"0000" when x"30BB",
			x"0000" when x"30BC",
			x"0000" when x"30BD",
			x"0000" when x"30BE",
			x"0000" when x"30BF",
			x"0000" when x"30C0",
			x"0000" when x"30C1",
			x"0000" when x"30C2",
			x"0000" when x"30C3",
			x"0000" when x"30C4",
			x"0000" when x"30C5",
			x"0000" when x"30C6",
			x"0000" when x"30C7",
			x"0000" when x"30C8",
			x"0000" when x"30C9",
			x"0000" when x"30CA",
			x"0000" when x"30CB",
			x"0000" when x"30CC",
			x"0000" when x"30CD",
			x"0000" when x"30CE",
			x"0000" when x"30CF",
			x"0000" when x"30D0",
			x"0000" when x"30D1",
			x"0000" when x"30D2",
			x"0000" when x"30D3",
			x"0000" when x"30D4",
			x"0000" when x"30D5",
			x"0000" when x"30D6",
			x"0000" when x"30D7",
			x"0000" when x"30D8",
			x"0000" when x"30D9",
			x"0000" when x"30DA",
			x"0000" when x"30DB",
			x"0000" when x"30DC",
			x"0000" when x"30DD",
			x"0000" when x"30DE",
			x"0000" when x"30DF",
			x"0000" when x"30E0",
			x"0000" when x"30E1",
			x"0000" when x"30E2",
			x"0000" when x"30E3",
			x"0000" when x"30E4",
			x"0000" when x"30E5",
			x"0000" when x"30E6",
			x"0000" when x"30E7",
			x"0000" when x"30E8",
			x"0000" when x"30E9",
			x"0000" when x"30EA",
			x"0000" when x"30EB",
			x"0000" when x"30EC",
			x"0000" when x"30ED",
			x"0000" when x"30EE",
			x"0000" when x"30EF",
			x"0000" when x"30F0",
			x"0000" when x"30F1",
			x"0000" when x"30F2",
			x"0000" when x"30F3",
			x"0000" when x"30F4",
			x"0000" when x"30F5",
			x"0000" when x"30F6",
			x"0000" when x"30F7",
			x"0000" when x"30F8",
			x"0000" when x"30F9",
			x"0000" when x"30FA",
			x"0000" when x"30FB",
			x"0000" when x"30FC",
			x"0000" when x"30FD",
			x"0000" when x"30FE",
			x"0000" when x"30FF",
			x"0000" when x"3100",
			x"0000" when x"3101",
			x"0000" when x"3102",
			x"0000" when x"3103",
			x"0000" when x"3104",
			x"0000" when x"3105",
			x"0000" when x"3106",
			x"0000" when x"3107",
			x"0000" when x"3108",
			x"0000" when x"3109",
			x"0000" when x"310A",
			x"0000" when x"310B",
			x"0000" when x"310C",
			x"0000" when x"310D",
			x"0000" when x"310E",
			x"0000" when x"310F",
			x"0000" when x"3110",
			x"0000" when x"3111",
			x"0000" when x"3112",
			x"0000" when x"3113",
			x"0000" when x"3114",
			x"0000" when x"3115",
			x"0000" when x"3116",
			x"0000" when x"3117",
			x"0000" when x"3118",
			x"0000" when x"3119",
			x"0000" when x"311A",
			x"0000" when x"311B",
			x"0000" when x"311C",
			x"0000" when x"311D",
			x"0000" when x"311E",
			x"0000" when x"311F",
			x"0000" when x"3120",
			x"0000" when x"3121",
			x"0000" when x"3122",
			x"0000" when x"3123",
			x"0000" when x"3124",
			x"0000" when x"3125",
			x"0000" when x"3126",
			x"0000" when x"3127",
			x"0000" when x"3128",
			x"0000" when x"3129",
			x"0000" when x"312A",
			x"0000" when x"312B",
			x"0000" when x"312C",
			x"0000" when x"312D",
			x"0000" when x"312E",
			x"0000" when x"312F",
			x"0000" when x"3130",
			x"0000" when x"3131",
			x"0000" when x"3132",
			x"0000" when x"3133",
			x"0000" when x"3134",
			x"0000" when x"3135",
			x"0000" when x"3136",
			x"0000" when x"3137",
			x"0000" when x"3138",
			x"0000" when x"3139",
			x"0000" when x"313A",
			x"0000" when x"313B",
			x"0000" when x"313C",
			x"0000" when x"313D",
			x"0000" when x"313E",
			x"0000" when x"313F",
			x"0000" when x"3140",
			x"0000" when x"3141",
			x"0000" when x"3142",
			x"0000" when x"3143",
			x"0000" when x"3144",
			x"0000" when x"3145",
			x"0000" when x"3146",
			x"0000" when x"3147",
			x"0000" when x"3148",
			x"0000" when x"3149",
			x"0000" when x"314A",
			x"0000" when x"314B",
			x"0000" when x"314C",
			x"0000" when x"314D",
			x"0000" when x"314E",
			x"0000" when x"314F",
			x"0000" when x"3150",
			x"0000" when x"3151",
			x"0000" when x"3152",
			x"0000" when x"3153",
			x"0000" when x"3154",
			x"0000" when x"3155",
			x"0000" when x"3156",
			x"0000" when x"3157",
			x"0000" when x"3158",
			x"0000" when x"3159",
			x"0000" when x"315A",
			x"0000" when x"315B",
			x"0000" when x"315C",
			x"0000" when x"315D",
			x"0000" when x"315E",
			x"0000" when x"315F",
			x"0000" when x"3160",
			x"0000" when x"3161",
			x"0000" when x"3162",
			x"0000" when x"3163",
			x"0000" when x"3164",
			x"0000" when x"3165",
			x"0000" when x"3166",
			x"0000" when x"3167",
			x"0000" when x"3168",
			x"0000" when x"3169",
			x"0000" when x"316A",
			x"0000" when x"316B",
			x"0000" when x"316C",
			x"0000" when x"316D",
			x"0000" when x"316E",
			x"0000" when x"316F",
			x"0000" when x"3170",
			x"0000" when x"3171",
			x"0000" when x"3172",
			x"0000" when x"3173",
			x"0000" when x"3174",
			x"0000" when x"3175",
			x"0000" when x"3176",
			x"0000" when x"3177",
			x"0000" when x"3178",
			x"0000" when x"3179",
			x"0000" when x"317A",
			x"0000" when x"317B",
			x"0000" when x"317C",
			x"0000" when x"317D",
			x"0000" when x"317E",
			x"0000" when x"317F",
			x"0000" when x"3180",
			x"0000" when x"3181",
			x"0000" when x"3182",
			x"0000" when x"3183",
			x"0000" when x"3184",
			x"0000" when x"3185",
			x"0000" when x"3186",
			x"0000" when x"3187",
			x"0000" when x"3188",
			x"0000" when x"3189",
			x"0000" when x"318A",
			x"0000" when x"318B",
			x"0000" when x"318C",
			x"0000" when x"318D",
			x"0000" when x"318E",
			x"0000" when x"318F",
			x"0000" when x"3190",
			x"0000" when x"3191",
			x"0000" when x"3192",
			x"0000" when x"3193",
			x"0000" when x"3194",
			x"0000" when x"3195",
			x"0000" when x"3196",
			x"0000" when x"3197",
			x"0000" when x"3198",
			x"0000" when x"3199",
			x"0000" when x"319A",
			x"0000" when x"319B",
			x"0000" when x"319C",
			x"0000" when x"319D",
			x"0000" when x"319E",
			x"0000" when x"319F",
			x"0000" when x"31A0",
			x"0000" when x"31A1",
			x"0000" when x"31A2",
			x"0000" when x"31A3",
			x"0000" when x"31A4",
			x"0000" when x"31A5",
			x"0000" when x"31A6",
			x"0000" when x"31A7",
			x"0000" when x"31A8",
			x"0000" when x"31A9",
			x"0000" when x"31AA",
			x"0000" when x"31AB",
			x"0000" when x"31AC",
			x"0000" when x"31AD",
			x"0000" when x"31AE",
			x"0000" when x"31AF",
			x"0000" when x"31B0",
			x"0000" when x"31B1",
			x"0000" when x"31B2",
			x"0000" when x"31B3",
			x"0000" when x"31B4",
			x"0000" when x"31B5",
			x"0000" when x"31B6",
			x"0000" when x"31B7",
			x"0000" when x"31B8",
			x"0000" when x"31B9",
			x"0000" when x"31BA",
			x"0000" when x"31BB",
			x"0000" when x"31BC",
			x"0000" when x"31BD",
			x"0000" when x"31BE",
			x"0000" when x"31BF",
			x"0000" when x"31C0",
			x"0000" when x"31C1",
			x"0000" when x"31C2",
			x"0000" when x"31C3",
			x"0000" when x"31C4",
			x"0000" when x"31C5",
			x"0000" when x"31C6",
			x"0000" when x"31C7",
			x"0000" when x"31C8",
			x"0000" when x"31C9",
			x"0000" when x"31CA",
			x"0000" when x"31CB",
			x"0000" when x"31CC",
			x"0000" when x"31CD",
			x"0000" when x"31CE",
			x"0000" when x"31CF",
			x"0000" when x"31D0",
			x"0000" when x"31D1",
			x"0000" when x"31D2",
			x"0000" when x"31D3",
			x"0000" when x"31D4",
			x"0000" when x"31D5",
			x"0000" when x"31D6",
			x"0000" when x"31D7",
			x"0000" when x"31D8",
			x"0000" when x"31D9",
			x"0000" when x"31DA",
			x"0000" when x"31DB",
			x"0000" when x"31DC",
			x"0000" when x"31DD",
			x"0000" when x"31DE",
			x"0000" when x"31DF",
			x"0000" when x"31E0",
			x"0000" when x"31E1",
			x"0000" when x"31E2",
			x"0000" when x"31E3",
			x"0000" when x"31E4",
			x"0000" when x"31E5",
			x"0000" when x"31E6",
			x"0000" when x"31E7",
			x"0000" when x"31E8",
			x"0000" when x"31E9",
			x"0000" when x"31EA",
			x"0000" when x"31EB",
			x"0000" when x"31EC",
			x"0000" when x"31ED",
			x"0000" when x"31EE",
			x"0000" when x"31EF",
			x"0000" when x"31F0",
			x"0000" when x"31F1",
			x"0000" when x"31F2",
			x"0000" when x"31F3",
			x"0000" when x"31F4",
			x"0000" when x"31F5",
			x"0000" when x"31F6",
			x"0000" when x"31F7",
			x"0000" when x"31F8",
			x"0000" when x"31F9",
			x"0000" when x"31FA",
			x"0000" when x"31FB",
			x"0000" when x"31FC",
			x"0000" when x"31FD",
			x"0000" when x"31FE",
			x"0000" when x"31FF",
			x"0000" when x"3200",
			x"0000" when x"3201",
			x"0000" when x"3202",
			x"0000" when x"3203",
			x"0000" when x"3204",
			x"0000" when x"3205",
			x"0000" when x"3206",
			x"0000" when x"3207",
			x"0000" when x"3208",
			x"0000" when x"3209",
			x"0000" when x"320A",
			x"0000" when x"320B",
			x"0000" when x"320C",
			x"0000" when x"320D",
			x"0000" when x"320E",
			x"0000" when x"320F",
			x"0000" when x"3210",
			x"0000" when x"3211",
			x"0000" when x"3212",
			x"0000" when x"3213",
			x"0000" when x"3214",
			x"0000" when x"3215",
			x"0000" when x"3216",
			x"0000" when x"3217",
			x"0000" when x"3218",
			x"0000" when x"3219",
			x"0000" when x"321A",
			x"0000" when x"321B",
			x"0000" when x"321C",
			x"0000" when x"321D",
			x"0000" when x"321E",
			x"0000" when x"321F",
			x"0000" when x"3220",
			x"0000" when x"3221",
			x"0000" when x"3222",
			x"0000" when x"3223",
			x"0000" when x"3224",
			x"0000" when x"3225",
			x"0000" when x"3226",
			x"0000" when x"3227",
			x"0000" when x"3228",
			x"0000" when x"3229",
			x"0000" when x"322A",
			x"0000" when x"322B",
			x"0000" when x"322C",
			x"0000" when x"322D",
			x"0000" when x"322E",
			x"0000" when x"322F",
			x"0000" when x"3230",
			x"0000" when x"3231",
			x"0000" when x"3232",
			x"0000" when x"3233",
			x"0000" when x"3234",
			x"0000" when x"3235",
			x"0000" when x"3236",
			x"0000" when x"3237",
			x"0000" when x"3238",
			x"0000" when x"3239",
			x"0000" when x"323A",
			x"0000" when x"323B",
			x"0000" when x"323C",
			x"0000" when x"323D",
			x"0000" when x"323E",
			x"0000" when x"323F",
			x"0000" when x"3240",
			x"0000" when x"3241",
			x"0000" when x"3242",
			x"0000" when x"3243",
			x"0000" when x"3244",
			x"0000" when x"3245",
			x"0000" when x"3246",
			x"0000" when x"3247",
			x"0000" when x"3248",
			x"0000" when x"3249",
			x"0000" when x"324A",
			x"0000" when x"324B",
			x"0000" when x"324C",
			x"0000" when x"324D",
			x"0000" when x"324E",
			x"0000" when x"324F",
			x"0000" when x"3250",
			x"0000" when x"3251",
			x"0000" when x"3252",
			x"0000" when x"3253",
			x"0000" when x"3254",
			x"0000" when x"3255",
			x"0000" when x"3256",
			x"0000" when x"3257",
			x"0000" when x"3258",
			x"0000" when x"3259",
			x"0000" when x"325A",
			x"0000" when x"325B",
			x"0000" when x"325C",
			x"0000" when x"325D",
			x"0000" when x"325E",
			x"0000" when x"325F",
			x"0000" when x"3260",
			x"0000" when x"3261",
			x"0000" when x"3262",
			x"0000" when x"3263",
			x"0000" when x"3264",
			x"0000" when x"3265",
			x"0000" when x"3266",
			x"0000" when x"3267",
			x"0000" when x"3268",
			x"0000" when x"3269",
			x"0000" when x"326A",
			x"0000" when x"326B",
			x"0000" when x"326C",
			x"0000" when x"326D",
			x"0000" when x"326E",
			x"0000" when x"326F",
			x"0000" when x"3270",
			x"0000" when x"3271",
			x"0000" when x"3272",
			x"0000" when x"3273",
			x"0000" when x"3274",
			x"0000" when x"3275",
			x"0000" when x"3276",
			x"0000" when x"3277",
			x"0000" when x"3278",
			x"0000" when x"3279",
			x"0000" when x"327A",
			x"0000" when x"327B",
			x"0000" when x"327C",
			x"0000" when x"327D",
			x"0000" when x"327E",
			x"0000" when x"327F",
			x"0000" when x"3280",
			x"0000" when x"3281",
			x"0000" when x"3282",
			x"0000" when x"3283",
			x"0000" when x"3284",
			x"0000" when x"3285",
			x"0000" when x"3286",
			x"0000" when x"3287",
			x"0000" when x"3288",
			x"0000" when x"3289",
			x"0000" when x"328A",
			x"0000" when x"328B",
			x"0000" when x"328C",
			x"0000" when x"328D",
			x"0000" when x"328E",
			x"0000" when x"328F",
			x"0000" when x"3290",
			x"0000" when x"3291",
			x"0000" when x"3292",
			x"0000" when x"3293",
			x"0000" when x"3294",
			x"0000" when x"3295",
			x"0000" when x"3296",
			x"0000" when x"3297",
			x"0000" when x"3298",
			x"0000" when x"3299",
			x"0000" when x"329A",
			x"0000" when x"329B",
			x"0000" when x"329C",
			x"0000" when x"329D",
			x"0000" when x"329E",
			x"0000" when x"329F",
			x"0000" when x"32A0",
			x"0000" when x"32A1",
			x"0000" when x"32A2",
			x"0000" when x"32A3",
			x"0000" when x"32A4",
			x"0000" when x"32A5",
			x"0000" when x"32A6",
			x"0000" when x"32A7",
			x"0000" when x"32A8",
			x"0000" when x"32A9",
			x"0000" when x"32AA",
			x"0000" when x"32AB",
			x"0000" when x"32AC",
			x"0000" when x"32AD",
			x"0000" when x"32AE",
			x"0000" when x"32AF",
			x"0000" when x"32B0",
			x"0000" when x"32B1",
			x"0000" when x"32B2",
			x"0000" when x"32B3",
			x"0000" when x"32B4",
			x"0000" when x"32B5",
			x"0000" when x"32B6",
			x"0000" when x"32B7",
			x"0000" when x"32B8",
			x"0000" when x"32B9",
			x"0000" when x"32BA",
			x"0000" when x"32BB",
			x"0000" when x"32BC",
			x"0000" when x"32BD",
			x"0000" when x"32BE",
			x"0000" when x"32BF",
			x"0000" when x"32C0",
			x"0000" when x"32C1",
			x"0000" when x"32C2",
			x"0000" when x"32C3",
			x"0000" when x"32C4",
			x"0000" when x"32C5",
			x"0000" when x"32C6",
			x"0000" when x"32C7",
			x"0000" when x"32C8",
			x"0000" when x"32C9",
			x"0000" when x"32CA",
			x"0000" when x"32CB",
			x"0000" when x"32CC",
			x"0000" when x"32CD",
			x"0000" when x"32CE",
			x"0000" when x"32CF",
			x"0000" when x"32D0",
			x"0000" when x"32D1",
			x"0000" when x"32D2",
			x"0000" when x"32D3",
			x"0000" when x"32D4",
			x"0000" when x"32D5",
			x"0000" when x"32D6",
			x"0000" when x"32D7",
			x"0000" when x"32D8",
			x"0000" when x"32D9",
			x"0000" when x"32DA",
			x"0000" when x"32DB",
			x"0000" when x"32DC",
			x"0000" when x"32DD",
			x"0000" when x"32DE",
			x"0000" when x"32DF",
			x"0000" when x"32E0",
			x"0000" when x"32E1",
			x"0000" when x"32E2",
			x"0000" when x"32E3",
			x"0000" when x"32E4",
			x"0000" when x"32E5",
			x"0000" when x"32E6",
			x"0000" when x"32E7",
			x"0000" when x"32E8",
			x"0000" when x"32E9",
			x"0000" when x"32EA",
			x"0000" when x"32EB",
			x"0000" when x"32EC",
			x"0000" when x"32ED",
			x"0000" when x"32EE",
			x"0000" when x"32EF",
			x"0000" when x"32F0",
			x"0000" when x"32F1",
			x"0000" when x"32F2",
			x"0000" when x"32F3",
			x"0000" when x"32F4",
			x"0000" when x"32F5",
			x"0000" when x"32F6",
			x"0000" when x"32F7",
			x"0000" when x"32F8",
			x"0000" when x"32F9",
			x"0000" when x"32FA",
			x"0000" when x"32FB",
			x"0000" when x"32FC",
			x"0000" when x"32FD",
			x"0000" when x"32FE",
			x"0000" when x"32FF",
			x"0000" when x"3300",
			x"0000" when x"3301",
			x"0000" when x"3302",
			x"0000" when x"3303",
			x"0000" when x"3304",
			x"0000" when x"3305",
			x"0000" when x"3306",
			x"0000" when x"3307",
			x"0000" when x"3308",
			x"0000" when x"3309",
			x"0000" when x"330A",
			x"0000" when x"330B",
			x"0000" when x"330C",
			x"0000" when x"330D",
			x"0000" when x"330E",
			x"0000" when x"330F",
			x"0000" when x"3310",
			x"0000" when x"3311",
			x"0000" when x"3312",
			x"0000" when x"3313",
			x"0000" when x"3314",
			x"0000" when x"3315",
			x"0000" when x"3316",
			x"0000" when x"3317",
			x"0000" when x"3318",
			x"0000" when x"3319",
			x"0000" when x"331A",
			x"0000" when x"331B",
			x"0000" when x"331C",
			x"0000" when x"331D",
			x"0000" when x"331E",
			x"0000" when x"331F",
			x"0000" when x"3320",
			x"0000" when x"3321",
			x"0000" when x"3322",
			x"0000" when x"3323",
			x"0000" when x"3324",
			x"0000" when x"3325",
			x"0000" when x"3326",
			x"0000" when x"3327",
			x"0000" when x"3328",
			x"0000" when x"3329",
			x"0000" when x"332A",
			x"0000" when x"332B",
			x"0000" when x"332C",
			x"0000" when x"332D",
			x"0000" when x"332E",
			x"0000" when x"332F",
			x"0000" when x"3330",
			x"0000" when x"3331",
			x"0000" when x"3332",
			x"0000" when x"3333",
			x"0000" when x"3334",
			x"0000" when x"3335",
			x"0000" when x"3336",
			x"0000" when x"3337",
			x"0000" when x"3338",
			x"0000" when x"3339",
			x"0000" when x"333A",
			x"0000" when x"333B",
			x"0000" when x"333C",
			x"0000" when x"333D",
			x"0000" when x"333E",
			x"0000" when x"333F",
			x"0000" when x"3340",
			x"0000" when x"3341",
			x"0000" when x"3342",
			x"0000" when x"3343",
			x"0000" when x"3344",
			x"0000" when x"3345",
			x"0000" when x"3346",
			x"0000" when x"3347",
			x"0000" when x"3348",
			x"0000" when x"3349",
			x"0000" when x"334A",
			x"0000" when x"334B",
			x"0000" when x"334C",
			x"0000" when x"334D",
			x"0000" when x"334E",
			x"0000" when x"334F",
			x"0000" when x"3350",
			x"0000" when x"3351",
			x"0000" when x"3352",
			x"0000" when x"3353",
			x"0000" when x"3354",
			x"0000" when x"3355",
			x"0000" when x"3356",
			x"0000" when x"3357",
			x"0000" when x"3358",
			x"0000" when x"3359",
			x"0000" when x"335A",
			x"0000" when x"335B",
			x"0000" when x"335C",
			x"0000" when x"335D",
			x"0000" when x"335E",
			x"0000" when x"335F",
			x"0000" when x"3360",
			x"0000" when x"3361",
			x"0000" when x"3362",
			x"0000" when x"3363",
			x"0000" when x"3364",
			x"0000" when x"3365",
			x"0000" when x"3366",
			x"0000" when x"3367",
			x"0000" when x"3368",
			x"0000" when x"3369",
			x"0000" when x"336A",
			x"0000" when x"336B",
			x"0000" when x"336C",
			x"0000" when x"336D",
			x"0000" when x"336E",
			x"0000" when x"336F",
			x"0000" when x"3370",
			x"0000" when x"3371",
			x"0000" when x"3372",
			x"0000" when x"3373",
			x"0000" when x"3374",
			x"0000" when x"3375",
			x"0000" when x"3376",
			x"0000" when x"3377",
			x"0000" when x"3378",
			x"0000" when x"3379",
			x"0000" when x"337A",
			x"0000" when x"337B",
			x"0000" when x"337C",
			x"0000" when x"337D",
			x"0000" when x"337E",
			x"0000" when x"337F",
			x"0000" when x"3380",
			x"0000" when x"3381",
			x"0000" when x"3382",
			x"0000" when x"3383",
			x"0000" when x"3384",
			x"0000" when x"3385",
			x"0000" when x"3386",
			x"0000" when x"3387",
			x"0000" when x"3388",
			x"0000" when x"3389",
			x"0000" when x"338A",
			x"0000" when x"338B",
			x"0000" when x"338C",
			x"0000" when x"338D",
			x"0000" when x"338E",
			x"0000" when x"338F",
			x"0000" when x"3390",
			x"0000" when x"3391",
			x"0000" when x"3392",
			x"0000" when x"3393",
			x"0000" when x"3394",
			x"0000" when x"3395",
			x"0000" when x"3396",
			x"0000" when x"3397",
			x"0000" when x"3398",
			x"0000" when x"3399",
			x"0000" when x"339A",
			x"0000" when x"339B",
			x"0000" when x"339C",
			x"0000" when x"339D",
			x"0000" when x"339E",
			x"0000" when x"339F",
			x"0000" when x"33A0",
			x"0000" when x"33A1",
			x"0000" when x"33A2",
			x"0000" when x"33A3",
			x"0000" when x"33A4",
			x"0000" when x"33A5",
			x"0000" when x"33A6",
			x"0000" when x"33A7",
			x"0000" when x"33A8",
			x"0000" when x"33A9",
			x"0000" when x"33AA",
			x"0000" when x"33AB",
			x"0000" when x"33AC",
			x"0000" when x"33AD",
			x"0000" when x"33AE",
			x"0000" when x"33AF",
			x"0000" when x"33B0",
			x"0000" when x"33B1",
			x"0000" when x"33B2",
			x"0000" when x"33B3",
			x"0000" when x"33B4",
			x"0000" when x"33B5",
			x"0000" when x"33B6",
			x"0000" when x"33B7",
			x"0000" when x"33B8",
			x"0000" when x"33B9",
			x"0000" when x"33BA",
			x"0000" when x"33BB",
			x"0000" when x"33BC",
			x"0000" when x"33BD",
			x"0000" when x"33BE",
			x"0000" when x"33BF",
			x"0000" when x"33C0",
			x"0000" when x"33C1",
			x"0000" when x"33C2",
			x"0000" when x"33C3",
			x"0000" when x"33C4",
			x"0000" when x"33C5",
			x"0000" when x"33C6",
			x"0000" when x"33C7",
			x"0000" when x"33C8",
			x"0000" when x"33C9",
			x"0000" when x"33CA",
			x"0000" when x"33CB",
			x"0000" when x"33CC",
			x"0000" when x"33CD",
			x"0000" when x"33CE",
			x"0000" when x"33CF",
			x"0000" when x"33D0",
			x"0000" when x"33D1",
			x"0000" when x"33D2",
			x"0000" when x"33D3",
			x"0000" when x"33D4",
			x"0000" when x"33D5",
			x"0000" when x"33D6",
			x"0000" when x"33D7",
			x"0000" when x"33D8",
			x"0000" when x"33D9",
			x"0000" when x"33DA",
			x"0000" when x"33DB",
			x"0000" when x"33DC",
			x"0000" when x"33DD",
			x"0000" when x"33DE",
			x"0000" when x"33DF",
			x"0000" when x"33E0",
			x"0000" when x"33E1",
			x"0000" when x"33E2",
			x"0000" when x"33E3",
			x"0000" when x"33E4",
			x"0000" when x"33E5",
			x"0000" when x"33E6",
			x"0000" when x"33E7",
			x"0000" when x"33E8",
			x"0000" when x"33E9",
			x"0000" when x"33EA",
			x"0000" when x"33EB",
			x"0000" when x"33EC",
			x"0000" when x"33ED",
			x"0000" when x"33EE",
			x"0000" when x"33EF",
			x"0000" when x"33F0",
			x"0000" when x"33F1",
			x"0000" when x"33F2",
			x"0000" when x"33F3",
			x"0000" when x"33F4",
			x"0000" when x"33F5",
			x"0000" when x"33F6",
			x"0000" when x"33F7",
			x"0000" when x"33F8",
			x"0000" when x"33F9",
			x"0000" when x"33FA",
			x"0000" when x"33FB",
			x"0000" when x"33FC",
			x"0000" when x"33FD",
			x"0000" when x"33FE",
			x"0000" when x"33FF",
			x"0000" when x"3400",
			x"0000" when x"3401",
			x"0000" when x"3402",
			x"0000" when x"3403",
			x"0000" when x"3404",
			x"0000" when x"3405",
			x"0000" when x"3406",
			x"0000" when x"3407",
			x"0000" when x"3408",
			x"0000" when x"3409",
			x"0000" when x"340A",
			x"0000" when x"340B",
			x"0000" when x"340C",
			x"0000" when x"340D",
			x"0000" when x"340E",
			x"0000" when x"340F",
			x"0000" when x"3410",
			x"0000" when x"3411",
			x"0000" when x"3412",
			x"0000" when x"3413",
			x"0000" when x"3414",
			x"0000" when x"3415",
			x"0000" when x"3416",
			x"0000" when x"3417",
			x"0000" when x"3418",
			x"0000" when x"3419",
			x"0000" when x"341A",
			x"0000" when x"341B",
			x"0000" when x"341C",
			x"0000" when x"341D",
			x"0000" when x"341E",
			x"0000" when x"341F",
			x"0000" when x"3420",
			x"0000" when x"3421",
			x"0000" when x"3422",
			x"0000" when x"3423",
			x"0000" when x"3424",
			x"0000" when x"3425",
			x"0000" when x"3426",
			x"0000" when x"3427",
			x"0000" when x"3428",
			x"0000" when x"3429",
			x"0000" when x"342A",
			x"0000" when x"342B",
			x"0000" when x"342C",
			x"0000" when x"342D",
			x"0000" when x"342E",
			x"0000" when x"342F",
			x"0000" when x"3430",
			x"0000" when x"3431",
			x"0000" when x"3432",
			x"0000" when x"3433",
			x"0000" when x"3434",
			x"0000" when x"3435",
			x"0000" when x"3436",
			x"0000" when x"3437",
			x"0000" when x"3438",
			x"0000" when x"3439",
			x"0000" when x"343A",
			x"0000" when x"343B",
			x"0000" when x"343C",
			x"0000" when x"343D",
			x"0000" when x"343E",
			x"0000" when x"343F",
			x"0000" when x"3440",
			x"0000" when x"3441",
			x"0000" when x"3442",
			x"0000" when x"3443",
			x"0000" when x"3444",
			x"0000" when x"3445",
			x"0000" when x"3446",
			x"0000" when x"3447",
			x"0000" when x"3448",
			x"0000" when x"3449",
			x"0000" when x"344A",
			x"0000" when x"344B",
			x"0000" when x"344C",
			x"0000" when x"344D",
			x"0000" when x"344E",
			x"0000" when x"344F",
			x"0000" when x"3450",
			x"0000" when x"3451",
			x"0000" when x"3452",
			x"0000" when x"3453",
			x"0000" when x"3454",
			x"0000" when x"3455",
			x"0000" when x"3456",
			x"0000" when x"3457",
			x"0000" when x"3458",
			x"0000" when x"3459",
			x"0000" when x"345A",
			x"0000" when x"345B",
			x"0000" when x"345C",
			x"0000" when x"345D",
			x"0000" when x"345E",
			x"0000" when x"345F",
			x"0000" when x"3460",
			x"0000" when x"3461",
			x"0000" when x"3462",
			x"0000" when x"3463",
			x"0000" when x"3464",
			x"0000" when x"3465",
			x"0000" when x"3466",
			x"0000" when x"3467",
			x"0000" when x"3468",
			x"0000" when x"3469",
			x"0000" when x"346A",
			x"0000" when x"346B",
			x"0000" when x"346C",
			x"0000" when x"346D",
			x"0000" when x"346E",
			x"0000" when x"346F",
			x"0000" when x"3470",
			x"0000" when x"3471",
			x"0000" when x"3472",
			x"0000" when x"3473",
			x"0000" when x"3474",
			x"0000" when x"3475",
			x"0000" when x"3476",
			x"0000" when x"3477",
			x"0000" when x"3478",
			x"0000" when x"3479",
			x"0000" when x"347A",
			x"0000" when x"347B",
			x"0000" when x"347C",
			x"0000" when x"347D",
			x"0000" when x"347E",
			x"0000" when x"347F",
			x"0000" when x"3480",
			x"0000" when x"3481",
			x"0000" when x"3482",
			x"0000" when x"3483",
			x"0000" when x"3484",
			x"0000" when x"3485",
			x"0000" when x"3486",
			x"0000" when x"3487",
			x"0000" when x"3488",
			x"0000" when x"3489",
			x"0000" when x"348A",
			x"0000" when x"348B",
			x"0000" when x"348C",
			x"0000" when x"348D",
			x"0000" when x"348E",
			x"0000" when x"348F",
			x"0000" when x"3490",
			x"0000" when x"3491",
			x"0000" when x"3492",
			x"0000" when x"3493",
			x"0000" when x"3494",
			x"0000" when x"3495",
			x"0000" when x"3496",
			x"0000" when x"3497",
			x"0000" when x"3498",
			x"0000" when x"3499",
			x"0000" when x"349A",
			x"0000" when x"349B",
			x"0000" when x"349C",
			x"0000" when x"349D",
			x"0000" when x"349E",
			x"0000" when x"349F",
			x"0000" when x"34A0",
			x"0000" when x"34A1",
			x"0000" when x"34A2",
			x"0000" when x"34A3",
			x"0000" when x"34A4",
			x"0000" when x"34A5",
			x"0000" when x"34A6",
			x"0000" when x"34A7",
			x"0000" when x"34A8",
			x"0000" when x"34A9",
			x"0000" when x"34AA",
			x"0000" when x"34AB",
			x"0000" when x"34AC",
			x"0000" when x"34AD",
			x"0000" when x"34AE",
			x"0000" when x"34AF",
			x"0000" when x"34B0",
			x"0000" when x"34B1",
			x"0000" when x"34B2",
			x"0000" when x"34B3",
			x"0000" when x"34B4",
			x"0000" when x"34B5",
			x"0000" when x"34B6",
			x"0000" when x"34B7",
			x"0000" when x"34B8",
			x"0000" when x"34B9",
			x"0000" when x"34BA",
			x"0000" when x"34BB",
			x"0000" when x"34BC",
			x"0000" when x"34BD",
			x"0000" when x"34BE",
			x"0000" when x"34BF",
			x"0000" when x"34C0",
			x"0000" when x"34C1",
			x"0000" when x"34C2",
			x"0000" when x"34C3",
			x"0000" when x"34C4",
			x"0000" when x"34C5",
			x"0000" when x"34C6",
			x"0000" when x"34C7",
			x"0000" when x"34C8",
			x"0000" when x"34C9",
			x"0000" when x"34CA",
			x"0000" when x"34CB",
			x"0000" when x"34CC",
			x"0000" when x"34CD",
			x"0000" when x"34CE",
			x"0000" when x"34CF",
			x"0000" when x"34D0",
			x"0000" when x"34D1",
			x"0000" when x"34D2",
			x"0000" when x"34D3",
			x"0000" when x"34D4",
			x"0000" when x"34D5",
			x"0000" when x"34D6",
			x"0000" when x"34D7",
			x"0000" when x"34D8",
			x"0000" when x"34D9",
			x"0000" when x"34DA",
			x"0000" when x"34DB",
			x"0000" when x"34DC",
			x"0000" when x"34DD",
			x"0000" when x"34DE",
			x"0000" when x"34DF",
			x"0000" when x"34E0",
			x"0000" when x"34E1",
			x"0000" when x"34E2",
			x"0000" when x"34E3",
			x"0000" when x"34E4",
			x"0000" when x"34E5",
			x"0000" when x"34E6",
			x"0000" when x"34E7",
			x"0000" when x"34E8",
			x"0000" when x"34E9",
			x"0000" when x"34EA",
			x"0000" when x"34EB",
			x"0000" when x"34EC",
			x"0000" when x"34ED",
			x"0000" when x"34EE",
			x"0000" when x"34EF",
			x"0000" when x"34F0",
			x"0000" when x"34F1",
			x"0000" when x"34F2",
			x"0000" when x"34F3",
			x"0000" when x"34F4",
			x"0000" when x"34F5",
			x"0000" when x"34F6",
			x"0000" when x"34F7",
			x"0000" when x"34F8",
			x"0000" when x"34F9",
			x"0000" when x"34FA",
			x"0000" when x"34FB",
			x"0000" when x"34FC",
			x"0000" when x"34FD",
			x"0000" when x"34FE",
			x"0000" when x"34FF",
			x"0000" when x"3500",
			x"0000" when x"3501",
			x"0000" when x"3502",
			x"0000" when x"3503",
			x"0000" when x"3504",
			x"0000" when x"3505",
			x"0000" when x"3506",
			x"0000" when x"3507",
			x"0000" when x"3508",
			x"0000" when x"3509",
			x"0000" when x"350A",
			x"0000" when x"350B",
			x"0000" when x"350C",
			x"0000" when x"350D",
			x"0000" when x"350E",
			x"0000" when x"350F",
			x"0000" when x"3510",
			x"0000" when x"3511",
			x"0000" when x"3512",
			x"0000" when x"3513",
			x"0000" when x"3514",
			x"0000" when x"3515",
			x"0000" when x"3516",
			x"0000" when x"3517",
			x"0000" when x"3518",
			x"0000" when x"3519",
			x"0000" when x"351A",
			x"0000" when x"351B",
			x"0000" when x"351C",
			x"0000" when x"351D",
			x"0000" when x"351E",
			x"0000" when x"351F",
			x"0000" when x"3520",
			x"0000" when x"3521",
			x"0000" when x"3522",
			x"0000" when x"3523",
			x"0000" when x"3524",
			x"0000" when x"3525",
			x"0000" when x"3526",
			x"0000" when x"3527",
			x"0000" when x"3528",
			x"0000" when x"3529",
			x"0000" when x"352A",
			x"0000" when x"352B",
			x"0000" when x"352C",
			x"0000" when x"352D",
			x"0000" when x"352E",
			x"0000" when x"352F",
			x"0000" when x"3530",
			x"0000" when x"3531",
			x"0000" when x"3532",
			x"0000" when x"3533",
			x"0000" when x"3534",
			x"0000" when x"3535",
			x"0000" when x"3536",
			x"0000" when x"3537",
			x"0000" when x"3538",
			x"0000" when x"3539",
			x"0000" when x"353A",
			x"0000" when x"353B",
			x"0000" when x"353C",
			x"0000" when x"353D",
			x"0000" when x"353E",
			x"0000" when x"353F",
			x"0000" when x"3540",
			x"0000" when x"3541",
			x"0000" when x"3542",
			x"0000" when x"3543",
			x"0000" when x"3544",
			x"0000" when x"3545",
			x"0000" when x"3546",
			x"0000" when x"3547",
			x"0000" when x"3548",
			x"0000" when x"3549",
			x"0000" when x"354A",
			x"0000" when x"354B",
			x"0000" when x"354C",
			x"0000" when x"354D",
			x"0000" when x"354E",
			x"0000" when x"354F",
			x"0000" when x"3550",
			x"0000" when x"3551",
			x"0000" when x"3552",
			x"0000" when x"3553",
			x"0000" when x"3554",
			x"0000" when x"3555",
			x"0000" when x"3556",
			x"0000" when x"3557",
			x"0000" when x"3558",
			x"0000" when x"3559",
			x"0000" when x"355A",
			x"0000" when x"355B",
			x"0000" when x"355C",
			x"0000" when x"355D",
			x"0000" when x"355E",
			x"0000" when x"355F",
			x"0000" when x"3560",
			x"0000" when x"3561",
			x"0000" when x"3562",
			x"0000" when x"3563",
			x"0000" when x"3564",
			x"0000" when x"3565",
			x"0000" when x"3566",
			x"0000" when x"3567",
			x"0000" when x"3568",
			x"0000" when x"3569",
			x"0000" when x"356A",
			x"0000" when x"356B",
			x"0000" when x"356C",
			x"0000" when x"356D",
			x"0000" when x"356E",
			x"0000" when x"356F",
			x"0000" when x"3570",
			x"0000" when x"3571",
			x"0000" when x"3572",
			x"0000" when x"3573",
			x"0000" when x"3574",
			x"0000" when x"3575",
			x"0000" when x"3576",
			x"0000" when x"3577",
			x"0000" when x"3578",
			x"0000" when x"3579",
			x"0000" when x"357A",
			x"0000" when x"357B",
			x"0000" when x"357C",
			x"0000" when x"357D",
			x"0000" when x"357E",
			x"0000" when x"357F",
			x"0000" when x"3580",
			x"0000" when x"3581",
			x"0000" when x"3582",
			x"0000" when x"3583",
			x"0000" when x"3584",
			x"0000" when x"3585",
			x"0000" when x"3586",
			x"0000" when x"3587",
			x"0000" when x"3588",
			x"0000" when x"3589",
			x"0000" when x"358A",
			x"0000" when x"358B",
			x"0000" when x"358C",
			x"0000" when x"358D",
			x"0000" when x"358E",
			x"0000" when x"358F",
			x"0000" when x"3590",
			x"0000" when x"3591",
			x"0000" when x"3592",
			x"0000" when x"3593",
			x"0000" when x"3594",
			x"0000" when x"3595",
			x"0000" when x"3596",
			x"0000" when x"3597",
			x"0000" when x"3598",
			x"0000" when x"3599",
			x"0000" when x"359A",
			x"0000" when x"359B",
			x"0000" when x"359C",
			x"0000" when x"359D",
			x"0000" when x"359E",
			x"0000" when x"359F",
			x"0000" when x"35A0",
			x"0000" when x"35A1",
			x"0000" when x"35A2",
			x"0000" when x"35A3",
			x"0000" when x"35A4",
			x"0000" when x"35A5",
			x"0000" when x"35A6",
			x"0000" when x"35A7",
			x"0000" when x"35A8",
			x"0000" when x"35A9",
			x"0000" when x"35AA",
			x"0000" when x"35AB",
			x"0000" when x"35AC",
			x"0000" when x"35AD",
			x"0000" when x"35AE",
			x"0000" when x"35AF",
			x"0000" when x"35B0",
			x"0000" when x"35B1",
			x"0000" when x"35B2",
			x"0000" when x"35B3",
			x"0000" when x"35B4",
			x"0000" when x"35B5",
			x"0000" when x"35B6",
			x"0000" when x"35B7",
			x"0000" when x"35B8",
			x"0000" when x"35B9",
			x"0000" when x"35BA",
			x"0000" when x"35BB",
			x"0000" when x"35BC",
			x"0000" when x"35BD",
			x"0000" when x"35BE",
			x"0000" when x"35BF",
			x"0000" when x"35C0",
			x"0000" when x"35C1",
			x"0000" when x"35C2",
			x"0000" when x"35C3",
			x"0000" when x"35C4",
			x"0000" when x"35C5",
			x"0000" when x"35C6",
			x"0000" when x"35C7",
			x"0000" when x"35C8",
			x"0000" when x"35C9",
			x"0000" when x"35CA",
			x"0000" when x"35CB",
			x"0000" when x"35CC",
			x"0000" when x"35CD",
			x"0000" when x"35CE",
			x"0000" when x"35CF",
			x"0000" when x"35D0",
			x"0000" when x"35D1",
			x"0000" when x"35D2",
			x"0000" when x"35D3",
			x"0000" when x"35D4",
			x"0000" when x"35D5",
			x"0000" when x"35D6",
			x"0000" when x"35D7",
			x"0000" when x"35D8",
			x"0000" when x"35D9",
			x"0000" when x"35DA",
			x"0000" when x"35DB",
			x"0000" when x"35DC",
			x"0000" when x"35DD",
			x"0000" when x"35DE",
			x"0000" when x"35DF",
			x"0000" when x"35E0",
			x"0000" when x"35E1",
			x"0000" when x"35E2",
			x"0000" when x"35E3",
			x"0000" when x"35E4",
			x"0000" when x"35E5",
			x"0000" when x"35E6",
			x"0000" when x"35E7",
			x"0000" when x"35E8",
			x"0000" when x"35E9",
			x"0000" when x"35EA",
			x"0000" when x"35EB",
			x"0000" when x"35EC",
			x"0000" when x"35ED",
			x"0000" when x"35EE",
			x"0000" when x"35EF",
			x"0000" when x"35F0",
			x"0000" when x"35F1",
			x"0000" when x"35F2",
			x"0000" when x"35F3",
			x"0000" when x"35F4",
			x"0000" when x"35F5",
			x"0000" when x"35F6",
			x"0000" when x"35F7",
			x"0000" when x"35F8",
			x"0000" when x"35F9",
			x"0000" when x"35FA",
			x"0000" when x"35FB",
			x"0000" when x"35FC",
			x"0000" when x"35FD",
			x"0000" when x"35FE",
			x"0000" when x"35FF",
			x"0000" when x"3600",
			x"0000" when x"3601",
			x"0000" when x"3602",
			x"0000" when x"3603",
			x"0000" when x"3604",
			x"0000" when x"3605",
			x"0000" when x"3606",
			x"0000" when x"3607",
			x"0000" when x"3608",
			x"0000" when x"3609",
			x"0000" when x"360A",
			x"0000" when x"360B",
			x"0000" when x"360C",
			x"0000" when x"360D",
			x"0000" when x"360E",
			x"0000" when x"360F",
			x"0000" when x"3610",
			x"0000" when x"3611",
			x"0000" when x"3612",
			x"0000" when x"3613",
			x"0000" when x"3614",
			x"0000" when x"3615",
			x"0000" when x"3616",
			x"0000" when x"3617",
			x"0000" when x"3618",
			x"0000" when x"3619",
			x"0000" when x"361A",
			x"0000" when x"361B",
			x"0000" when x"361C",
			x"0000" when x"361D",
			x"0000" when x"361E",
			x"0000" when x"361F",
			x"0000" when x"3620",
			x"0000" when x"3621",
			x"0000" when x"3622",
			x"0000" when x"3623",
			x"0000" when x"3624",
			x"0000" when x"3625",
			x"0000" when x"3626",
			x"0000" when x"3627",
			x"0000" when x"3628",
			x"0000" when x"3629",
			x"0000" when x"362A",
			x"0000" when x"362B",
			x"0000" when x"362C",
			x"0000" when x"362D",
			x"0000" when x"362E",
			x"0000" when x"362F",
			x"0000" when x"3630",
			x"0000" when x"3631",
			x"0000" when x"3632",
			x"0000" when x"3633",
			x"0000" when x"3634",
			x"0000" when x"3635",
			x"0000" when x"3636",
			x"0000" when x"3637",
			x"0000" when x"3638",
			x"0000" when x"3639",
			x"0000" when x"363A",
			x"0000" when x"363B",
			x"0000" when x"363C",
			x"0000" when x"363D",
			x"0000" when x"363E",
			x"0000" when x"363F",
			x"0000" when x"3640",
			x"0000" when x"3641",
			x"0000" when x"3642",
			x"0000" when x"3643",
			x"0000" when x"3644",
			x"0000" when x"3645",
			x"0000" when x"3646",
			x"0000" when x"3647",
			x"0000" when x"3648",
			x"0000" when x"3649",
			x"0000" when x"364A",
			x"0000" when x"364B",
			x"0000" when x"364C",
			x"0000" when x"364D",
			x"0000" when x"364E",
			x"0000" when x"364F",
			x"0000" when x"3650",
			x"0000" when x"3651",
			x"0000" when x"3652",
			x"0000" when x"3653",
			x"0000" when x"3654",
			x"0000" when x"3655",
			x"0000" when x"3656",
			x"0000" when x"3657",
			x"0000" when x"3658",
			x"0000" when x"3659",
			x"0000" when x"365A",
			x"0000" when x"365B",
			x"0000" when x"365C",
			x"0000" when x"365D",
			x"0000" when x"365E",
			x"0000" when x"365F",
			x"0000" when x"3660",
			x"0000" when x"3661",
			x"0000" when x"3662",
			x"0000" when x"3663",
			x"0000" when x"3664",
			x"0000" when x"3665",
			x"0000" when x"3666",
			x"0000" when x"3667",
			x"0000" when x"3668",
			x"0000" when x"3669",
			x"0000" when x"366A",
			x"0000" when x"366B",
			x"0000" when x"366C",
			x"0000" when x"366D",
			x"0000" when x"366E",
			x"0000" when x"366F",
			x"0000" when x"3670",
			x"0000" when x"3671",
			x"0000" when x"3672",
			x"0000" when x"3673",
			x"0000" when x"3674",
			x"0000" when x"3675",
			x"0000" when x"3676",
			x"0000" when x"3677",
			x"0000" when x"3678",
			x"0000" when x"3679",
			x"0000" when x"367A",
			x"0000" when x"367B",
			x"0000" when x"367C",
			x"0000" when x"367D",
			x"0000" when x"367E",
			x"0000" when x"367F",
			x"0000" when x"3680",
			x"0000" when x"3681",
			x"0000" when x"3682",
			x"0000" when x"3683",
			x"0000" when x"3684",
			x"0000" when x"3685",
			x"0000" when x"3686",
			x"0000" when x"3687",
			x"0000" when x"3688",
			x"0000" when x"3689",
			x"0000" when x"368A",
			x"0000" when x"368B",
			x"0000" when x"368C",
			x"0000" when x"368D",
			x"0000" when x"368E",
			x"0000" when x"368F",
			x"0000" when x"3690",
			x"0000" when x"3691",
			x"0000" when x"3692",
			x"0000" when x"3693",
			x"0000" when x"3694",
			x"0000" when x"3695",
			x"0000" when x"3696",
			x"0000" when x"3697",
			x"0000" when x"3698",
			x"0000" when x"3699",
			x"0000" when x"369A",
			x"0000" when x"369B",
			x"0000" when x"369C",
			x"0000" when x"369D",
			x"0000" when x"369E",
			x"0000" when x"369F",
			x"0000" when x"36A0",
			x"0000" when x"36A1",
			x"0000" when x"36A2",
			x"0000" when x"36A3",
			x"0000" when x"36A4",
			x"0000" when x"36A5",
			x"0000" when x"36A6",
			x"0000" when x"36A7",
			x"0000" when x"36A8",
			x"0000" when x"36A9",
			x"0000" when x"36AA",
			x"0000" when x"36AB",
			x"0000" when x"36AC",
			x"0000" when x"36AD",
			x"0000" when x"36AE",
			x"0000" when x"36AF",
			x"0000" when x"36B0",
			x"0000" when x"36B1",
			x"0000" when x"36B2",
			x"0000" when x"36B3",
			x"0000" when x"36B4",
			x"0000" when x"36B5",
			x"0000" when x"36B6",
			x"0000" when x"36B7",
			x"0000" when x"36B8",
			x"0000" when x"36B9",
			x"0000" when x"36BA",
			x"0000" when x"36BB",
			x"0000" when x"36BC",
			x"0000" when x"36BD",
			x"0000" when x"36BE",
			x"0000" when x"36BF",
			x"0000" when x"36C0",
			x"0000" when x"36C1",
			x"0000" when x"36C2",
			x"0000" when x"36C3",
			x"0000" when x"36C4",
			x"0000" when x"36C5",
			x"0000" when x"36C6",
			x"0000" when x"36C7",
			x"0000" when x"36C8",
			x"0000" when x"36C9",
			x"0000" when x"36CA",
			x"0000" when x"36CB",
			x"0000" when x"36CC",
			x"0000" when x"36CD",
			x"0000" when x"36CE",
			x"0000" when x"36CF",
			x"0000" when x"36D0",
			x"0000" when x"36D1",
			x"0000" when x"36D2",
			x"0000" when x"36D3",
			x"0000" when x"36D4",
			x"0000" when x"36D5",
			x"0000" when x"36D6",
			x"0000" when x"36D7",
			x"0000" when x"36D8",
			x"0000" when x"36D9",
			x"0000" when x"36DA",
			x"0000" when x"36DB",
			x"0000" when x"36DC",
			x"0000" when x"36DD",
			x"0000" when x"36DE",
			x"0000" when x"36DF",
			x"0000" when x"36E0",
			x"0000" when x"36E1",
			x"0000" when x"36E2",
			x"0000" when x"36E3",
			x"0000" when x"36E4",
			x"0000" when x"36E5",
			x"0000" when x"36E6",
			x"0000" when x"36E7",
			x"0000" when x"36E8",
			x"0000" when x"36E9",
			x"0000" when x"36EA",
			x"0000" when x"36EB",
			x"0000" when x"36EC",
			x"0000" when x"36ED",
			x"0000" when x"36EE",
			x"0000" when x"36EF",
			x"0000" when x"36F0",
			x"0000" when x"36F1",
			x"0000" when x"36F2",
			x"0000" when x"36F3",
			x"0000" when x"36F4",
			x"0000" when x"36F5",
			x"0000" when x"36F6",
			x"0000" when x"36F7",
			x"0000" when x"36F8",
			x"0000" when x"36F9",
			x"0000" when x"36FA",
			x"0000" when x"36FB",
			x"0000" when x"36FC",
			x"0000" when x"36FD",
			x"0000" when x"36FE",
			x"0000" when x"36FF",
			x"0000" when x"3700",
			x"0000" when x"3701",
			x"0000" when x"3702",
			x"0000" when x"3703",
			x"0000" when x"3704",
			x"0000" when x"3705",
			x"0000" when x"3706",
			x"0000" when x"3707",
			x"0000" when x"3708",
			x"0000" when x"3709",
			x"0000" when x"370A",
			x"0000" when x"370B",
			x"0000" when x"370C",
			x"0000" when x"370D",
			x"0000" when x"370E",
			x"0000" when x"370F",
			x"0000" when x"3710",
			x"0000" when x"3711",
			x"0000" when x"3712",
			x"0000" when x"3713",
			x"0000" when x"3714",
			x"0000" when x"3715",
			x"0000" when x"3716",
			x"0000" when x"3717",
			x"0000" when x"3718",
			x"0000" when x"3719",
			x"0000" when x"371A",
			x"0000" when x"371B",
			x"0000" when x"371C",
			x"0000" when x"371D",
			x"0000" when x"371E",
			x"0000" when x"371F",
			x"0000" when x"3720",
			x"0000" when x"3721",
			x"0000" when x"3722",
			x"0000" when x"3723",
			x"0000" when x"3724",
			x"0000" when x"3725",
			x"0000" when x"3726",
			x"0000" when x"3727",
			x"0000" when x"3728",
			x"0000" when x"3729",
			x"0000" when x"372A",
			x"0000" when x"372B",
			x"0000" when x"372C",
			x"0000" when x"372D",
			x"0000" when x"372E",
			x"0000" when x"372F",
			x"0000" when x"3730",
			x"0000" when x"3731",
			x"0000" when x"3732",
			x"0000" when x"3733",
			x"0000" when x"3734",
			x"0000" when x"3735",
			x"0000" when x"3736",
			x"0000" when x"3737",
			x"0000" when x"3738",
			x"0000" when x"3739",
			x"0000" when x"373A",
			x"0000" when x"373B",
			x"0000" when x"373C",
			x"0000" when x"373D",
			x"0000" when x"373E",
			x"0000" when x"373F",
			x"0000" when x"3740",
			x"0000" when x"3741",
			x"0000" when x"3742",
			x"0000" when x"3743",
			x"0000" when x"3744",
			x"0000" when x"3745",
			x"0000" when x"3746",
			x"0000" when x"3747",
			x"0000" when x"3748",
			x"0000" when x"3749",
			x"0000" when x"374A",
			x"0000" when x"374B",
			x"0000" when x"374C",
			x"0000" when x"374D",
			x"0000" when x"374E",
			x"0000" when x"374F",
			x"0000" when x"3750",
			x"0000" when x"3751",
			x"0000" when x"3752",
			x"0000" when x"3753",
			x"0000" when x"3754",
			x"0000" when x"3755",
			x"0000" when x"3756",
			x"0000" when x"3757",
			x"0000" when x"3758",
			x"0000" when x"3759",
			x"0000" when x"375A",
			x"0000" when x"375B",
			x"0000" when x"375C",
			x"0000" when x"375D",
			x"0000" when x"375E",
			x"0000" when x"375F",
			x"0000" when x"3760",
			x"0000" when x"3761",
			x"0000" when x"3762",
			x"0000" when x"3763",
			x"0000" when x"3764",
			x"0000" when x"3765",
			x"0000" when x"3766",
			x"0000" when x"3767",
			x"0000" when x"3768",
			x"0000" when x"3769",
			x"0000" when x"376A",
			x"0000" when x"376B",
			x"0000" when x"376C",
			x"0000" when x"376D",
			x"0000" when x"376E",
			x"0000" when x"376F",
			x"0000" when x"3770",
			x"0000" when x"3771",
			x"0000" when x"3772",
			x"0000" when x"3773",
			x"0000" when x"3774",
			x"0000" when x"3775",
			x"0000" when x"3776",
			x"0000" when x"3777",
			x"0000" when x"3778",
			x"0000" when x"3779",
			x"0000" when x"377A",
			x"0000" when x"377B",
			x"0000" when x"377C",
			x"0000" when x"377D",
			x"0000" when x"377E",
			x"0000" when x"377F",
			x"0000" when x"3780",
			x"0000" when x"3781",
			x"0000" when x"3782",
			x"0000" when x"3783",
			x"0000" when x"3784",
			x"0000" when x"3785",
			x"0000" when x"3786",
			x"0000" when x"3787",
			x"0000" when x"3788",
			x"0000" when x"3789",
			x"0000" when x"378A",
			x"0000" when x"378B",
			x"0000" when x"378C",
			x"0000" when x"378D",
			x"0000" when x"378E",
			x"0000" when x"378F",
			x"0000" when x"3790",
			x"0000" when x"3791",
			x"0000" when x"3792",
			x"0000" when x"3793",
			x"0000" when x"3794",
			x"0000" when x"3795",
			x"0000" when x"3796",
			x"0000" when x"3797",
			x"0000" when x"3798",
			x"0000" when x"3799",
			x"0000" when x"379A",
			x"0000" when x"379B",
			x"0000" when x"379C",
			x"0000" when x"379D",
			x"0000" when x"379E",
			x"0000" when x"379F",
			x"0000" when x"37A0",
			x"0000" when x"37A1",
			x"0000" when x"37A2",
			x"0000" when x"37A3",
			x"0000" when x"37A4",
			x"0000" when x"37A5",
			x"0000" when x"37A6",
			x"0000" when x"37A7",
			x"0000" when x"37A8",
			x"0000" when x"37A9",
			x"0000" when x"37AA",
			x"0000" when x"37AB",
			x"0000" when x"37AC",
			x"0000" when x"37AD",
			x"0000" when x"37AE",
			x"0000" when x"37AF",
			x"0000" when x"37B0",
			x"0000" when x"37B1",
			x"0000" when x"37B2",
			x"0000" when x"37B3",
			x"0000" when x"37B4",
			x"0000" when x"37B5",
			x"0000" when x"37B6",
			x"0000" when x"37B7",
			x"0000" when x"37B8",
			x"0000" when x"37B9",
			x"0000" when x"37BA",
			x"0000" when x"37BB",
			x"0000" when x"37BC",
			x"0000" when x"37BD",
			x"0000" when x"37BE",
			x"0000" when x"37BF",
			x"0000" when x"37C0",
			x"0000" when x"37C1",
			x"0000" when x"37C2",
			x"0000" when x"37C3",
			x"0000" when x"37C4",
			x"0000" when x"37C5",
			x"0000" when x"37C6",
			x"0000" when x"37C7",
			x"0000" when x"37C8",
			x"0000" when x"37C9",
			x"0000" when x"37CA",
			x"0000" when x"37CB",
			x"0000" when x"37CC",
			x"0000" when x"37CD",
			x"0000" when x"37CE",
			x"0000" when x"37CF",
			x"0000" when x"37D0",
			x"0000" when x"37D1",
			x"0000" when x"37D2",
			x"0000" when x"37D3",
			x"0000" when x"37D4",
			x"0000" when x"37D5",
			x"0000" when x"37D6",
			x"0000" when x"37D7",
			x"0000" when x"37D8",
			x"0000" when x"37D9",
			x"0000" when x"37DA",
			x"0000" when x"37DB",
			x"0000" when x"37DC",
			x"0000" when x"37DD",
			x"0000" when x"37DE",
			x"0000" when x"37DF",
			x"0000" when x"37E0",
			x"0000" when x"37E1",
			x"0000" when x"37E2",
			x"0000" when x"37E3",
			x"0000" when x"37E4",
			x"0000" when x"37E5",
			x"0000" when x"37E6",
			x"0000" when x"37E7",
			x"0000" when x"37E8",
			x"0000" when x"37E9",
			x"0000" when x"37EA",
			x"0000" when x"37EB",
			x"0000" when x"37EC",
			x"0000" when x"37ED",
			x"0000" when x"37EE",
			x"0000" when x"37EF",
			x"0000" when x"37F0",
			x"0000" when x"37F1",
			x"0000" when x"37F2",
			x"0000" when x"37F3",
			x"0000" when x"37F4",
			x"0000" when x"37F5",
			x"0000" when x"37F6",
			x"0000" when x"37F7",
			x"0000" when x"37F8",
			x"0000" when x"37F9",
			x"0000" when x"37FA",
			x"0000" when x"37FB",
			x"0000" when x"37FC",
			x"0000" when x"37FD",
			x"0000" when x"37FE",
			x"0000" when x"37FF",
			x"0000" when x"3800",
			x"0000" when x"3801",
			x"0000" when x"3802",
			x"0000" when x"3803",
			x"0000" when x"3804",
			x"0000" when x"3805",
			x"0000" when x"3806",
			x"0000" when x"3807",
			x"0000" when x"3808",
			x"0000" when x"3809",
			x"0000" when x"380A",
			x"0000" when x"380B",
			x"0000" when x"380C",
			x"0000" when x"380D",
			x"0000" when x"380E",
			x"0000" when x"380F",
			x"0000" when x"3810",
			x"0000" when x"3811",
			x"0000" when x"3812",
			x"0000" when x"3813",
			x"0000" when x"3814",
			x"0000" when x"3815",
			x"0000" when x"3816",
			x"0000" when x"3817",
			x"0000" when x"3818",
			x"0000" when x"3819",
			x"0000" when x"381A",
			x"0000" when x"381B",
			x"0000" when x"381C",
			x"0000" when x"381D",
			x"0000" when x"381E",
			x"0000" when x"381F",
			x"0000" when x"3820",
			x"0000" when x"3821",
			x"0000" when x"3822",
			x"0000" when x"3823",
			x"0000" when x"3824",
			x"0000" when x"3825",
			x"0000" when x"3826",
			x"0000" when x"3827",
			x"0000" when x"3828",
			x"0000" when x"3829",
			x"0000" when x"382A",
			x"0000" when x"382B",
			x"0000" when x"382C",
			x"0000" when x"382D",
			x"0000" when x"382E",
			x"0000" when x"382F",
			x"0000" when x"3830",
			x"0000" when x"3831",
			x"0000" when x"3832",
			x"0000" when x"3833",
			x"0000" when x"3834",
			x"0000" when x"3835",
			x"0000" when x"3836",
			x"0000" when x"3837",
			x"0000" when x"3838",
			x"0000" when x"3839",
			x"0000" when x"383A",
			x"0000" when x"383B",
			x"0000" when x"383C",
			x"0000" when x"383D",
			x"0000" when x"383E",
			x"0000" when x"383F",
			x"0000" when x"3840",
			x"0000" when x"3841",
			x"0000" when x"3842",
			x"0000" when x"3843",
			x"0000" when x"3844",
			x"0000" when x"3845",
			x"0000" when x"3846",
			x"0000" when x"3847",
			x"0000" when x"3848",
			x"0000" when x"3849",
			x"0000" when x"384A",
			x"0000" when x"384B",
			x"0000" when x"384C",
			x"0000" when x"384D",
			x"0000" when x"384E",
			x"0000" when x"384F",
			x"0000" when x"3850",
			x"0000" when x"3851",
			x"0000" when x"3852",
			x"0000" when x"3853",
			x"0000" when x"3854",
			x"0000" when x"3855",
			x"0000" when x"3856",
			x"0000" when x"3857",
			x"0000" when x"3858",
			x"0000" when x"3859",
			x"0000" when x"385A",
			x"0000" when x"385B",
			x"0000" when x"385C",
			x"0000" when x"385D",
			x"0000" when x"385E",
			x"0000" when x"385F",
			x"0000" when x"3860",
			x"0000" when x"3861",
			x"0000" when x"3862",
			x"0000" when x"3863",
			x"0000" when x"3864",
			x"0000" when x"3865",
			x"0000" when x"3866",
			x"0000" when x"3867",
			x"0000" when x"3868",
			x"0000" when x"3869",
			x"0000" when x"386A",
			x"0000" when x"386B",
			x"0000" when x"386C",
			x"0000" when x"386D",
			x"0000" when x"386E",
			x"0000" when x"386F",
			x"0000" when x"3870",
			x"0000" when x"3871",
			x"0000" when x"3872",
			x"0000" when x"3873",
			x"0000" when x"3874",
			x"0000" when x"3875",
			x"0000" when x"3876",
			x"0000" when x"3877",
			x"0000" when x"3878",
			x"0000" when x"3879",
			x"0000" when x"387A",
			x"0000" when x"387B",
			x"0000" when x"387C",
			x"0000" when x"387D",
			x"0000" when x"387E",
			x"0000" when x"387F",
			x"0000" when x"3880",
			x"0000" when x"3881",
			x"0000" when x"3882",
			x"0000" when x"3883",
			x"0000" when x"3884",
			x"0000" when x"3885",
			x"0000" when x"3886",
			x"0000" when x"3887",
			x"0000" when x"3888",
			x"0000" when x"3889",
			x"0000" when x"388A",
			x"0000" when x"388B",
			x"0000" when x"388C",
			x"0000" when x"388D",
			x"0000" when x"388E",
			x"0000" when x"388F",
			x"0000" when x"3890",
			x"0000" when x"3891",
			x"0000" when x"3892",
			x"0000" when x"3893",
			x"0000" when x"3894",
			x"0000" when x"3895",
			x"0000" when x"3896",
			x"0000" when x"3897",
			x"0000" when x"3898",
			x"0000" when x"3899",
			x"0000" when x"389A",
			x"0000" when x"389B",
			x"0000" when x"389C",
			x"0000" when x"389D",
			x"0000" when x"389E",
			x"0000" when x"389F",
			x"0000" when x"38A0",
			x"0000" when x"38A1",
			x"0000" when x"38A2",
			x"0000" when x"38A3",
			x"0000" when x"38A4",
			x"0000" when x"38A5",
			x"0000" when x"38A6",
			x"0000" when x"38A7",
			x"0000" when x"38A8",
			x"0000" when x"38A9",
			x"0000" when x"38AA",
			x"0000" when x"38AB",
			x"0000" when x"38AC",
			x"0000" when x"38AD",
			x"0000" when x"38AE",
			x"0000" when x"38AF",
			x"0000" when x"38B0",
			x"0000" when x"38B1",
			x"0000" when x"38B2",
			x"0000" when x"38B3",
			x"0000" when x"38B4",
			x"0000" when x"38B5",
			x"0000" when x"38B6",
			x"0000" when x"38B7",
			x"0000" when x"38B8",
			x"0000" when x"38B9",
			x"0000" when x"38BA",
			x"0000" when x"38BB",
			x"0000" when x"38BC",
			x"0000" when x"38BD",
			x"0000" when x"38BE",
			x"0000" when x"38BF",
			x"0000" when x"38C0",
			x"0000" when x"38C1",
			x"0000" when x"38C2",
			x"0000" when x"38C3",
			x"0000" when x"38C4",
			x"0000" when x"38C5",
			x"0000" when x"38C6",
			x"0000" when x"38C7",
			x"0000" when x"38C8",
			x"0000" when x"38C9",
			x"0000" when x"38CA",
			x"0000" when x"38CB",
			x"0000" when x"38CC",
			x"0000" when x"38CD",
			x"0000" when x"38CE",
			x"0000" when x"38CF",
			x"0000" when x"38D0",
			x"0000" when x"38D1",
			x"0000" when x"38D2",
			x"0000" when x"38D3",
			x"0000" when x"38D4",
			x"0000" when x"38D5",
			x"0000" when x"38D6",
			x"0000" when x"38D7",
			x"0000" when x"38D8",
			x"0000" when x"38D9",
			x"0000" when x"38DA",
			x"0000" when x"38DB",
			x"0000" when x"38DC",
			x"0000" when x"38DD",
			x"0000" when x"38DE",
			x"0000" when x"38DF",
			x"0000" when x"38E0",
			x"0000" when x"38E1",
			x"0000" when x"38E2",
			x"0000" when x"38E3",
			x"0000" when x"38E4",
			x"0000" when x"38E5",
			x"0000" when x"38E6",
			x"0000" when x"38E7",
			x"0000" when x"38E8",
			x"0000" when x"38E9",
			x"0000" when x"38EA",
			x"0000" when x"38EB",
			x"0000" when x"38EC",
			x"0000" when x"38ED",
			x"0000" when x"38EE",
			x"0000" when x"38EF",
			x"0000" when x"38F0",
			x"0000" when x"38F1",
			x"0000" when x"38F2",
			x"0000" when x"38F3",
			x"0000" when x"38F4",
			x"0000" when x"38F5",
			x"0000" when x"38F6",
			x"0000" when x"38F7",
			x"0000" when x"38F8",
			x"0000" when x"38F9",
			x"0000" when x"38FA",
			x"0000" when x"38FB",
			x"0000" when x"38FC",
			x"0000" when x"38FD",
			x"0000" when x"38FE",
			x"0000" when x"38FF",
			x"0000" when x"3900",
			x"0000" when x"3901",
			x"0000" when x"3902",
			x"0000" when x"3903",
			x"0000" when x"3904",
			x"0000" when x"3905",
			x"0000" when x"3906",
			x"0000" when x"3907",
			x"0000" when x"3908",
			x"0000" when x"3909",
			x"0000" when x"390A",
			x"0000" when x"390B",
			x"0000" when x"390C",
			x"0000" when x"390D",
			x"0000" when x"390E",
			x"0000" when x"390F",
			x"0000" when x"3910",
			x"0000" when x"3911",
			x"0000" when x"3912",
			x"0000" when x"3913",
			x"0000" when x"3914",
			x"0000" when x"3915",
			x"0000" when x"3916",
			x"0000" when x"3917",
			x"0000" when x"3918",
			x"0000" when x"3919",
			x"0000" when x"391A",
			x"0000" when x"391B",
			x"0000" when x"391C",
			x"0000" when x"391D",
			x"0000" when x"391E",
			x"0000" when x"391F",
			x"0000" when x"3920",
			x"0000" when x"3921",
			x"0000" when x"3922",
			x"0000" when x"3923",
			x"0000" when x"3924",
			x"0000" when x"3925",
			x"0000" when x"3926",
			x"0000" when x"3927",
			x"0000" when x"3928",
			x"0000" when x"3929",
			x"0000" when x"392A",
			x"0000" when x"392B",
			x"0000" when x"392C",
			x"0000" when x"392D",
			x"0000" when x"392E",
			x"0000" when x"392F",
			x"0000" when x"3930",
			x"0000" when x"3931",
			x"0000" when x"3932",
			x"0000" when x"3933",
			x"0000" when x"3934",
			x"0000" when x"3935",
			x"0000" when x"3936",
			x"0000" when x"3937",
			x"0000" when x"3938",
			x"0000" when x"3939",
			x"0000" when x"393A",
			x"0000" when x"393B",
			x"0000" when x"393C",
			x"0000" when x"393D",
			x"0000" when x"393E",
			x"0000" when x"393F",
			x"0000" when x"3940",
			x"0000" when x"3941",
			x"0000" when x"3942",
			x"0000" when x"3943",
			x"0000" when x"3944",
			x"0000" when x"3945",
			x"0000" when x"3946",
			x"0000" when x"3947",
			x"0000" when x"3948",
			x"0000" when x"3949",
			x"0000" when x"394A",
			x"0000" when x"394B",
			x"0000" when x"394C",
			x"0000" when x"394D",
			x"0000" when x"394E",
			x"0000" when x"394F",
			x"0000" when x"3950",
			x"0000" when x"3951",
			x"0000" when x"3952",
			x"0000" when x"3953",
			x"0000" when x"3954",
			x"0000" when x"3955",
			x"0000" when x"3956",
			x"0000" when x"3957",
			x"0000" when x"3958",
			x"0000" when x"3959",
			x"0000" when x"395A",
			x"0000" when x"395B",
			x"0000" when x"395C",
			x"0000" when x"395D",
			x"0000" when x"395E",
			x"0000" when x"395F",
			x"0000" when x"3960",
			x"0000" when x"3961",
			x"0000" when x"3962",
			x"0000" when x"3963",
			x"0000" when x"3964",
			x"0000" when x"3965",
			x"0000" when x"3966",
			x"0000" when x"3967",
			x"0000" when x"3968",
			x"0000" when x"3969",
			x"0000" when x"396A",
			x"0000" when x"396B",
			x"0000" when x"396C",
			x"0000" when x"396D",
			x"0000" when x"396E",
			x"0000" when x"396F",
			x"0000" when x"3970",
			x"0000" when x"3971",
			x"0000" when x"3972",
			x"0000" when x"3973",
			x"0000" when x"3974",
			x"0000" when x"3975",
			x"0000" when x"3976",
			x"0000" when x"3977",
			x"0000" when x"3978",
			x"0000" when x"3979",
			x"0000" when x"397A",
			x"0000" when x"397B",
			x"0000" when x"397C",
			x"0000" when x"397D",
			x"0000" when x"397E",
			x"0000" when x"397F",
			x"0000" when x"3980",
			x"0000" when x"3981",
			x"0000" when x"3982",
			x"0000" when x"3983",
			x"0000" when x"3984",
			x"0000" when x"3985",
			x"0000" when x"3986",
			x"0000" when x"3987",
			x"0000" when x"3988",
			x"0000" when x"3989",
			x"0000" when x"398A",
			x"0000" when x"398B",
			x"0000" when x"398C",
			x"0000" when x"398D",
			x"0000" when x"398E",
			x"0000" when x"398F",
			x"0000" when x"3990",
			x"0000" when x"3991",
			x"0000" when x"3992",
			x"0000" when x"3993",
			x"0000" when x"3994",
			x"0000" when x"3995",
			x"0000" when x"3996",
			x"0000" when x"3997",
			x"0000" when x"3998",
			x"0000" when x"3999",
			x"0000" when x"399A",
			x"0000" when x"399B",
			x"0000" when x"399C",
			x"0000" when x"399D",
			x"0000" when x"399E",
			x"0000" when x"399F",
			x"0000" when x"39A0",
			x"0000" when x"39A1",
			x"0000" when x"39A2",
			x"0000" when x"39A3",
			x"0000" when x"39A4",
			x"0000" when x"39A5",
			x"0000" when x"39A6",
			x"0000" when x"39A7",
			x"0000" when x"39A8",
			x"0000" when x"39A9",
			x"0000" when x"39AA",
			x"0000" when x"39AB",
			x"0000" when x"39AC",
			x"0000" when x"39AD",
			x"0000" when x"39AE",
			x"0000" when x"39AF",
			x"0000" when x"39B0",
			x"0000" when x"39B1",
			x"0000" when x"39B2",
			x"0000" when x"39B3",
			x"0000" when x"39B4",
			x"0000" when x"39B5",
			x"0000" when x"39B6",
			x"0000" when x"39B7",
			x"0000" when x"39B8",
			x"0000" when x"39B9",
			x"0000" when x"39BA",
			x"0000" when x"39BB",
			x"0000" when x"39BC",
			x"0000" when x"39BD",
			x"0000" when x"39BE",
			x"0000" when x"39BF",
			x"0000" when x"39C0",
			x"0000" when x"39C1",
			x"0000" when x"39C2",
			x"0000" when x"39C3",
			x"0000" when x"39C4",
			x"0000" when x"39C5",
			x"0000" when x"39C6",
			x"0000" when x"39C7",
			x"0000" when x"39C8",
			x"0000" when x"39C9",
			x"0000" when x"39CA",
			x"0000" when x"39CB",
			x"0000" when x"39CC",
			x"0000" when x"39CD",
			x"0000" when x"39CE",
			x"0000" when x"39CF",
			x"0000" when x"39D0",
			x"0000" when x"39D1",
			x"0000" when x"39D2",
			x"0000" when x"39D3",
			x"0000" when x"39D4",
			x"0000" when x"39D5",
			x"0000" when x"39D6",
			x"0000" when x"39D7",
			x"0000" when x"39D8",
			x"0000" when x"39D9",
			x"0000" when x"39DA",
			x"0000" when x"39DB",
			x"0000" when x"39DC",
			x"0000" when x"39DD",
			x"0000" when x"39DE",
			x"0000" when x"39DF",
			x"0000" when x"39E0",
			x"0000" when x"39E1",
			x"0000" when x"39E2",
			x"0000" when x"39E3",
			x"0000" when x"39E4",
			x"0000" when x"39E5",
			x"0000" when x"39E6",
			x"0000" when x"39E7",
			x"0000" when x"39E8",
			x"0000" when x"39E9",
			x"0000" when x"39EA",
			x"0000" when x"39EB",
			x"0000" when x"39EC",
			x"0000" when x"39ED",
			x"0000" when x"39EE",
			x"0000" when x"39EF",
			x"0000" when x"39F0",
			x"0000" when x"39F1",
			x"0000" when x"39F2",
			x"0000" when x"39F3",
			x"0000" when x"39F4",
			x"0000" when x"39F5",
			x"0000" when x"39F6",
			x"0000" when x"39F7",
			x"0000" when x"39F8",
			x"0000" when x"39F9",
			x"0000" when x"39FA",
			x"0000" when x"39FB",
			x"0000" when x"39FC",
			x"0000" when x"39FD",
			x"0000" when x"39FE",
			x"0000" when x"39FF",
			x"0000" when x"3A00",
			x"0000" when x"3A01",
			x"0000" when x"3A02",
			x"0000" when x"3A03",
			x"0000" when x"3A04",
			x"0000" when x"3A05",
			x"0000" when x"3A06",
			x"0000" when x"3A07",
			x"0000" when x"3A08",
			x"0000" when x"3A09",
			x"0000" when x"3A0A",
			x"0000" when x"3A0B",
			x"0000" when x"3A0C",
			x"0000" when x"3A0D",
			x"0000" when x"3A0E",
			x"0000" when x"3A0F",
			x"0000" when x"3A10",
			x"0000" when x"3A11",
			x"0000" when x"3A12",
			x"0000" when x"3A13",
			x"0000" when x"3A14",
			x"0000" when x"3A15",
			x"0000" when x"3A16",
			x"0000" when x"3A17",
			x"0000" when x"3A18",
			x"0000" when x"3A19",
			x"0000" when x"3A1A",
			x"0000" when x"3A1B",
			x"0000" when x"3A1C",
			x"0000" when x"3A1D",
			x"0000" when x"3A1E",
			x"0000" when x"3A1F",
			x"0000" when x"3A20",
			x"0000" when x"3A21",
			x"0000" when x"3A22",
			x"0000" when x"3A23",
			x"0000" when x"3A24",
			x"0000" when x"3A25",
			x"0000" when x"3A26",
			x"0000" when x"3A27",
			x"0000" when x"3A28",
			x"0000" when x"3A29",
			x"0000" when x"3A2A",
			x"0000" when x"3A2B",
			x"0000" when x"3A2C",
			x"0000" when x"3A2D",
			x"0000" when x"3A2E",
			x"0000" when x"3A2F",
			x"0000" when x"3A30",
			x"0000" when x"3A31",
			x"0000" when x"3A32",
			x"0000" when x"3A33",
			x"0000" when x"3A34",
			x"0000" when x"3A35",
			x"0000" when x"3A36",
			x"0000" when x"3A37",
			x"0000" when x"3A38",
			x"0000" when x"3A39",
			x"0000" when x"3A3A",
			x"0000" when x"3A3B",
			x"0000" when x"3A3C",
			x"0000" when x"3A3D",
			x"0000" when x"3A3E",
			x"0000" when x"3A3F",
			x"0000" when x"3A40",
			x"0000" when x"3A41",
			x"0000" when x"3A42",
			x"0000" when x"3A43",
			x"0000" when x"3A44",
			x"0000" when x"3A45",
			x"0000" when x"3A46",
			x"0000" when x"3A47",
			x"0000" when x"3A48",
			x"0000" when x"3A49",
			x"0000" when x"3A4A",
			x"0000" when x"3A4B",
			x"0000" when x"3A4C",
			x"0000" when x"3A4D",
			x"0000" when x"3A4E",
			x"0000" when x"3A4F",
			x"0000" when x"3A50",
			x"0000" when x"3A51",
			x"0000" when x"3A52",
			x"0000" when x"3A53",
			x"0000" when x"3A54",
			x"0000" when x"3A55",
			x"0000" when x"3A56",
			x"0000" when x"3A57",
			x"0000" when x"3A58",
			x"0000" when x"3A59",
			x"0000" when x"3A5A",
			x"0000" when x"3A5B",
			x"0000" when x"3A5C",
			x"0000" when x"3A5D",
			x"0000" when x"3A5E",
			x"0000" when x"3A5F",
			x"0000" when x"3A60",
			x"0000" when x"3A61",
			x"0000" when x"3A62",
			x"0000" when x"3A63",
			x"0000" when x"3A64",
			x"0000" when x"3A65",
			x"0000" when x"3A66",
			x"0000" when x"3A67",
			x"0000" when x"3A68",
			x"0000" when x"3A69",
			x"0000" when x"3A6A",
			x"0000" when x"3A6B",
			x"0000" when x"3A6C",
			x"0000" when x"3A6D",
			x"0000" when x"3A6E",
			x"0000" when x"3A6F",
			x"0000" when x"3A70",
			x"0000" when x"3A71",
			x"0000" when x"3A72",
			x"0000" when x"3A73",
			x"0000" when x"3A74",
			x"0000" when x"3A75",
			x"0000" when x"3A76",
			x"0000" when x"3A77",
			x"0000" when x"3A78",
			x"0000" when x"3A79",
			x"0000" when x"3A7A",
			x"0000" when x"3A7B",
			x"0000" when x"3A7C",
			x"0000" when x"3A7D",
			x"0000" when x"3A7E",
			x"0000" when x"3A7F",
			x"0000" when x"3A80",
			x"0000" when x"3A81",
			x"0000" when x"3A82",
			x"0000" when x"3A83",
			x"0000" when x"3A84",
			x"0000" when x"3A85",
			x"0000" when x"3A86",
			x"0000" when x"3A87",
			x"0000" when x"3A88",
			x"0000" when x"3A89",
			x"0000" when x"3A8A",
			x"0000" when x"3A8B",
			x"0000" when x"3A8C",
			x"0000" when x"3A8D",
			x"0000" when x"3A8E",
			x"0000" when x"3A8F",
			x"0000" when x"3A90",
			x"0000" when x"3A91",
			x"0000" when x"3A92",
			x"0000" when x"3A93",
			x"0000" when x"3A94",
			x"0000" when x"3A95",
			x"0000" when x"3A96",
			x"0000" when x"3A97",
			x"0000" when x"3A98",
			x"0000" when x"3A99",
			x"0000" when x"3A9A",
			x"0000" when x"3A9B",
			x"0000" when x"3A9C",
			x"0000" when x"3A9D",
			x"0000" when x"3A9E",
			x"0000" when x"3A9F",
			x"0000" when x"3AA0",
			x"0000" when x"3AA1",
			x"0000" when x"3AA2",
			x"0000" when x"3AA3",
			x"0000" when x"3AA4",
			x"0000" when x"3AA5",
			x"0000" when x"3AA6",
			x"0000" when x"3AA7",
			x"0000" when x"3AA8",
			x"0000" when x"3AA9",
			x"0000" when x"3AAA",
			x"0000" when x"3AAB",
			x"0000" when x"3AAC",
			x"0000" when x"3AAD",
			x"0000" when x"3AAE",
			x"0000" when x"3AAF",
			x"0000" when x"3AB0",
			x"0000" when x"3AB1",
			x"0000" when x"3AB2",
			x"0000" when x"3AB3",
			x"0000" when x"3AB4",
			x"0000" when x"3AB5",
			x"0000" when x"3AB6",
			x"0000" when x"3AB7",
			x"0000" when x"3AB8",
			x"0000" when x"3AB9",
			x"0000" when x"3ABA",
			x"0000" when x"3ABB",
			x"0000" when x"3ABC",
			x"0000" when x"3ABD",
			x"0000" when x"3ABE",
			x"0000" when x"3ABF",
			x"0000" when x"3AC0",
			x"0000" when x"3AC1",
			x"0000" when x"3AC2",
			x"0000" when x"3AC3",
			x"0000" when x"3AC4",
			x"0000" when x"3AC5",
			x"0000" when x"3AC6",
			x"0000" when x"3AC7",
			x"0000" when x"3AC8",
			x"0000" when x"3AC9",
			x"0000" when x"3ACA",
			x"0000" when x"3ACB",
			x"0000" when x"3ACC",
			x"0000" when x"3ACD",
			x"0000" when x"3ACE",
			x"0000" when x"3ACF",
			x"0000" when x"3AD0",
			x"0000" when x"3AD1",
			x"0000" when x"3AD2",
			x"0000" when x"3AD3",
			x"0000" when x"3AD4",
			x"0000" when x"3AD5",
			x"0000" when x"3AD6",
			x"0000" when x"3AD7",
			x"0000" when x"3AD8",
			x"0000" when x"3AD9",
			x"0000" when x"3ADA",
			x"0000" when x"3ADB",
			x"0000" when x"3ADC",
			x"0000" when x"3ADD",
			x"0000" when x"3ADE",
			x"0000" when x"3ADF",
			x"0000" when x"3AE0",
			x"0000" when x"3AE1",
			x"0000" when x"3AE2",
			x"0000" when x"3AE3",
			x"0000" when x"3AE4",
			x"0000" when x"3AE5",
			x"0000" when x"3AE6",
			x"0000" when x"3AE7",
			x"0000" when x"3AE8",
			x"0000" when x"3AE9",
			x"0000" when x"3AEA",
			x"0000" when x"3AEB",
			x"0000" when x"3AEC",
			x"0000" when x"3AED",
			x"0000" when x"3AEE",
			x"0000" when x"3AEF",
			x"0000" when x"3AF0",
			x"0000" when x"3AF1",
			x"0000" when x"3AF2",
			x"0000" when x"3AF3",
			x"0000" when x"3AF4",
			x"0000" when x"3AF5",
			x"0000" when x"3AF6",
			x"0000" when x"3AF7",
			x"0000" when x"3AF8",
			x"0000" when x"3AF9",
			x"0000" when x"3AFA",
			x"0000" when x"3AFB",
			x"0000" when x"3AFC",
			x"0000" when x"3AFD",
			x"0000" when x"3AFE",
			x"0000" when x"3AFF",
			x"0000" when x"3B00",
			x"0000" when x"3B01",
			x"0000" when x"3B02",
			x"0000" when x"3B03",
			x"0000" when x"3B04",
			x"0000" when x"3B05",
			x"0000" when x"3B06",
			x"0000" when x"3B07",
			x"0000" when x"3B08",
			x"0000" when x"3B09",
			x"0000" when x"3B0A",
			x"0000" when x"3B0B",
			x"0000" when x"3B0C",
			x"0000" when x"3B0D",
			x"0000" when x"3B0E",
			x"0000" when x"3B0F",
			x"0000" when x"3B10",
			x"0000" when x"3B11",
			x"0000" when x"3B12",
			x"0000" when x"3B13",
			x"0000" when x"3B14",
			x"0000" when x"3B15",
			x"0000" when x"3B16",
			x"0000" when x"3B17",
			x"0000" when x"3B18",
			x"0000" when x"3B19",
			x"0000" when x"3B1A",
			x"0000" when x"3B1B",
			x"0000" when x"3B1C",
			x"0000" when x"3B1D",
			x"0000" when x"3B1E",
			x"0000" when x"3B1F",
			x"0000" when x"3B20",
			x"0000" when x"3B21",
			x"0000" when x"3B22",
			x"0000" when x"3B23",
			x"0000" when x"3B24",
			x"0000" when x"3B25",
			x"0000" when x"3B26",
			x"0000" when x"3B27",
			x"0000" when x"3B28",
			x"0000" when x"3B29",
			x"0000" when x"3B2A",
			x"0000" when x"3B2B",
			x"0000" when x"3B2C",
			x"0000" when x"3B2D",
			x"0000" when x"3B2E",
			x"0000" when x"3B2F",
			x"0000" when x"3B30",
			x"0000" when x"3B31",
			x"0000" when x"3B32",
			x"0000" when x"3B33",
			x"0000" when x"3B34",
			x"0000" when x"3B35",
			x"0000" when x"3B36",
			x"0000" when x"3B37",
			x"0000" when x"3B38",
			x"0000" when x"3B39",
			x"0000" when x"3B3A",
			x"0000" when x"3B3B",
			x"0000" when x"3B3C",
			x"0000" when x"3B3D",
			x"0000" when x"3B3E",
			x"0000" when x"3B3F",
			x"0000" when x"3B40",
			x"0000" when x"3B41",
			x"0000" when x"3B42",
			x"0000" when x"3B43",
			x"0000" when x"3B44",
			x"0000" when x"3B45",
			x"0000" when x"3B46",
			x"0000" when x"3B47",
			x"0000" when x"3B48",
			x"0000" when x"3B49",
			x"0000" when x"3B4A",
			x"0000" when x"3B4B",
			x"0000" when x"3B4C",
			x"0000" when x"3B4D",
			x"0000" when x"3B4E",
			x"0000" when x"3B4F",
			x"0000" when x"3B50",
			x"0000" when x"3B51",
			x"0000" when x"3B52",
			x"0000" when x"3B53",
			x"0000" when x"3B54",
			x"0000" when x"3B55",
			x"0000" when x"3B56",
			x"0000" when x"3B57",
			x"0000" when x"3B58",
			x"0000" when x"3B59",
			x"0000" when x"3B5A",
			x"0000" when x"3B5B",
			x"0000" when x"3B5C",
			x"0000" when x"3B5D",
			x"0000" when x"3B5E",
			x"0000" when x"3B5F",
			x"0000" when x"3B60",
			x"0000" when x"3B61",
			x"0000" when x"3B62",
			x"0000" when x"3B63",
			x"0000" when x"3B64",
			x"0000" when x"3B65",
			x"0000" when x"3B66",
			x"0000" when x"3B67",
			x"0000" when x"3B68",
			x"0000" when x"3B69",
			x"0000" when x"3B6A",
			x"0000" when x"3B6B",
			x"0000" when x"3B6C",
			x"0000" when x"3B6D",
			x"0000" when x"3B6E",
			x"0000" when x"3B6F",
			x"0000" when x"3B70",
			x"0000" when x"3B71",
			x"0000" when x"3B72",
			x"0000" when x"3B73",
			x"0000" when x"3B74",
			x"0000" when x"3B75",
			x"0000" when x"3B76",
			x"0000" when x"3B77",
			x"0000" when x"3B78",
			x"0000" when x"3B79",
			x"0000" when x"3B7A",
			x"0000" when x"3B7B",
			x"0000" when x"3B7C",
			x"0000" when x"3B7D",
			x"0000" when x"3B7E",
			x"0000" when x"3B7F",
			x"0000" when x"3B80",
			x"0000" when x"3B81",
			x"0000" when x"3B82",
			x"0000" when x"3B83",
			x"0000" when x"3B84",
			x"0000" when x"3B85",
			x"0000" when x"3B86",
			x"0000" when x"3B87",
			x"0000" when x"3B88",
			x"0000" when x"3B89",
			x"0000" when x"3B8A",
			x"0000" when x"3B8B",
			x"0000" when x"3B8C",
			x"0000" when x"3B8D",
			x"0000" when x"3B8E",
			x"0000" when x"3B8F",
			x"0000" when x"3B90",
			x"0000" when x"3B91",
			x"0000" when x"3B92",
			x"0000" when x"3B93",
			x"0000" when x"3B94",
			x"0000" when x"3B95",
			x"0000" when x"3B96",
			x"0000" when x"3B97",
			x"0000" when x"3B98",
			x"0000" when x"3B99",
			x"0000" when x"3B9A",
			x"0000" when x"3B9B",
			x"0000" when x"3B9C",
			x"0000" when x"3B9D",
			x"0000" when x"3B9E",
			x"0000" when x"3B9F",
			x"0000" when x"3BA0",
			x"0000" when x"3BA1",
			x"0000" when x"3BA2",
			x"0000" when x"3BA3",
			x"0000" when x"3BA4",
			x"0000" when x"3BA5",
			x"0000" when x"3BA6",
			x"0000" when x"3BA7",
			x"0000" when x"3BA8",
			x"0000" when x"3BA9",
			x"0000" when x"3BAA",
			x"0000" when x"3BAB",
			x"0000" when x"3BAC",
			x"0000" when x"3BAD",
			x"0000" when x"3BAE",
			x"0000" when x"3BAF",
			x"0000" when x"3BB0",
			x"0000" when x"3BB1",
			x"0000" when x"3BB2",
			x"0000" when x"3BB3",
			x"0000" when x"3BB4",
			x"0000" when x"3BB5",
			x"0000" when x"3BB6",
			x"0000" when x"3BB7",
			x"0000" when x"3BB8",
			x"0000" when x"3BB9",
			x"0000" when x"3BBA",
			x"0000" when x"3BBB",
			x"0000" when x"3BBC",
			x"0000" when x"3BBD",
			x"0000" when x"3BBE",
			x"0000" when x"3BBF",
			x"0000" when x"3BC0",
			x"0000" when x"3BC1",
			x"0000" when x"3BC2",
			x"0000" when x"3BC3",
			x"0000" when x"3BC4",
			x"0000" when x"3BC5",
			x"0000" when x"3BC6",
			x"0000" when x"3BC7",
			x"0000" when x"3BC8",
			x"0000" when x"3BC9",
			x"0000" when x"3BCA",
			x"0000" when x"3BCB",
			x"0000" when x"3BCC",
			x"0000" when x"3BCD",
			x"0000" when x"3BCE",
			x"0000" when x"3BCF",
			x"0000" when x"3BD0",
			x"0000" when x"3BD1",
			x"0000" when x"3BD2",
			x"0000" when x"3BD3",
			x"0000" when x"3BD4",
			x"0000" when x"3BD5",
			x"0000" when x"3BD6",
			x"0000" when x"3BD7",
			x"0000" when x"3BD8",
			x"0000" when x"3BD9",
			x"0000" when x"3BDA",
			x"0000" when x"3BDB",
			x"0000" when x"3BDC",
			x"0000" when x"3BDD",
			x"0000" when x"3BDE",
			x"0000" when x"3BDF",
			x"0000" when x"3BE0",
			x"0000" when x"3BE1",
			x"0000" when x"3BE2",
			x"0000" when x"3BE3",
			x"0000" when x"3BE4",
			x"0000" when x"3BE5",
			x"0000" when x"3BE6",
			x"0000" when x"3BE7",
			x"0000" when x"3BE8",
			x"0000" when x"3BE9",
			x"0000" when x"3BEA",
			x"0000" when x"3BEB",
			x"0000" when x"3BEC",
			x"0000" when x"3BED",
			x"0000" when x"3BEE",
			x"0000" when x"3BEF",
			x"0000" when x"3BF0",
			x"0000" when x"3BF1",
			x"0000" when x"3BF2",
			x"0000" when x"3BF3",
			x"0000" when x"3BF4",
			x"0000" when x"3BF5",
			x"0000" when x"3BF6",
			x"0000" when x"3BF7",
			x"0000" when x"3BF8",
			x"0000" when x"3BF9",
			x"0000" when x"3BFA",
			x"0000" when x"3BFB",
			x"0000" when x"3BFC",
			x"0000" when x"3BFD",
			x"0000" when x"3BFE",
			x"0000" when x"3BFF",
			x"0000" when x"3C00",
			x"0000" when x"3C01",
			x"0000" when x"3C02",
			x"0000" when x"3C03",
			x"0000" when x"3C04",
			x"0000" when x"3C05",
			x"0000" when x"3C06",
			x"0000" when x"3C07",
			x"0000" when x"3C08",
			x"0000" when x"3C09",
			x"0000" when x"3C0A",
			x"0000" when x"3C0B",
			x"0000" when x"3C0C",
			x"0000" when x"3C0D",
			x"0000" when x"3C0E",
			x"0000" when x"3C0F",
			x"0000" when x"3C10",
			x"0000" when x"3C11",
			x"0000" when x"3C12",
			x"0000" when x"3C13",
			x"0000" when x"3C14",
			x"0000" when x"3C15",
			x"0000" when x"3C16",
			x"0000" when x"3C17",
			x"0000" when x"3C18",
			x"0000" when x"3C19",
			x"0000" when x"3C1A",
			x"0000" when x"3C1B",
			x"0000" when x"3C1C",
			x"0000" when x"3C1D",
			x"0000" when x"3C1E",
			x"0000" when x"3C1F",
			x"0000" when x"3C20",
			x"0000" when x"3C21",
			x"0000" when x"3C22",
			x"0000" when x"3C23",
			x"0000" when x"3C24",
			x"0000" when x"3C25",
			x"0000" when x"3C26",
			x"0000" when x"3C27",
			x"0000" when x"3C28",
			x"0000" when x"3C29",
			x"0000" when x"3C2A",
			x"0000" when x"3C2B",
			x"0000" when x"3C2C",
			x"0000" when x"3C2D",
			x"0000" when x"3C2E",
			x"0000" when x"3C2F",
			x"0000" when x"3C30",
			x"0000" when x"3C31",
			x"0000" when x"3C32",
			x"0000" when x"3C33",
			x"0000" when x"3C34",
			x"0000" when x"3C35",
			x"0000" when x"3C36",
			x"0000" when x"3C37",
			x"0000" when x"3C38",
			x"0000" when x"3C39",
			x"0000" when x"3C3A",
			x"0000" when x"3C3B",
			x"0000" when x"3C3C",
			x"0000" when x"3C3D",
			x"0000" when x"3C3E",
			x"0000" when x"3C3F",
			x"0000" when x"3C40",
			x"0000" when x"3C41",
			x"0000" when x"3C42",
			x"0000" when x"3C43",
			x"0000" when x"3C44",
			x"0000" when x"3C45",
			x"0000" when x"3C46",
			x"0000" when x"3C47",
			x"0000" when x"3C48",
			x"0000" when x"3C49",
			x"0000" when x"3C4A",
			x"0000" when x"3C4B",
			x"0000" when x"3C4C",
			x"0000" when x"3C4D",
			x"0000" when x"3C4E",
			x"0000" when x"3C4F",
			x"0000" when x"3C50",
			x"0000" when x"3C51",
			x"0000" when x"3C52",
			x"0000" when x"3C53",
			x"0000" when x"3C54",
			x"0000" when x"3C55",
			x"0000" when x"3C56",
			x"0000" when x"3C57",
			x"0000" when x"3C58",
			x"0000" when x"3C59",
			x"0000" when x"3C5A",
			x"0000" when x"3C5B",
			x"0000" when x"3C5C",
			x"0000" when x"3C5D",
			x"0000" when x"3C5E",
			x"0000" when x"3C5F",
			x"0000" when x"3C60",
			x"0000" when x"3C61",
			x"0000" when x"3C62",
			x"0000" when x"3C63",
			x"0000" when x"3C64",
			x"0000" when x"3C65",
			x"0000" when x"3C66",
			x"0000" when x"3C67",
			x"0000" when x"3C68",
			x"0000" when x"3C69",
			x"0000" when x"3C6A",
			x"0000" when x"3C6B",
			x"0000" when x"3C6C",
			x"0000" when x"3C6D",
			x"0000" when x"3C6E",
			x"0000" when x"3C6F",
			x"0000" when x"3C70",
			x"0000" when x"3C71",
			x"0000" when x"3C72",
			x"0000" when x"3C73",
			x"0000" when x"3C74",
			x"0000" when x"3C75",
			x"0000" when x"3C76",
			x"0000" when x"3C77",
			x"0000" when x"3C78",
			x"0000" when x"3C79",
			x"0000" when x"3C7A",
			x"0000" when x"3C7B",
			x"0000" when x"3C7C",
			x"0000" when x"3C7D",
			x"0000" when x"3C7E",
			x"0000" when x"3C7F",
			x"0000" when x"3C80",
			x"0000" when x"3C81",
			x"0000" when x"3C82",
			x"0000" when x"3C83",
			x"0000" when x"3C84",
			x"0000" when x"3C85",
			x"0000" when x"3C86",
			x"0000" when x"3C87",
			x"0000" when x"3C88",
			x"0000" when x"3C89",
			x"0000" when x"3C8A",
			x"0000" when x"3C8B",
			x"0000" when x"3C8C",
			x"0000" when x"3C8D",
			x"0000" when x"3C8E",
			x"0000" when x"3C8F",
			x"0000" when x"3C90",
			x"0000" when x"3C91",
			x"0000" when x"3C92",
			x"0000" when x"3C93",
			x"0000" when x"3C94",
			x"0000" when x"3C95",
			x"0000" when x"3C96",
			x"0000" when x"3C97",
			x"0000" when x"3C98",
			x"0000" when x"3C99",
			x"0000" when x"3C9A",
			x"0000" when x"3C9B",
			x"0000" when x"3C9C",
			x"0000" when x"3C9D",
			x"0000" when x"3C9E",
			x"0000" when x"3C9F",
			x"0000" when x"3CA0",
			x"0000" when x"3CA1",
			x"0000" when x"3CA2",
			x"0000" when x"3CA3",
			x"0000" when x"3CA4",
			x"0000" when x"3CA5",
			x"0000" when x"3CA6",
			x"0000" when x"3CA7",
			x"0000" when x"3CA8",
			x"0000" when x"3CA9",
			x"0000" when x"3CAA",
			x"0000" when x"3CAB",
			x"0000" when x"3CAC",
			x"0000" when x"3CAD",
			x"0000" when x"3CAE",
			x"0000" when x"3CAF",
			x"0000" when x"3CB0",
			x"0000" when x"3CB1",
			x"0000" when x"3CB2",
			x"0000" when x"3CB3",
			x"0000" when x"3CB4",
			x"0000" when x"3CB5",
			x"0000" when x"3CB6",
			x"0000" when x"3CB7",
			x"0000" when x"3CB8",
			x"0000" when x"3CB9",
			x"0000" when x"3CBA",
			x"0000" when x"3CBB",
			x"0000" when x"3CBC",
			x"0000" when x"3CBD",
			x"0000" when x"3CBE",
			x"0000" when x"3CBF",
			x"0000" when x"3CC0",
			x"0000" when x"3CC1",
			x"0000" when x"3CC2",
			x"0000" when x"3CC3",
			x"0000" when x"3CC4",
			x"0000" when x"3CC5",
			x"0000" when x"3CC6",
			x"0000" when x"3CC7",
			x"0000" when x"3CC8",
			x"0000" when x"3CC9",
			x"0000" when x"3CCA",
			x"0000" when x"3CCB",
			x"0000" when x"3CCC",
			x"0000" when x"3CCD",
			x"0000" when x"3CCE",
			x"0000" when x"3CCF",
			x"0000" when x"3CD0",
			x"0000" when x"3CD1",
			x"0000" when x"3CD2",
			x"0000" when x"3CD3",
			x"0000" when x"3CD4",
			x"0000" when x"3CD5",
			x"0000" when x"3CD6",
			x"0000" when x"3CD7",
			x"0000" when x"3CD8",
			x"0000" when x"3CD9",
			x"0000" when x"3CDA",
			x"0000" when x"3CDB",
			x"0000" when x"3CDC",
			x"0000" when x"3CDD",
			x"0000" when x"3CDE",
			x"0000" when x"3CDF",
			x"0000" when x"3CE0",
			x"0000" when x"3CE1",
			x"0000" when x"3CE2",
			x"0000" when x"3CE3",
			x"0000" when x"3CE4",
			x"0000" when x"3CE5",
			x"0000" when x"3CE6",
			x"0000" when x"3CE7",
			x"0000" when x"3CE8",
			x"0000" when x"3CE9",
			x"0000" when x"3CEA",
			x"0000" when x"3CEB",
			x"0000" when x"3CEC",
			x"0000" when x"3CED",
			x"0000" when x"3CEE",
			x"0000" when x"3CEF",
			x"0000" when x"3CF0",
			x"0000" when x"3CF1",
			x"0000" when x"3CF2",
			x"0000" when x"3CF3",
			x"0000" when x"3CF4",
			x"0000" when x"3CF5",
			x"0000" when x"3CF6",
			x"0000" when x"3CF7",
			x"0000" when x"3CF8",
			x"0000" when x"3CF9",
			x"0000" when x"3CFA",
			x"0000" when x"3CFB",
			x"0000" when x"3CFC",
			x"0000" when x"3CFD",
			x"0000" when x"3CFE",
			x"0000" when x"3CFF",
			x"0000" when x"3D00",
			x"0000" when x"3D01",
			x"0000" when x"3D02",
			x"0000" when x"3D03",
			x"0000" when x"3D04",
			x"0000" when x"3D05",
			x"0000" when x"3D06",
			x"0000" when x"3D07",
			x"0000" when x"3D08",
			x"0000" when x"3D09",
			x"0000" when x"3D0A",
			x"0000" when x"3D0B",
			x"0000" when x"3D0C",
			x"0000" when x"3D0D",
			x"0000" when x"3D0E",
			x"0000" when x"3D0F",
			x"0000" when x"3D10",
			x"0000" when x"3D11",
			x"0000" when x"3D12",
			x"0000" when x"3D13",
			x"0000" when x"3D14",
			x"0000" when x"3D15",
			x"0000" when x"3D16",
			x"0000" when x"3D17",
			x"0000" when x"3D18",
			x"0000" when x"3D19",
			x"0000" when x"3D1A",
			x"0000" when x"3D1B",
			x"0000" when x"3D1C",
			x"0000" when x"3D1D",
			x"0000" when x"3D1E",
			x"0000" when x"3D1F",
			x"0000" when x"3D20",
			x"0000" when x"3D21",
			x"0000" when x"3D22",
			x"0000" when x"3D23",
			x"0000" when x"3D24",
			x"0000" when x"3D25",
			x"0000" when x"3D26",
			x"0000" when x"3D27",
			x"0000" when x"3D28",
			x"0000" when x"3D29",
			x"0000" when x"3D2A",
			x"0000" when x"3D2B",
			x"0000" when x"3D2C",
			x"0000" when x"3D2D",
			x"0000" when x"3D2E",
			x"0000" when x"3D2F",
			x"0000" when x"3D30",
			x"0000" when x"3D31",
			x"0000" when x"3D32",
			x"0000" when x"3D33",
			x"0000" when x"3D34",
			x"0000" when x"3D35",
			x"0000" when x"3D36",
			x"0000" when x"3D37",
			x"0000" when x"3D38",
			x"0000" when x"3D39",
			x"0000" when x"3D3A",
			x"0000" when x"3D3B",
			x"0000" when x"3D3C",
			x"0000" when x"3D3D",
			x"0000" when x"3D3E",
			x"0000" when x"3D3F",
			x"0000" when x"3D40",
			x"0000" when x"3D41",
			x"0000" when x"3D42",
			x"0000" when x"3D43",
			x"0000" when x"3D44",
			x"0000" when x"3D45",
			x"0000" when x"3D46",
			x"0000" when x"3D47",
			x"0000" when x"3D48",
			x"0000" when x"3D49",
			x"0000" when x"3D4A",
			x"0000" when x"3D4B",
			x"0000" when x"3D4C",
			x"0000" when x"3D4D",
			x"0000" when x"3D4E",
			x"0000" when x"3D4F",
			x"0000" when x"3D50",
			x"0000" when x"3D51",
			x"0000" when x"3D52",
			x"0000" when x"3D53",
			x"0000" when x"3D54",
			x"0000" when x"3D55",
			x"0000" when x"3D56",
			x"0000" when x"3D57",
			x"0000" when x"3D58",
			x"0000" when x"3D59",
			x"0000" when x"3D5A",
			x"0000" when x"3D5B",
			x"0000" when x"3D5C",
			x"0000" when x"3D5D",
			x"0000" when x"3D5E",
			x"0000" when x"3D5F",
			x"0000" when x"3D60",
			x"0000" when x"3D61",
			x"0000" when x"3D62",
			x"0000" when x"3D63",
			x"0000" when x"3D64",
			x"0000" when x"3D65",
			x"0000" when x"3D66",
			x"0000" when x"3D67",
			x"0000" when x"3D68",
			x"0000" when x"3D69",
			x"0000" when x"3D6A",
			x"0000" when x"3D6B",
			x"0000" when x"3D6C",
			x"0000" when x"3D6D",
			x"0000" when x"3D6E",
			x"0000" when x"3D6F",
			x"0000" when x"3D70",
			x"0000" when x"3D71",
			x"0000" when x"3D72",
			x"0000" when x"3D73",
			x"0000" when x"3D74",
			x"0000" when x"3D75",
			x"0000" when x"3D76",
			x"0000" when x"3D77",
			x"0000" when x"3D78",
			x"0000" when x"3D79",
			x"0000" when x"3D7A",
			x"0000" when x"3D7B",
			x"0000" when x"3D7C",
			x"0000" when x"3D7D",
			x"0000" when x"3D7E",
			x"0000" when x"3D7F",
			x"0000" when x"3D80",
			x"0000" when x"3D81",
			x"0000" when x"3D82",
			x"0000" when x"3D83",
			x"0000" when x"3D84",
			x"0000" when x"3D85",
			x"0000" when x"3D86",
			x"0000" when x"3D87",
			x"0000" when x"3D88",
			x"0000" when x"3D89",
			x"0000" when x"3D8A",
			x"0000" when x"3D8B",
			x"0000" when x"3D8C",
			x"0000" when x"3D8D",
			x"0000" when x"3D8E",
			x"0000" when x"3D8F",
			x"0000" when x"3D90",
			x"0000" when x"3D91",
			x"0000" when x"3D92",
			x"0000" when x"3D93",
			x"0000" when x"3D94",
			x"0000" when x"3D95",
			x"0000" when x"3D96",
			x"0000" when x"3D97",
			x"0000" when x"3D98",
			x"0000" when x"3D99",
			x"0000" when x"3D9A",
			x"0000" when x"3D9B",
			x"0000" when x"3D9C",
			x"0000" when x"3D9D",
			x"0000" when x"3D9E",
			x"0000" when x"3D9F",
			x"0000" when x"3DA0",
			x"0000" when x"3DA1",
			x"0000" when x"3DA2",
			x"0000" when x"3DA3",
			x"0000" when x"3DA4",
			x"0000" when x"3DA5",
			x"0000" when x"3DA6",
			x"0000" when x"3DA7",
			x"0000" when x"3DA8",
			x"0000" when x"3DA9",
			x"0000" when x"3DAA",
			x"0000" when x"3DAB",
			x"0000" when x"3DAC",
			x"0000" when x"3DAD",
			x"0000" when x"3DAE",
			x"0000" when x"3DAF",
			x"0000" when x"3DB0",
			x"0000" when x"3DB1",
			x"0000" when x"3DB2",
			x"0000" when x"3DB3",
			x"0000" when x"3DB4",
			x"0000" when x"3DB5",
			x"0000" when x"3DB6",
			x"0000" when x"3DB7",
			x"0000" when x"3DB8",
			x"0000" when x"3DB9",
			x"0000" when x"3DBA",
			x"0000" when x"3DBB",
			x"0000" when x"3DBC",
			x"0000" when x"3DBD",
			x"0000" when x"3DBE",
			x"0000" when x"3DBF",
			x"0000" when x"3DC0",
			x"0000" when x"3DC1",
			x"0000" when x"3DC2",
			x"0000" when x"3DC3",
			x"0000" when x"3DC4",
			x"0000" when x"3DC5",
			x"0000" when x"3DC6",
			x"0000" when x"3DC7",
			x"0000" when x"3DC8",
			x"0000" when x"3DC9",
			x"0000" when x"3DCA",
			x"0000" when x"3DCB",
			x"0000" when x"3DCC",
			x"0000" when x"3DCD",
			x"0000" when x"3DCE",
			x"0000" when x"3DCF",
			x"0000" when x"3DD0",
			x"0000" when x"3DD1",
			x"0000" when x"3DD2",
			x"0000" when x"3DD3",
			x"0000" when x"3DD4",
			x"0000" when x"3DD5",
			x"0000" when x"3DD6",
			x"0000" when x"3DD7",
			x"0000" when x"3DD8",
			x"0000" when x"3DD9",
			x"0000" when x"3DDA",
			x"0000" when x"3DDB",
			x"0000" when x"3DDC",
			x"0000" when x"3DDD",
			x"0000" when x"3DDE",
			x"0000" when x"3DDF",
			x"0000" when x"3DE0",
			x"0000" when x"3DE1",
			x"0000" when x"3DE2",
			x"0000" when x"3DE3",
			x"0000" when x"3DE4",
			x"0000" when x"3DE5",
			x"0000" when x"3DE6",
			x"0000" when x"3DE7",
			x"0000" when x"3DE8",
			x"0000" when x"3DE9",
			x"0000" when x"3DEA",
			x"0000" when x"3DEB",
			x"0000" when x"3DEC",
			x"0000" when x"3DED",
			x"0000" when x"3DEE",
			x"0000" when x"3DEF",
			x"0000" when x"3DF0",
			x"0000" when x"3DF1",
			x"0000" when x"3DF2",
			x"0000" when x"3DF3",
			x"0000" when x"3DF4",
			x"0000" when x"3DF5",
			x"0000" when x"3DF6",
			x"0000" when x"3DF7",
			x"0000" when x"3DF8",
			x"0000" when x"3DF9",
			x"0000" when x"3DFA",
			x"0000" when x"3DFB",
			x"0000" when x"3DFC",
			x"0000" when x"3DFD",
			x"0000" when x"3DFE",
			x"0000" when x"3DFF",
			x"0000" when x"3E00",
			x"0000" when x"3E01",
			x"0000" when x"3E02",
			x"0000" when x"3E03",
			x"0000" when x"3E04",
			x"0000" when x"3E05",
			x"0000" when x"3E06",
			x"0000" when x"3E07",
			x"0000" when x"3E08",
			x"0000" when x"3E09",
			x"0000" when x"3E0A",
			x"0000" when x"3E0B",
			x"0000" when x"3E0C",
			x"0000" when x"3E0D",
			x"0000" when x"3E0E",
			x"0000" when x"3E0F",
			x"0000" when x"3E10",
			x"0000" when x"3E11",
			x"0000" when x"3E12",
			x"0000" when x"3E13",
			x"0000" when x"3E14",
			x"0000" when x"3E15",
			x"0000" when x"3E16",
			x"0000" when x"3E17",
			x"0000" when x"3E18",
			x"0000" when x"3E19",
			x"0000" when x"3E1A",
			x"0000" when x"3E1B",
			x"0000" when x"3E1C",
			x"0000" when x"3E1D",
			x"0000" when x"3E1E",
			x"0000" when x"3E1F",
			x"0000" when x"3E20",
			x"0000" when x"3E21",
			x"0000" when x"3E22",
			x"0000" when x"3E23",
			x"0000" when x"3E24",
			x"0000" when x"3E25",
			x"0000" when x"3E26",
			x"0000" when x"3E27",
			x"0000" when x"3E28",
			x"0000" when x"3E29",
			x"0000" when x"3E2A",
			x"0000" when x"3E2B",
			x"0000" when x"3E2C",
			x"0000" when x"3E2D",
			x"0000" when x"3E2E",
			x"0000" when x"3E2F",
			x"0000" when x"3E30",
			x"0000" when x"3E31",
			x"0000" when x"3E32",
			x"0000" when x"3E33",
			x"0000" when x"3E34",
			x"0000" when x"3E35",
			x"0000" when x"3E36",
			x"0000" when x"3E37",
			x"0000" when x"3E38",
			x"0000" when x"3E39",
			x"0000" when x"3E3A",
			x"0000" when x"3E3B",
			x"0000" when x"3E3C",
			x"0000" when x"3E3D",
			x"0000" when x"3E3E",
			x"0000" when x"3E3F",
			x"0000" when x"3E40",
			x"0000" when x"3E41",
			x"0000" when x"3E42",
			x"0000" when x"3E43",
			x"0000" when x"3E44",
			x"0000" when x"3E45",
			x"0000" when x"3E46",
			x"0000" when x"3E47",
			x"0000" when x"3E48",
			x"0000" when x"3E49",
			x"0000" when x"3E4A",
			x"0000" when x"3E4B",
			x"0000" when x"3E4C",
			x"0000" when x"3E4D",
			x"0000" when x"3E4E",
			x"0000" when x"3E4F",
			x"0000" when x"3E50",
			x"0000" when x"3E51",
			x"0000" when x"3E52",
			x"0000" when x"3E53",
			x"0000" when x"3E54",
			x"0000" when x"3E55",
			x"0000" when x"3E56",
			x"0000" when x"3E57",
			x"0000" when x"3E58",
			x"0000" when x"3E59",
			x"0000" when x"3E5A",
			x"0000" when x"3E5B",
			x"0000" when x"3E5C",
			x"0000" when x"3E5D",
			x"0000" when x"3E5E",
			x"0000" when x"3E5F",
			x"0000" when x"3E60",
			x"0000" when x"3E61",
			x"0000" when x"3E62",
			x"0000" when x"3E63",
			x"0000" when x"3E64",
			x"0000" when x"3E65",
			x"0000" when x"3E66",
			x"0000" when x"3E67",
			x"0000" when x"3E68",
			x"0000" when x"3E69",
			x"0000" when x"3E6A",
			x"0000" when x"3E6B",
			x"0000" when x"3E6C",
			x"0000" when x"3E6D",
			x"0000" when x"3E6E",
			x"0000" when x"3E6F",
			x"0000" when x"3E70",
			x"0000" when x"3E71",
			x"0000" when x"3E72",
			x"0000" when x"3E73",
			x"0000" when x"3E74",
			x"0000" when x"3E75",
			x"0000" when x"3E76",
			x"0000" when x"3E77",
			x"0000" when x"3E78",
			x"0000" when x"3E79",
			x"0000" when x"3E7A",
			x"0000" when x"3E7B",
			x"0000" when x"3E7C",
			x"0000" when x"3E7D",
			x"0000" when x"3E7E",
			x"0000" when x"3E7F",
			x"0000" when x"3E80",
			x"0000" when x"3E81",
			x"0000" when x"3E82",
			x"0000" when x"3E83",
			x"0000" when x"3E84",
			x"0000" when x"3E85",
			x"0000" when x"3E86",
			x"0000" when x"3E87",
			x"0000" when x"3E88",
			x"0000" when x"3E89",
			x"0000" when x"3E8A",
			x"0000" when x"3E8B",
			x"0000" when x"3E8C",
			x"0000" when x"3E8D",
			x"0000" when x"3E8E",
			x"0000" when x"3E8F",
			x"0000" when x"3E90",
			x"0000" when x"3E91",
			x"0000" when x"3E92",
			x"0000" when x"3E93",
			x"0000" when x"3E94",
			x"0000" when x"3E95",
			x"0000" when x"3E96",
			x"0000" when x"3E97",
			x"0000" when x"3E98",
			x"0000" when x"3E99",
			x"0000" when x"3E9A",
			x"0000" when x"3E9B",
			x"0000" when x"3E9C",
			x"0000" when x"3E9D",
			x"0000" when x"3E9E",
			x"0000" when x"3E9F",
			x"0000" when x"3EA0",
			x"0000" when x"3EA1",
			x"0000" when x"3EA2",
			x"0000" when x"3EA3",
			x"0000" when x"3EA4",
			x"0000" when x"3EA5",
			x"0000" when x"3EA6",
			x"0000" when x"3EA7",
			x"0000" when x"3EA8",
			x"0000" when x"3EA9",
			x"0000" when x"3EAA",
			x"0000" when x"3EAB",
			x"0000" when x"3EAC",
			x"0000" when x"3EAD",
			x"0000" when x"3EAE",
			x"0000" when x"3EAF",
			x"0000" when x"3EB0",
			x"0000" when x"3EB1",
			x"0000" when x"3EB2",
			x"0000" when x"3EB3",
			x"0000" when x"3EB4",
			x"0000" when x"3EB5",
			x"0000" when x"3EB6",
			x"0000" when x"3EB7",
			x"0000" when x"3EB8",
			x"0000" when x"3EB9",
			x"0000" when x"3EBA",
			x"0000" when x"3EBB",
			x"0000" when x"3EBC",
			x"0000" when x"3EBD",
			x"0000" when x"3EBE",
			x"0000" when x"3EBF",
			x"0000" when x"3EC0",
			x"0000" when x"3EC1",
			x"0000" when x"3EC2",
			x"0000" when x"3EC3",
			x"0000" when x"3EC4",
			x"0000" when x"3EC5",
			x"0000" when x"3EC6",
			x"0000" when x"3EC7",
			x"0000" when x"3EC8",
			x"0000" when x"3EC9",
			x"0000" when x"3ECA",
			x"0000" when x"3ECB",
			x"0000" when x"3ECC",
			x"0000" when x"3ECD",
			x"0000" when x"3ECE",
			x"0000" when x"3ECF",
			x"0000" when x"3ED0",
			x"0000" when x"3ED1",
			x"0000" when x"3ED2",
			x"0000" when x"3ED3",
			x"0000" when x"3ED4",
			x"0000" when x"3ED5",
			x"0000" when x"3ED6",
			x"0000" when x"3ED7",
			x"0000" when x"3ED8",
			x"0000" when x"3ED9",
			x"0000" when x"3EDA",
			x"0000" when x"3EDB",
			x"0000" when x"3EDC",
			x"0000" when x"3EDD",
			x"0000" when x"3EDE",
			x"0000" when x"3EDF",
			x"0000" when x"3EE0",
			x"0000" when x"3EE1",
			x"0000" when x"3EE2",
			x"0000" when x"3EE3",
			x"0000" when x"3EE4",
			x"0000" when x"3EE5",
			x"0000" when x"3EE6",
			x"0000" when x"3EE7",
			x"0000" when x"3EE8",
			x"0000" when x"3EE9",
			x"0000" when x"3EEA",
			x"0000" when x"3EEB",
			x"0000" when x"3EEC",
			x"0000" when x"3EED",
			x"0000" when x"3EEE",
			x"0000" when x"3EEF",
			x"0000" when x"3EF0",
			x"0000" when x"3EF1",
			x"0000" when x"3EF2",
			x"0000" when x"3EF3",
			x"0000" when x"3EF4",
			x"0000" when x"3EF5",
			x"0000" when x"3EF6",
			x"0000" when x"3EF7",
			x"0000" when x"3EF8",
			x"0000" when x"3EF9",
			x"0000" when x"3EFA",
			x"0000" when x"3EFB",
			x"0000" when x"3EFC",
			x"0000" when x"3EFD",
			x"0000" when x"3EFE",
			x"0000" when x"3EFF",
			x"0000" when x"3F00",
			x"0000" when x"3F01",
			x"0000" when x"3F02",
			x"0000" when x"3F03",
			x"0000" when x"3F04",
			x"0000" when x"3F05",
			x"0000" when x"3F06",
			x"0000" when x"3F07",
			x"0000" when x"3F08",
			x"0000" when x"3F09",
			x"0000" when x"3F0A",
			x"0000" when x"3F0B",
			x"0000" when x"3F0C",
			x"0000" when x"3F0D",
			x"0000" when x"3F0E",
			x"0000" when x"3F0F",
			x"0000" when x"3F10",
			x"0000" when x"3F11",
			x"0000" when x"3F12",
			x"0000" when x"3F13",
			x"0000" when x"3F14",
			x"0000" when x"3F15",
			x"0000" when x"3F16",
			x"0000" when x"3F17",
			x"0000" when x"3F18",
			x"0000" when x"3F19",
			x"0000" when x"3F1A",
			x"0000" when x"3F1B",
			x"0000" when x"3F1C",
			x"0000" when x"3F1D",
			x"0000" when x"3F1E",
			x"0000" when x"3F1F",
			x"0000" when x"3F20",
			x"0000" when x"3F21",
			x"0000" when x"3F22",
			x"0000" when x"3F23",
			x"0000" when x"3F24",
			x"0000" when x"3F25",
			x"0000" when x"3F26",
			x"0000" when x"3F27",
			x"0000" when x"3F28",
			x"0000" when x"3F29",
			x"0000" when x"3F2A",
			x"0000" when x"3F2B",
			x"0000" when x"3F2C",
			x"0000" when x"3F2D",
			x"0000" when x"3F2E",
			x"0000" when x"3F2F",
			x"0000" when x"3F30",
			x"0000" when x"3F31",
			x"0000" when x"3F32",
			x"0000" when x"3F33",
			x"0000" when x"3F34",
			x"0000" when x"3F35",
			x"0000" when x"3F36",
			x"0000" when x"3F37",
			x"0000" when x"3F38",
			x"0000" when x"3F39",
			x"0000" when x"3F3A",
			x"0000" when x"3F3B",
			x"0000" when x"3F3C",
			x"0000" when x"3F3D",
			x"0000" when x"3F3E",
			x"0000" when x"3F3F",
			x"0000" when x"3F40",
			x"0000" when x"3F41",
			x"0000" when x"3F42",
			x"0000" when x"3F43",
			x"0000" when x"3F44",
			x"0000" when x"3F45",
			x"0000" when x"3F46",
			x"0000" when x"3F47",
			x"0000" when x"3F48",
			x"0000" when x"3F49",
			x"0000" when x"3F4A",
			x"0000" when x"3F4B",
			x"0000" when x"3F4C",
			x"0000" when x"3F4D",
			x"0000" when x"3F4E",
			x"0000" when x"3F4F",
			x"0000" when x"3F50",
			x"0000" when x"3F51",
			x"0000" when x"3F52",
			x"0000" when x"3F53",
			x"0000" when x"3F54",
			x"0000" when x"3F55",
			x"0000" when x"3F56",
			x"0000" when x"3F57",
			x"0000" when x"3F58",
			x"0000" when x"3F59",
			x"0000" when x"3F5A",
			x"0000" when x"3F5B",
			x"0000" when x"3F5C",
			x"0000" when x"3F5D",
			x"0000" when x"3F5E",
			x"0000" when x"3F5F",
			x"0000" when x"3F60",
			x"0000" when x"3F61",
			x"0000" when x"3F62",
			x"0000" when x"3F63",
			x"0000" when x"3F64",
			x"0000" when x"3F65",
			x"0000" when x"3F66",
			x"0000" when x"3F67",
			x"0000" when x"3F68",
			x"0000" when x"3F69",
			x"0000" when x"3F6A",
			x"0000" when x"3F6B",
			x"0000" when x"3F6C",
			x"0000" when x"3F6D",
			x"0000" when x"3F6E",
			x"0000" when x"3F6F",
			x"0000" when x"3F70",
			x"0000" when x"3F71",
			x"0000" when x"3F72",
			x"0000" when x"3F73",
			x"0000" when x"3F74",
			x"0000" when x"3F75",
			x"0000" when x"3F76",
			x"0000" when x"3F77",
			x"0000" when x"3F78",
			x"0000" when x"3F79",
			x"0000" when x"3F7A",
			x"0000" when x"3F7B",
			x"0000" when x"3F7C",
			x"0000" when x"3F7D",
			x"0000" when x"3F7E",
			x"0000" when x"3F7F",
			x"0000" when x"3F80",
			x"0000" when x"3F81",
			x"0000" when x"3F82",
			x"0000" when x"3F83",
			x"0000" when x"3F84",
			x"0000" when x"3F85",
			x"0000" when x"3F86",
			x"0000" when x"3F87",
			x"0000" when x"3F88",
			x"0000" when x"3F89",
			x"0000" when x"3F8A",
			x"0000" when x"3F8B",
			x"0000" when x"3F8C",
			x"0000" when x"3F8D",
			x"0000" when x"3F8E",
			x"0000" when x"3F8F",
			x"0000" when x"3F90",
			x"0000" when x"3F91",
			x"0000" when x"3F92",
			x"0000" when x"3F93",
			x"0000" when x"3F94",
			x"0000" when x"3F95",
			x"0000" when x"3F96",
			x"0000" when x"3F97",
			x"0000" when x"3F98",
			x"0000" when x"3F99",
			x"0000" when x"3F9A",
			x"0000" when x"3F9B",
			x"0000" when x"3F9C",
			x"0000" when x"3F9D",
			x"0000" when x"3F9E",
			x"0000" when x"3F9F",
			x"0000" when x"3FA0",
			x"0000" when x"3FA1",
			x"0000" when x"3FA2",
			x"0000" when x"3FA3",
			x"0000" when x"3FA4",
			x"0000" when x"3FA5",
			x"0000" when x"3FA6",
			x"0000" when x"3FA7",
			x"0000" when x"3FA8",
			x"0000" when x"3FA9",
			x"0000" when x"3FAA",
			x"0000" when x"3FAB",
			x"0000" when x"3FAC",
			x"0000" when x"3FAD",
			x"0000" when x"3FAE",
			x"0000" when x"3FAF",
			x"0000" when x"3FB0",
			x"0000" when x"3FB1",
			x"0000" when x"3FB2",
			x"0000" when x"3FB3",
			x"0000" when x"3FB4",
			x"0000" when x"3FB5",
			x"0000" when x"3FB6",
			x"0000" when x"3FB7",
			x"0000" when x"3FB8",
			x"0000" when x"3FB9",
			x"0000" when x"3FBA",
			x"0000" when x"3FBB",
			x"0000" when x"3FBC",
			x"0000" when x"3FBD",
			x"0000" when x"3FBE",
			x"0000" when x"3FBF",
			x"0000" when x"3FC0",
			x"0000" when x"3FC1",
			x"0000" when x"3FC2",
			x"0000" when x"3FC3",
			x"0000" when x"3FC4",
			x"0000" when x"3FC5",
			x"0000" when x"3FC6",
			x"0000" when x"3FC7",
			x"0000" when x"3FC8",
			x"0000" when x"3FC9",
			x"0000" when x"3FCA",
			x"0000" when x"3FCB",
			x"0000" when x"3FCC",
			x"0000" when x"3FCD",
			x"0000" when x"3FCE",
			x"0000" when x"3FCF",
			x"0000" when x"3FD0",
			x"0000" when x"3FD1",
			x"0000" when x"3FD2",
			x"0000" when x"3FD3",
			x"0000" when x"3FD4",
			x"0000" when x"3FD5",
			x"0000" when x"3FD6",
			x"0000" when x"3FD7",
			x"0000" when x"3FD8",
			x"0000" when x"3FD9",
			x"0000" when x"3FDA",
			x"0000" when x"3FDB",
			x"0000" when x"3FDC",
			x"0000" when x"3FDD",
			x"0000" when x"3FDE",
			x"0000" when x"3FDF",
			x"0000" when x"3FE0",
			x"0000" when x"3FE1",
			x"0000" when x"3FE2",
			x"0000" when x"3FE3",
			x"0000" when x"3FE4",
			x"0000" when x"3FE5",
			x"0000" when x"3FE6",
			x"0000" when x"3FE7",
			x"0000" when x"3FE8",
			x"0000" when x"3FE9",
			x"0000" when x"3FEA",
			x"0000" when x"3FEB",
			x"0000" when x"3FEC",
			x"0000" when x"3FED",
			x"0000" when x"3FEE",
			x"0000" when x"3FEF",
			x"0000" when x"3FF0",
			x"0000" when x"3FF1",
			x"0000" when x"3FF2",
			x"0000" when x"3FF3",
			x"0000" when x"3FF4",
			x"0000" when x"3FF5",
			x"0000" when x"3FF6",
			x"0000" when x"3FF7",
			x"0000" when x"3FF8",
			x"0000" when x"3FF9",
			x"0000" when x"3FFA",
			x"0000" when x"3FFB",
			x"0000" when x"3FFC",
			x"0000" when x"3FFD",
			x"0000" when x"3FFE",
			x"0000" when x"3FFF",
			x"0000" when x"4000",
			x"0000" when x"4001",
			x"0000" when x"4002",
			x"0000" when x"4003",
			x"0000" when x"4004",
			x"0000" when x"4005",
			x"0000" when x"4006",
			x"0000" when x"4007",
			x"0000" when x"4008",
			x"0000" when x"4009",
			x"0000" when x"400A",
			x"0000" when x"400B",
			x"0000" when x"400C",
			x"0000" when x"400D",
			x"0000" when x"400E",
			x"0000" when x"400F",
			x"0000" when x"4010",
			x"0000" when x"4011",
			x"0000" when x"4012",
			x"0000" when x"4013",
			x"0000" when x"4014",
			x"0000" when x"4015",
			x"0000" when x"4016",
			x"0000" when x"4017",
			x"0000" when x"4018",
			x"0000" when x"4019",
			x"0000" when x"401A",
			x"0000" when x"401B",
			x"0000" when x"401C",
			x"0000" when x"401D",
			x"0000" when x"401E",
			x"0000" when x"401F",
			x"0000" when x"4020",
			x"0000" when x"4021",
			x"0000" when x"4022",
			x"0000" when x"4023",
			x"0000" when x"4024",
			x"0000" when x"4025",
			x"0000" when x"4026",
			x"0000" when x"4027",
			x"0000" when x"4028",
			x"0000" when x"4029",
			x"0000" when x"402A",
			x"0000" when x"402B",
			x"0000" when x"402C",
			x"0000" when x"402D",
			x"0000" when x"402E",
			x"0000" when x"402F",
			x"0000" when x"4030",
			x"0000" when x"4031",
			x"0000" when x"4032",
			x"0000" when x"4033",
			x"0000" when x"4034",
			x"0000" when x"4035",
			x"0000" when x"4036",
			x"0000" when x"4037",
			x"0000" when x"4038",
			x"0000" when x"4039",
			x"0000" when x"403A",
			x"0000" when x"403B",
			x"0000" when x"403C",
			x"0000" when x"403D",
			x"0000" when x"403E",
			x"0000" when x"403F",
			x"0000" when x"4040",
			x"0000" when x"4041",
			x"0000" when x"4042",
			x"0000" when x"4043",
			x"0000" when x"4044",
			x"0000" when x"4045",
			x"0000" when x"4046",
			x"0000" when x"4047",
			x"0000" when x"4048",
			x"0000" when x"4049",
			x"0000" when x"404A",
			x"0000" when x"404B",
			x"0000" when x"404C",
			x"0000" when x"404D",
			x"0000" when x"404E",
			x"0000" when x"404F",
			x"0000" when x"4050",
			x"0000" when x"4051",
			x"0000" when x"4052",
			x"0000" when x"4053",
			x"0000" when x"4054",
			x"0000" when x"4055",
			x"0000" when x"4056",
			x"0000" when x"4057",
			x"0000" when x"4058",
			x"0000" when x"4059",
			x"0000" when x"405A",
			x"0000" when x"405B",
			x"0000" when x"405C",
			x"0000" when x"405D",
			x"0000" when x"405E",
			x"0000" when x"405F",
			x"0000" when x"4060",
			x"0000" when x"4061",
			x"0000" when x"4062",
			x"0000" when x"4063",
			x"0000" when x"4064",
			x"0000" when x"4065",
			x"0000" when x"4066",
			x"0000" when x"4067",
			x"0000" when x"4068",
			x"0000" when x"4069",
			x"0000" when x"406A",
			x"0000" when x"406B",
			x"0000" when x"406C",
			x"0000" when x"406D",
			x"0000" when x"406E",
			x"0000" when x"406F",
			x"0000" when x"4070",
			x"0000" when x"4071",
			x"0000" when x"4072",
			x"0000" when x"4073",
			x"0000" when x"4074",
			x"0000" when x"4075",
			x"0000" when x"4076",
			x"0000" when x"4077",
			x"0000" when x"4078",
			x"0000" when x"4079",
			x"0000" when x"407A",
			x"0000" when x"407B",
			x"0000" when x"407C",
			x"0000" when x"407D",
			x"0000" when x"407E",
			x"0000" when x"407F",
			x"0000" when x"4080",
			x"0000" when x"4081",
			x"0000" when x"4082",
			x"0000" when x"4083",
			x"0000" when x"4084",
			x"0000" when x"4085",
			x"0000" when x"4086",
			x"0000" when x"4087",
			x"0000" when x"4088",
			x"0000" when x"4089",
			x"0000" when x"408A",
			x"0000" when x"408B",
			x"0000" when x"408C",
			x"0000" when x"408D",
			x"0000" when x"408E",
			x"0000" when x"408F",
			x"0000" when x"4090",
			x"0000" when x"4091",
			x"0000" when x"4092",
			x"0000" when x"4093",
			x"0000" when x"4094",
			x"0000" when x"4095",
			x"0000" when x"4096",
			x"0000" when x"4097",
			x"0000" when x"4098",
			x"0000" when x"4099",
			x"0000" when x"409A",
			x"0000" when x"409B",
			x"0000" when x"409C",
			x"0000" when x"409D",
			x"0000" when x"409E",
			x"0000" when x"409F",
			x"0000" when x"40A0",
			x"0000" when x"40A1",
			x"0000" when x"40A2",
			x"0000" when x"40A3",
			x"0000" when x"40A4",
			x"0000" when x"40A5",
			x"0000" when x"40A6",
			x"0000" when x"40A7",
			x"0000" when x"40A8",
			x"0000" when x"40A9",
			x"0000" when x"40AA",
			x"0000" when x"40AB",
			x"0000" when x"40AC",
			x"0000" when x"40AD",
			x"0000" when x"40AE",
			x"0000" when x"40AF",
			x"0000" when x"40B0",
			x"0000" when x"40B1",
			x"0000" when x"40B2",
			x"0000" when x"40B3",
			x"0000" when x"40B4",
			x"0000" when x"40B5",
			x"0000" when x"40B6",
			x"0000" when x"40B7",
			x"0000" when x"40B8",
			x"0000" when x"40B9",
			x"0000" when x"40BA",
			x"0000" when x"40BB",
			x"0000" when x"40BC",
			x"0000" when x"40BD",
			x"0000" when x"40BE",
			x"0000" when x"40BF",
			x"0000" when x"40C0",
			x"0000" when x"40C1",
			x"0000" when x"40C2",
			x"0000" when x"40C3",
			x"0000" when x"40C4",
			x"0000" when x"40C5",
			x"0000" when x"40C6",
			x"0000" when x"40C7",
			x"0000" when x"40C8",
			x"0000" when x"40C9",
			x"0000" when x"40CA",
			x"0000" when x"40CB",
			x"0000" when x"40CC",
			x"0000" when x"40CD",
			x"0000" when x"40CE",
			x"0000" when x"40CF",
			x"0000" when x"40D0",
			x"0000" when x"40D1",
			x"0000" when x"40D2",
			x"0000" when x"40D3",
			x"0000" when x"40D4",
			x"0000" when x"40D5",
			x"0000" when x"40D6",
			x"0000" when x"40D7",
			x"0000" when x"40D8",
			x"0000" when x"40D9",
			x"0000" when x"40DA",
			x"0000" when x"40DB",
			x"0000" when x"40DC",
			x"0000" when x"40DD",
			x"0000" when x"40DE",
			x"0000" when x"40DF",
			x"0000" when x"40E0",
			x"0000" when x"40E1",
			x"0000" when x"40E2",
			x"0000" when x"40E3",
			x"0000" when x"40E4",
			x"0000" when x"40E5",
			x"0000" when x"40E6",
			x"0000" when x"40E7",
			x"0000" when x"40E8",
			x"0000" when x"40E9",
			x"0000" when x"40EA",
			x"0000" when x"40EB",
			x"0000" when x"40EC",
			x"0000" when x"40ED",
			x"0000" when x"40EE",
			x"0000" when x"40EF",
			x"0000" when x"40F0",
			x"0000" when x"40F1",
			x"0000" when x"40F2",
			x"0000" when x"40F3",
			x"0000" when x"40F4",
			x"0000" when x"40F5",
			x"0000" when x"40F6",
			x"0000" when x"40F7",
			x"0000" when x"40F8",
			x"0000" when x"40F9",
			x"0000" when x"40FA",
			x"0000" when x"40FB",
			x"0000" when x"40FC",
			x"0000" when x"40FD",
			x"0000" when x"40FE",
			x"0000" when x"40FF",
			x"0000" when x"4100",
			x"0000" when x"4101",
			x"0000" when x"4102",
			x"0000" when x"4103",
			x"0000" when x"4104",
			x"0000" when x"4105",
			x"0000" when x"4106",
			x"0000" when x"4107",
			x"0000" when x"4108",
			x"0000" when x"4109",
			x"0000" when x"410A",
			x"0000" when x"410B",
			x"0000" when x"410C",
			x"0000" when x"410D",
			x"0000" when x"410E",
			x"0000" when x"410F",
			x"0000" when x"4110",
			x"0000" when x"4111",
			x"0000" when x"4112",
			x"0000" when x"4113",
			x"0000" when x"4114",
			x"0000" when x"4115",
			x"0000" when x"4116",
			x"0000" when x"4117",
			x"0000" when x"4118",
			x"0000" when x"4119",
			x"0000" when x"411A",
			x"0000" when x"411B",
			x"0000" when x"411C",
			x"0000" when x"411D",
			x"0000" when x"411E",
			x"0000" when x"411F",
			x"0000" when x"4120",
			x"0000" when x"4121",
			x"0000" when x"4122",
			x"0000" when x"4123",
			x"0000" when x"4124",
			x"0000" when x"4125",
			x"0000" when x"4126",
			x"0000" when x"4127",
			x"0000" when x"4128",
			x"0000" when x"4129",
			x"0000" when x"412A",
			x"0000" when x"412B",
			x"0000" when x"412C",
			x"0000" when x"412D",
			x"0000" when x"412E",
			x"0000" when x"412F",
			x"0000" when x"4130",
			x"0000" when x"4131",
			x"0000" when x"4132",
			x"0000" when x"4133",
			x"0000" when x"4134",
			x"0000" when x"4135",
			x"0000" when x"4136",
			x"0000" when x"4137",
			x"0000" when x"4138",
			x"0000" when x"4139",
			x"0000" when x"413A",
			x"0000" when x"413B",
			x"0000" when x"413C",
			x"0000" when x"413D",
			x"0000" when x"413E",
			x"0000" when x"413F",
			x"0000" when x"4140",
			x"0000" when x"4141",
			x"0000" when x"4142",
			x"0000" when x"4143",
			x"0000" when x"4144",
			x"0000" when x"4145",
			x"0000" when x"4146",
			x"0000" when x"4147",
			x"0000" when x"4148",
			x"0000" when x"4149",
			x"0000" when x"414A",
			x"0000" when x"414B",
			x"0000" when x"414C",
			x"0000" when x"414D",
			x"0000" when x"414E",
			x"0000" when x"414F",
			x"0000" when x"4150",
			x"0000" when x"4151",
			x"0000" when x"4152",
			x"0000" when x"4153",
			x"0000" when x"4154",
			x"0000" when x"4155",
			x"0000" when x"4156",
			x"0000" when x"4157",
			x"0000" when x"4158",
			x"0000" when x"4159",
			x"0000" when x"415A",
			x"0000" when x"415B",
			x"0000" when x"415C",
			x"0000" when x"415D",
			x"0000" when x"415E",
			x"0000" when x"415F",
			x"0000" when x"4160",
			x"0000" when x"4161",
			x"0000" when x"4162",
			x"0000" when x"4163",
			x"0000" when x"4164",
			x"0000" when x"4165",
			x"0000" when x"4166",
			x"0000" when x"4167",
			x"0000" when x"4168",
			x"0000" when x"4169",
			x"0000" when x"416A",
			x"0000" when x"416B",
			x"0000" when x"416C",
			x"0000" when x"416D",
			x"0000" when x"416E",
			x"0000" when x"416F",
			x"0000" when x"4170",
			x"0000" when x"4171",
			x"0000" when x"4172",
			x"0000" when x"4173",
			x"0000" when x"4174",
			x"0000" when x"4175",
			x"0000" when x"4176",
			x"0000" when x"4177",
			x"0000" when x"4178",
			x"0000" when x"4179",
			x"0000" when x"417A",
			x"0000" when x"417B",
			x"0000" when x"417C",
			x"0000" when x"417D",
			x"0000" when x"417E",
			x"0000" when x"417F",
			x"0000" when x"4180",
			x"0000" when x"4181",
			x"0000" when x"4182",
			x"0000" when x"4183",
			x"0000" when x"4184",
			x"0000" when x"4185",
			x"0000" when x"4186",
			x"0000" when x"4187",
			x"0000" when x"4188",
			x"0000" when x"4189",
			x"0000" when x"418A",
			x"0000" when x"418B",
			x"0000" when x"418C",
			x"0000" when x"418D",
			x"0000" when x"418E",
			x"0000" when x"418F",
			x"0000" when x"4190",
			x"0000" when x"4191",
			x"0000" when x"4192",
			x"0000" when x"4193",
			x"0000" when x"4194",
			x"0000" when x"4195",
			x"0000" when x"4196",
			x"0000" when x"4197",
			x"0000" when x"4198",
			x"0000" when x"4199",
			x"0000" when x"419A",
			x"0000" when x"419B",
			x"0000" when x"419C",
			x"0000" when x"419D",
			x"0000" when x"419E",
			x"0000" when x"419F",
			x"0000" when x"41A0",
			x"0000" when x"41A1",
			x"0000" when x"41A2",
			x"0000" when x"41A3",
			x"0000" when x"41A4",
			x"0000" when x"41A5",
			x"0000" when x"41A6",
			x"0000" when x"41A7",
			x"0000" when x"41A8",
			x"0000" when x"41A9",
			x"0000" when x"41AA",
			x"0000" when x"41AB",
			x"0000" when x"41AC",
			x"0000" when x"41AD",
			x"0000" when x"41AE",
			x"0000" when x"41AF",
			x"0000" when x"41B0",
			x"0000" when x"41B1",
			x"0000" when x"41B2",
			x"0000" when x"41B3",
			x"0000" when x"41B4",
			x"0000" when x"41B5",
			x"0000" when x"41B6",
			x"0000" when x"41B7",
			x"0000" when x"41B8",
			x"0000" when x"41B9",
			x"0000" when x"41BA",
			x"0000" when x"41BB",
			x"0000" when x"41BC",
			x"0000" when x"41BD",
			x"0000" when x"41BE",
			x"0000" when x"41BF",
			x"0000" when x"41C0",
			x"0000" when x"41C1",
			x"0000" when x"41C2",
			x"0000" when x"41C3",
			x"0000" when x"41C4",
			x"0000" when x"41C5",
			x"0000" when x"41C6",
			x"0000" when x"41C7",
			x"0000" when x"41C8",
			x"0000" when x"41C9",
			x"0000" when x"41CA",
			x"0000" when x"41CB",
			x"0000" when x"41CC",
			x"0000" when x"41CD",
			x"0000" when x"41CE",
			x"0000" when x"41CF",
			x"0000" when x"41D0",
			x"0000" when x"41D1",
			x"0000" when x"41D2",
			x"0000" when x"41D3",
			x"0000" when x"41D4",
			x"0000" when x"41D5",
			x"0000" when x"41D6",
			x"0000" when x"41D7",
			x"0000" when x"41D8",
			x"0000" when x"41D9",
			x"0000" when x"41DA",
			x"0000" when x"41DB",
			x"0000" when x"41DC",
			x"0000" when x"41DD",
			x"0000" when x"41DE",
			x"0000" when x"41DF",
			x"0000" when x"41E0",
			x"0000" when x"41E1",
			x"0000" when x"41E2",
			x"0000" when x"41E3",
			x"0000" when x"41E4",
			x"0000" when x"41E5",
			x"0000" when x"41E6",
			x"0000" when x"41E7",
			x"0000" when x"41E8",
			x"0000" when x"41E9",
			x"0000" when x"41EA",
			x"0000" when x"41EB",
			x"0000" when x"41EC",
			x"0000" when x"41ED",
			x"0000" when x"41EE",
			x"0000" when x"41EF",
			x"0000" when x"41F0",
			x"0000" when x"41F1",
			x"0000" when x"41F2",
			x"0000" when x"41F3",
			x"0000" when x"41F4",
			x"0000" when x"41F5",
			x"0000" when x"41F6",
			x"0000" when x"41F7",
			x"0000" when x"41F8",
			x"0000" when x"41F9",
			x"0000" when x"41FA",
			x"0000" when x"41FB",
			x"0000" when x"41FC",
			x"0000" when x"41FD",
			x"0000" when x"41FE",
			x"0000" when x"41FF",
			x"0000" when x"4200",
			x"0000" when x"4201",
			x"0000" when x"4202",
			x"0000" when x"4203",
			x"0000" when x"4204",
			x"0000" when x"4205",
			x"0000" when x"4206",
			x"0000" when x"4207",
			x"0000" when x"4208",
			x"0000" when x"4209",
			x"0000" when x"420A",
			x"0000" when x"420B",
			x"0000" when x"420C",
			x"0000" when x"420D",
			x"0000" when x"420E",
			x"0000" when x"420F",
			x"0000" when x"4210",
			x"0000" when x"4211",
			x"0000" when x"4212",
			x"0000" when x"4213",
			x"0000" when x"4214",
			x"0000" when x"4215",
			x"0000" when x"4216",
			x"0000" when x"4217",
			x"0000" when x"4218",
			x"0000" when x"4219",
			x"0000" when x"421A",
			x"0000" when x"421B",
			x"0000" when x"421C",
			x"0000" when x"421D",
			x"0000" when x"421E",
			x"0000" when x"421F",
			x"0000" when x"4220",
			x"0000" when x"4221",
			x"0000" when x"4222",
			x"0000" when x"4223",
			x"0000" when x"4224",
			x"0000" when x"4225",
			x"0000" when x"4226",
			x"0000" when x"4227",
			x"0000" when x"4228",
			x"0000" when x"4229",
			x"0000" when x"422A",
			x"0000" when x"422B",
			x"0000" when x"422C",
			x"0000" when x"422D",
			x"0000" when x"422E",
			x"0000" when x"422F",
			x"0000" when x"4230",
			x"0000" when x"4231",
			x"0000" when x"4232",
			x"0000" when x"4233",
			x"0000" when x"4234",
			x"0000" when x"4235",
			x"0000" when x"4236",
			x"0000" when x"4237",
			x"0000" when x"4238",
			x"0000" when x"4239",
			x"0000" when x"423A",
			x"0000" when x"423B",
			x"0000" when x"423C",
			x"0000" when x"423D",
			x"0000" when x"423E",
			x"0000" when x"423F",
			x"0000" when x"4240",
			x"0000" when x"4241",
			x"0000" when x"4242",
			x"0000" when x"4243",
			x"0000" when x"4244",
			x"0000" when x"4245",
			x"0000" when x"4246",
			x"0000" when x"4247",
			x"0000" when x"4248",
			x"0000" when x"4249",
			x"0000" when x"424A",
			x"0000" when x"424B",
			x"0000" when x"424C",
			x"0000" when x"424D",
			x"0000" when x"424E",
			x"0000" when x"424F",
			x"0000" when x"4250",
			x"0000" when x"4251",
			x"0000" when x"4252",
			x"0000" when x"4253",
			x"0000" when x"4254",
			x"0000" when x"4255",
			x"0000" when x"4256",
			x"0000" when x"4257",
			x"0000" when x"4258",
			x"0000" when x"4259",
			x"0000" when x"425A",
			x"0000" when x"425B",
			x"0000" when x"425C",
			x"0000" when x"425D",
			x"0000" when x"425E",
			x"0000" when x"425F",
			x"0000" when x"4260",
			x"0000" when x"4261",
			x"0000" when x"4262",
			x"0000" when x"4263",
			x"0000" when x"4264",
			x"0000" when x"4265",
			x"0000" when x"4266",
			x"0000" when x"4267",
			x"0000" when x"4268",
			x"0000" when x"4269",
			x"0000" when x"426A",
			x"0000" when x"426B",
			x"0000" when x"426C",
			x"0000" when x"426D",
			x"0000" when x"426E",
			x"0000" when x"426F",
			x"0000" when x"4270",
			x"0000" when x"4271",
			x"0000" when x"4272",
			x"0000" when x"4273",
			x"0000" when x"4274",
			x"0000" when x"4275",
			x"0000" when x"4276",
			x"0000" when x"4277",
			x"0000" when x"4278",
			x"0000" when x"4279",
			x"0000" when x"427A",
			x"0000" when x"427B",
			x"0000" when x"427C",
			x"0000" when x"427D",
			x"0000" when x"427E",
			x"0000" when x"427F",
			x"0000" when x"4280",
			x"0000" when x"4281",
			x"0000" when x"4282",
			x"0000" when x"4283",
			x"0000" when x"4284",
			x"0000" when x"4285",
			x"0000" when x"4286",
			x"0000" when x"4287",
			x"0000" when x"4288",
			x"0000" when x"4289",
			x"0000" when x"428A",
			x"0000" when x"428B",
			x"0000" when x"428C",
			x"0000" when x"428D",
			x"0000" when x"428E",
			x"0000" when x"428F",
			x"0000" when x"4290",
			x"0000" when x"4291",
			x"0000" when x"4292",
			x"0000" when x"4293",
			x"0000" when x"4294",
			x"0000" when x"4295",
			x"0000" when x"4296",
			x"0000" when x"4297",
			x"0000" when x"4298",
			x"0000" when x"4299",
			x"0000" when x"429A",
			x"0000" when x"429B",
			x"0000" when x"429C",
			x"0000" when x"429D",
			x"0000" when x"429E",
			x"0000" when x"429F",
			x"0000" when x"42A0",
			x"0000" when x"42A1",
			x"0000" when x"42A2",
			x"0000" when x"42A3",
			x"0000" when x"42A4",
			x"0000" when x"42A5",
			x"0000" when x"42A6",
			x"0000" when x"42A7",
			x"0000" when x"42A8",
			x"0000" when x"42A9",
			x"0000" when x"42AA",
			x"0000" when x"42AB",
			x"0000" when x"42AC",
			x"0000" when x"42AD",
			x"0000" when x"42AE",
			x"0000" when x"42AF",
			x"0000" when x"42B0",
			x"0000" when x"42B1",
			x"0000" when x"42B2",
			x"0000" when x"42B3",
			x"0000" when x"42B4",
			x"0000" when x"42B5",
			x"0000" when x"42B6",
			x"0000" when x"42B7",
			x"0000" when x"42B8",
			x"0000" when x"42B9",
			x"0000" when x"42BA",
			x"0000" when x"42BB",
			x"0000" when x"42BC",
			x"0000" when x"42BD",
			x"0000" when x"42BE",
			x"0000" when x"42BF",
			x"0000" when x"42C0",
			x"0000" when x"42C1",
			x"0000" when x"42C2",
			x"0000" when x"42C3",
			x"0000" when x"42C4",
			x"0000" when x"42C5",
			x"0000" when x"42C6",
			x"0000" when x"42C7",
			x"0000" when x"42C8",
			x"0000" when x"42C9",
			x"0000" when x"42CA",
			x"0000" when x"42CB",
			x"0000" when x"42CC",
			x"0000" when x"42CD",
			x"0000" when x"42CE",
			x"0000" when x"42CF",
			x"0000" when x"42D0",
			x"0000" when x"42D1",
			x"0000" when x"42D2",
			x"0000" when x"42D3",
			x"0000" when x"42D4",
			x"0000" when x"42D5",
			x"0000" when x"42D6",
			x"0000" when x"42D7",
			x"0000" when x"42D8",
			x"0000" when x"42D9",
			x"0000" when x"42DA",
			x"0000" when x"42DB",
			x"0000" when x"42DC",
			x"0000" when x"42DD",
			x"0000" when x"42DE",
			x"0000" when x"42DF",
			x"0000" when x"42E0",
			x"0000" when x"42E1",
			x"0000" when x"42E2",
			x"0000" when x"42E3",
			x"0000" when x"42E4",
			x"0000" when x"42E5",
			x"0000" when x"42E6",
			x"0000" when x"42E7",
			x"0000" when x"42E8",
			x"0000" when x"42E9",
			x"0000" when x"42EA",
			x"0000" when x"42EB",
			x"0000" when x"42EC",
			x"0000" when x"42ED",
			x"0000" when x"42EE",
			x"0000" when x"42EF",
			x"0000" when x"42F0",
			x"0000" when x"42F1",
			x"0000" when x"42F2",
			x"0000" when x"42F3",
			x"0000" when x"42F4",
			x"0000" when x"42F5",
			x"0000" when x"42F6",
			x"0000" when x"42F7",
			x"0000" when x"42F8",
			x"0000" when x"42F9",
			x"0000" when x"42FA",
			x"0000" when x"42FB",
			x"0000" when x"42FC",
			x"0000" when x"42FD",
			x"0000" when x"42FE",
			x"0000" when x"42FF",
			x"0000" when x"4300",
			x"0000" when x"4301",
			x"0000" when x"4302",
			x"0000" when x"4303",
			x"0000" when x"4304",
			x"0000" when x"4305",
			x"0000" when x"4306",
			x"0000" when x"4307",
			x"0000" when x"4308",
			x"0000" when x"4309",
			x"0000" when x"430A",
			x"0000" when x"430B",
			x"0000" when x"430C",
			x"0000" when x"430D",
			x"0000" when x"430E",
			x"0000" when x"430F",
			x"0000" when x"4310",
			x"0000" when x"4311",
			x"0000" when x"4312",
			x"0000" when x"4313",
			x"0000" when x"4314",
			x"0000" when x"4315",
			x"0000" when x"4316",
			x"0000" when x"4317",
			x"0000" when x"4318",
			x"0000" when x"4319",
			x"0000" when x"431A",
			x"0000" when x"431B",
			x"0000" when x"431C",
			x"0000" when x"431D",
			x"0000" when x"431E",
			x"0000" when x"431F",
			x"0000" when x"4320",
			x"0000" when x"4321",
			x"0000" when x"4322",
			x"0000" when x"4323",
			x"0000" when x"4324",
			x"0000" when x"4325",
			x"0000" when x"4326",
			x"0000" when x"4327",
			x"0000" when x"4328",
			x"0000" when x"4329",
			x"0000" when x"432A",
			x"0000" when x"432B",
			x"0000" when x"432C",
			x"0000" when x"432D",
			x"0000" when x"432E",
			x"0000" when x"432F",
			x"0000" when x"4330",
			x"0000" when x"4331",
			x"0000" when x"4332",
			x"0000" when x"4333",
			x"0000" when x"4334",
			x"0000" when x"4335",
			x"0000" when x"4336",
			x"0000" when x"4337",
			x"0000" when x"4338",
			x"0000" when x"4339",
			x"0000" when x"433A",
			x"0000" when x"433B",
			x"0000" when x"433C",
			x"0000" when x"433D",
			x"0000" when x"433E",
			x"0000" when x"433F",
			x"0000" when x"4340",
			x"0000" when x"4341",
			x"0000" when x"4342",
			x"0000" when x"4343",
			x"0000" when x"4344",
			x"0000" when x"4345",
			x"0000" when x"4346",
			x"0000" when x"4347",
			x"0000" when x"4348",
			x"0000" when x"4349",
			x"0000" when x"434A",
			x"0000" when x"434B",
			x"0000" when x"434C",
			x"0000" when x"434D",
			x"0000" when x"434E",
			x"0000" when x"434F",
			x"0000" when x"4350",
			x"0000" when x"4351",
			x"0000" when x"4352",
			x"0000" when x"4353",
			x"0000" when x"4354",
			x"0000" when x"4355",
			x"0000" when x"4356",
			x"0000" when x"4357",
			x"0000" when x"4358",
			x"0000" when x"4359",
			x"0000" when x"435A",
			x"0000" when x"435B",
			x"0000" when x"435C",
			x"0000" when x"435D",
			x"0000" when x"435E",
			x"0000" when x"435F",
			x"0000" when x"4360",
			x"0000" when x"4361",
			x"0000" when x"4362",
			x"0000" when x"4363",
			x"0000" when x"4364",
			x"0000" when x"4365",
			x"0000" when x"4366",
			x"0000" when x"4367",
			x"0000" when x"4368",
			x"0000" when x"4369",
			x"0000" when x"436A",
			x"0000" when x"436B",
			x"0000" when x"436C",
			x"0000" when x"436D",
			x"0000" when x"436E",
			x"0000" when x"436F",
			x"0000" when x"4370",
			x"0000" when x"4371",
			x"0000" when x"4372",
			x"0000" when x"4373",
			x"0000" when x"4374",
			x"0000" when x"4375",
			x"0000" when x"4376",
			x"0000" when x"4377",
			x"0000" when x"4378",
			x"0000" when x"4379",
			x"0000" when x"437A",
			x"0000" when x"437B",
			x"0000" when x"437C",
			x"0000" when x"437D",
			x"0000" when x"437E",
			x"0000" when x"437F",
			x"0000" when x"4380",
			x"0000" when x"4381",
			x"0000" when x"4382",
			x"0000" when x"4383",
			x"0000" when x"4384",
			x"0000" when x"4385",
			x"0000" when x"4386",
			x"0000" when x"4387",
			x"0000" when x"4388",
			x"0000" when x"4389",
			x"0000" when x"438A",
			x"0000" when x"438B",
			x"0000" when x"438C",
			x"0000" when x"438D",
			x"0000" when x"438E",
			x"0000" when x"438F",
			x"0000" when x"4390",
			x"0000" when x"4391",
			x"0000" when x"4392",
			x"0000" when x"4393",
			x"0000" when x"4394",
			x"0000" when x"4395",
			x"0000" when x"4396",
			x"0000" when x"4397",
			x"0000" when x"4398",
			x"0000" when x"4399",
			x"0000" when x"439A",
			x"0000" when x"439B",
			x"0000" when x"439C",
			x"0000" when x"439D",
			x"0000" when x"439E",
			x"0000" when x"439F",
			x"0000" when x"43A0",
			x"0000" when x"43A1",
			x"0000" when x"43A2",
			x"0000" when x"43A3",
			x"0000" when x"43A4",
			x"0000" when x"43A5",
			x"0000" when x"43A6",
			x"0000" when x"43A7",
			x"0000" when x"43A8",
			x"0000" when x"43A9",
			x"0000" when x"43AA",
			x"0000" when x"43AB",
			x"0000" when x"43AC",
			x"0000" when x"43AD",
			x"0000" when x"43AE",
			x"0000" when x"43AF",
			x"0000" when x"43B0",
			x"0000" when x"43B1",
			x"0000" when x"43B2",
			x"0000" when x"43B3",
			x"0000" when x"43B4",
			x"0000" when x"43B5",
			x"0000" when x"43B6",
			x"0000" when x"43B7",
			x"0000" when x"43B8",
			x"0000" when x"43B9",
			x"0000" when x"43BA",
			x"0000" when x"43BB",
			x"0000" when x"43BC",
			x"0000" when x"43BD",
			x"0000" when x"43BE",
			x"0000" when x"43BF",
			x"0000" when x"43C0",
			x"0000" when x"43C1",
			x"0000" when x"43C2",
			x"0000" when x"43C3",
			x"0000" when x"43C4",
			x"0000" when x"43C5",
			x"0000" when x"43C6",
			x"0000" when x"43C7",
			x"0000" when x"43C8",
			x"0000" when x"43C9",
			x"0000" when x"43CA",
			x"0000" when x"43CB",
			x"0000" when x"43CC",
			x"0000" when x"43CD",
			x"0000" when x"43CE",
			x"0000" when x"43CF",
			x"0000" when x"43D0",
			x"0000" when x"43D1",
			x"0000" when x"43D2",
			x"0000" when x"43D3",
			x"0000" when x"43D4",
			x"0000" when x"43D5",
			x"0000" when x"43D6",
			x"0000" when x"43D7",
			x"0000" when x"43D8",
			x"0000" when x"43D9",
			x"0000" when x"43DA",
			x"0000" when x"43DB",
			x"0000" when x"43DC",
			x"0000" when x"43DD",
			x"0000" when x"43DE",
			x"0000" when x"43DF",
			x"0000" when x"43E0",
			x"0000" when x"43E1",
			x"0000" when x"43E2",
			x"0000" when x"43E3",
			x"0000" when x"43E4",
			x"0000" when x"43E5",
			x"0000" when x"43E6",
			x"0000" when x"43E7",
			x"0000" when x"43E8",
			x"0000" when x"43E9",
			x"0000" when x"43EA",
			x"0000" when x"43EB",
			x"0000" when x"43EC",
			x"0000" when x"43ED",
			x"0000" when x"43EE",
			x"0000" when x"43EF",
			x"0000" when x"43F0",
			x"0000" when x"43F1",
			x"0000" when x"43F2",
			x"0000" when x"43F3",
			x"0000" when x"43F4",
			x"0000" when x"43F5",
			x"0000" when x"43F6",
			x"0000" when x"43F7",
			x"0000" when x"43F8",
			x"0000" when x"43F9",
			x"0000" when x"43FA",
			x"0000" when x"43FB",
			x"0000" when x"43FC",
			x"0000" when x"43FD",
			x"0000" when x"43FE",
			x"0000" when x"43FF",
			x"0000" when x"4400",
			x"0000" when x"4401",
			x"0000" when x"4402",
			x"0000" when x"4403",
			x"0000" when x"4404",
			x"0000" when x"4405",
			x"0000" when x"4406",
			x"0000" when x"4407",
			x"0000" when x"4408",
			x"0000" when x"4409",
			x"0000" when x"440A",
			x"0000" when x"440B",
			x"0000" when x"440C",
			x"0000" when x"440D",
			x"0000" when x"440E",
			x"0000" when x"440F",
			x"0000" when x"4410",
			x"0000" when x"4411",
			x"0000" when x"4412",
			x"0000" when x"4413",
			x"0000" when x"4414",
			x"0000" when x"4415",
			x"0000" when x"4416",
			x"0000" when x"4417",
			x"0000" when x"4418",
			x"0000" when x"4419",
			x"0000" when x"441A",
			x"0000" when x"441B",
			x"0000" when x"441C",
			x"0000" when x"441D",
			x"0000" when x"441E",
			x"0000" when x"441F",
			x"0000" when x"4420",
			x"0000" when x"4421",
			x"0000" when x"4422",
			x"0000" when x"4423",
			x"0000" when x"4424",
			x"0000" when x"4425",
			x"0000" when x"4426",
			x"0000" when x"4427",
			x"0000" when x"4428",
			x"0000" when x"4429",
			x"0000" when x"442A",
			x"0000" when x"442B",
			x"0000" when x"442C",
			x"0000" when x"442D",
			x"0000" when x"442E",
			x"0000" when x"442F",
			x"0000" when x"4430",
			x"0000" when x"4431",
			x"0000" when x"4432",
			x"0000" when x"4433",
			x"0000" when x"4434",
			x"0000" when x"4435",
			x"0000" when x"4436",
			x"0000" when x"4437",
			x"0000" when x"4438",
			x"0000" when x"4439",
			x"0000" when x"443A",
			x"0000" when x"443B",
			x"0000" when x"443C",
			x"0000" when x"443D",
			x"0000" when x"443E",
			x"0000" when x"443F",
			x"0000" when x"4440",
			x"0000" when x"4441",
			x"0000" when x"4442",
			x"0000" when x"4443",
			x"0000" when x"4444",
			x"0000" when x"4445",
			x"0000" when x"4446",
			x"0000" when x"4447",
			x"0000" when x"4448",
			x"0000" when x"4449",
			x"0000" when x"444A",
			x"0000" when x"444B",
			x"0000" when x"444C",
			x"0000" when x"444D",
			x"0000" when x"444E",
			x"0000" when x"444F",
			x"0000" when x"4450",
			x"0000" when x"4451",
			x"0000" when x"4452",
			x"0000" when x"4453",
			x"0000" when x"4454",
			x"0000" when x"4455",
			x"0000" when x"4456",
			x"0000" when x"4457",
			x"0000" when x"4458",
			x"0000" when x"4459",
			x"0000" when x"445A",
			x"0000" when x"445B",
			x"0000" when x"445C",
			x"0000" when x"445D",
			x"0000" when x"445E",
			x"0000" when x"445F",
			x"0000" when x"4460",
			x"0000" when x"4461",
			x"0000" when x"4462",
			x"0000" when x"4463",
			x"0000" when x"4464",
			x"0000" when x"4465",
			x"0000" when x"4466",
			x"0000" when x"4467",
			x"0000" when x"4468",
			x"0000" when x"4469",
			x"0000" when x"446A",
			x"0000" when x"446B",
			x"0000" when x"446C",
			x"0000" when x"446D",
			x"0000" when x"446E",
			x"0000" when x"446F",
			x"0000" when x"4470",
			x"0000" when x"4471",
			x"0000" when x"4472",
			x"0000" when x"4473",
			x"0000" when x"4474",
			x"0000" when x"4475",
			x"0000" when x"4476",
			x"0000" when x"4477",
			x"0000" when x"4478",
			x"0000" when x"4479",
			x"0000" when x"447A",
			x"0000" when x"447B",
			x"0000" when x"447C",
			x"0000" when x"447D",
			x"0000" when x"447E",
			x"0000" when x"447F",
			x"0000" when x"4480",
			x"0000" when x"4481",
			x"0000" when x"4482",
			x"0000" when x"4483",
			x"0000" when x"4484",
			x"0000" when x"4485",
			x"0000" when x"4486",
			x"0000" when x"4487",
			x"0000" when x"4488",
			x"0000" when x"4489",
			x"0000" when x"448A",
			x"0000" when x"448B",
			x"0000" when x"448C",
			x"0000" when x"448D",
			x"0000" when x"448E",
			x"0000" when x"448F",
			x"0000" when x"4490",
			x"0000" when x"4491",
			x"0000" when x"4492",
			x"0000" when x"4493",
			x"0000" when x"4494",
			x"0000" when x"4495",
			x"0000" when x"4496",
			x"0000" when x"4497",
			x"0000" when x"4498",
			x"0000" when x"4499",
			x"0000" when x"449A",
			x"0000" when x"449B",
			x"0000" when x"449C",
			x"0000" when x"449D",
			x"0000" when x"449E",
			x"0000" when x"449F",
			x"0000" when x"44A0",
			x"0000" when x"44A1",
			x"0000" when x"44A2",
			x"0000" when x"44A3",
			x"0000" when x"44A4",
			x"0000" when x"44A5",
			x"0000" when x"44A6",
			x"0000" when x"44A7",
			x"0000" when x"44A8",
			x"0000" when x"44A9",
			x"0000" when x"44AA",
			x"0000" when x"44AB",
			x"0000" when x"44AC",
			x"0000" when x"44AD",
			x"0000" when x"44AE",
			x"0000" when x"44AF",
			x"0000" when x"44B0",
			x"0000" when x"44B1",
			x"0000" when x"44B2",
			x"0000" when x"44B3",
			x"0000" when x"44B4",
			x"0000" when x"44B5",
			x"0000" when x"44B6",
			x"0000" when x"44B7",
			x"0000" when x"44B8",
			x"0000" when x"44B9",
			x"0000" when x"44BA",
			x"0000" when x"44BB",
			x"0000" when x"44BC",
			x"0000" when x"44BD",
			x"0000" when x"44BE",
			x"0000" when x"44BF",
			x"0000" when x"44C0",
			x"0000" when x"44C1",
			x"0000" when x"44C2",
			x"0000" when x"44C3",
			x"0000" when x"44C4",
			x"0000" when x"44C5",
			x"0000" when x"44C6",
			x"0000" when x"44C7",
			x"0000" when x"44C8",
			x"0000" when x"44C9",
			x"0000" when x"44CA",
			x"0000" when x"44CB",
			x"0000" when x"44CC",
			x"0000" when x"44CD",
			x"0000" when x"44CE",
			x"0000" when x"44CF",
			x"0000" when x"44D0",
			x"0000" when x"44D1",
			x"0000" when x"44D2",
			x"0000" when x"44D3",
			x"0000" when x"44D4",
			x"0000" when x"44D5",
			x"0000" when x"44D6",
			x"0000" when x"44D7",
			x"0000" when x"44D8",
			x"0000" when x"44D9",
			x"0000" when x"44DA",
			x"0000" when x"44DB",
			x"0000" when x"44DC",
			x"0000" when x"44DD",
			x"0000" when x"44DE",
			x"0000" when x"44DF",
			x"0000" when x"44E0",
			x"0000" when x"44E1",
			x"0000" when x"44E2",
			x"0000" when x"44E3",
			x"0000" when x"44E4",
			x"0000" when x"44E5",
			x"0000" when x"44E6",
			x"0000" when x"44E7",
			x"0000" when x"44E8",
			x"0000" when x"44E9",
			x"0000" when x"44EA",
			x"0000" when x"44EB",
			x"0000" when x"44EC",
			x"0000" when x"44ED",
			x"0000" when x"44EE",
			x"0000" when x"44EF",
			x"0000" when x"44F0",
			x"0000" when x"44F1",
			x"0000" when x"44F2",
			x"0000" when x"44F3",
			x"0000" when x"44F4",
			x"0000" when x"44F5",
			x"0000" when x"44F6",
			x"0000" when x"44F7",
			x"0000" when x"44F8",
			x"0000" when x"44F9",
			x"0000" when x"44FA",
			x"0000" when x"44FB",
			x"0000" when x"44FC",
			x"0000" when x"44FD",
			x"0000" when x"44FE",
			x"0000" when x"44FF",
			x"0000" when x"4500",
			x"0000" when x"4501",
			x"0000" when x"4502",
			x"0000" when x"4503",
			x"0000" when x"4504",
			x"0000" when x"4505",
			x"0000" when x"4506",
			x"0000" when x"4507",
			x"0000" when x"4508",
			x"0000" when x"4509",
			x"0000" when x"450A",
			x"0000" when x"450B",
			x"0000" when x"450C",
			x"0000" when x"450D",
			x"0000" when x"450E",
			x"0000" when x"450F",
			x"0000" when x"4510",
			x"0000" when x"4511",
			x"0000" when x"4512",
			x"0000" when x"4513",
			x"0000" when x"4514",
			x"0000" when x"4515",
			x"0000" when x"4516",
			x"0000" when x"4517",
			x"0000" when x"4518",
			x"0000" when x"4519",
			x"0000" when x"451A",
			x"0000" when x"451B",
			x"0000" when x"451C",
			x"0000" when x"451D",
			x"0000" when x"451E",
			x"0000" when x"451F",
			x"0000" when x"4520",
			x"0000" when x"4521",
			x"0000" when x"4522",
			x"0000" when x"4523",
			x"0000" when x"4524",
			x"0000" when x"4525",
			x"0000" when x"4526",
			x"0000" when x"4527",
			x"0000" when x"4528",
			x"0000" when x"4529",
			x"0000" when x"452A",
			x"0000" when x"452B",
			x"0000" when x"452C",
			x"0000" when x"452D",
			x"0000" when x"452E",
			x"0000" when x"452F",
			x"0000" when x"4530",
			x"0000" when x"4531",
			x"0000" when x"4532",
			x"0000" when x"4533",
			x"0000" when x"4534",
			x"0000" when x"4535",
			x"0000" when x"4536",
			x"0000" when x"4537",
			x"0000" when x"4538",
			x"0000" when x"4539",
			x"0000" when x"453A",
			x"0000" when x"453B",
			x"0000" when x"453C",
			x"0000" when x"453D",
			x"0000" when x"453E",
			x"0000" when x"453F",
			x"0000" when x"4540",
			x"0000" when x"4541",
			x"0000" when x"4542",
			x"0000" when x"4543",
			x"0000" when x"4544",
			x"0000" when x"4545",
			x"0000" when x"4546",
			x"0000" when x"4547",
			x"0000" when x"4548",
			x"0000" when x"4549",
			x"0000" when x"454A",
			x"0000" when x"454B",
			x"0000" when x"454C",
			x"0000" when x"454D",
			x"0000" when x"454E",
			x"0000" when x"454F",
			x"0000" when x"4550",
			x"0000" when x"4551",
			x"0000" when x"4552",
			x"0000" when x"4553",
			x"0000" when x"4554",
			x"0000" when x"4555",
			x"0000" when x"4556",
			x"0000" when x"4557",
			x"0000" when x"4558",
			x"0000" when x"4559",
			x"0000" when x"455A",
			x"0000" when x"455B",
			x"0000" when x"455C",
			x"0000" when x"455D",
			x"0000" when x"455E",
			x"0000" when x"455F",
			x"0000" when x"4560",
			x"0000" when x"4561",
			x"0000" when x"4562",
			x"0000" when x"4563",
			x"0000" when x"4564",
			x"0000" when x"4565",
			x"0000" when x"4566",
			x"0000" when x"4567",
			x"0000" when x"4568",
			x"0000" when x"4569",
			x"0000" when x"456A",
			x"0000" when x"456B",
			x"0000" when x"456C",
			x"0000" when x"456D",
			x"0000" when x"456E",
			x"0000" when x"456F",
			x"0000" when x"4570",
			x"0000" when x"4571",
			x"0000" when x"4572",
			x"0000" when x"4573",
			x"0000" when x"4574",
			x"0000" when x"4575",
			x"0000" when x"4576",
			x"0000" when x"4577",
			x"0000" when x"4578",
			x"0000" when x"4579",
			x"0000" when x"457A",
			x"0000" when x"457B",
			x"0000" when x"457C",
			x"0000" when x"457D",
			x"0000" when x"457E",
			x"0000" when x"457F",
			x"0000" when x"4580",
			x"0000" when x"4581",
			x"0000" when x"4582",
			x"0000" when x"4583",
			x"0000" when x"4584",
			x"0000" when x"4585",
			x"0000" when x"4586",
			x"0000" when x"4587",
			x"0000" when x"4588",
			x"0000" when x"4589",
			x"0000" when x"458A",
			x"0000" when x"458B",
			x"0000" when x"458C",
			x"0000" when x"458D",
			x"0000" when x"458E",
			x"0000" when x"458F",
			x"0000" when x"4590",
			x"0000" when x"4591",
			x"0000" when x"4592",
			x"0000" when x"4593",
			x"0000" when x"4594",
			x"0000" when x"4595",
			x"0000" when x"4596",
			x"0000" when x"4597",
			x"0000" when x"4598",
			x"0000" when x"4599",
			x"0000" when x"459A",
			x"0000" when x"459B",
			x"0000" when x"459C",
			x"0000" when x"459D",
			x"0000" when x"459E",
			x"0000" when x"459F",
			x"0000" when x"45A0",
			x"0000" when x"45A1",
			x"0000" when x"45A2",
			x"0000" when x"45A3",
			x"0000" when x"45A4",
			x"0000" when x"45A5",
			x"0000" when x"45A6",
			x"0000" when x"45A7",
			x"0000" when x"45A8",
			x"0000" when x"45A9",
			x"0000" when x"45AA",
			x"0000" when x"45AB",
			x"0000" when x"45AC",
			x"0000" when x"45AD",
			x"0000" when x"45AE",
			x"0000" when x"45AF",
			x"0000" when x"45B0",
			x"0000" when x"45B1",
			x"0000" when x"45B2",
			x"0000" when x"45B3",
			x"0000" when x"45B4",
			x"0000" when x"45B5",
			x"0000" when x"45B6",
			x"0000" when x"45B7",
			x"0000" when x"45B8",
			x"0000" when x"45B9",
			x"0000" when x"45BA",
			x"0000" when x"45BB",
			x"0000" when x"45BC",
			x"0000" when x"45BD",
			x"0000" when x"45BE",
			x"0000" when x"45BF",
			x"0000" when x"45C0",
			x"0000" when x"45C1",
			x"0000" when x"45C2",
			x"0000" when x"45C3",
			x"0000" when x"45C4",
			x"0000" when x"45C5",
			x"0000" when x"45C6",
			x"0000" when x"45C7",
			x"0000" when x"45C8",
			x"0000" when x"45C9",
			x"0000" when x"45CA",
			x"0000" when x"45CB",
			x"0000" when x"45CC",
			x"0000" when x"45CD",
			x"0000" when x"45CE",
			x"0000" when x"45CF",
			x"0000" when x"45D0",
			x"0000" when x"45D1",
			x"0000" when x"45D2",
			x"0000" when x"45D3",
			x"0000" when x"45D4",
			x"0000" when x"45D5",
			x"0000" when x"45D6",
			x"0000" when x"45D7",
			x"0000" when x"45D8",
			x"0000" when x"45D9",
			x"0000" when x"45DA",
			x"0000" when x"45DB",
			x"0000" when x"45DC",
			x"0000" when x"45DD",
			x"0000" when x"45DE",
			x"0000" when x"45DF",
			x"0000" when x"45E0",
			x"0000" when x"45E1",
			x"0000" when x"45E2",
			x"0000" when x"45E3",
			x"0000" when x"45E4",
			x"0000" when x"45E5",
			x"0000" when x"45E6",
			x"0000" when x"45E7",
			x"0000" when x"45E8",
			x"0000" when x"45E9",
			x"0000" when x"45EA",
			x"0000" when x"45EB",
			x"0000" when x"45EC",
			x"0000" when x"45ED",
			x"0000" when x"45EE",
			x"0000" when x"45EF",
			x"0000" when x"45F0",
			x"0000" when x"45F1",
			x"0000" when x"45F2",
			x"0000" when x"45F3",
			x"0000" when x"45F4",
			x"0000" when x"45F5",
			x"0000" when x"45F6",
			x"0000" when x"45F7",
			x"0000" when x"45F8",
			x"0000" when x"45F9",
			x"0000" when x"45FA",
			x"0000" when x"45FB",
			x"0000" when x"45FC",
			x"0000" when x"45FD",
			x"0000" when x"45FE",
			x"0000" when x"45FF",
			x"0000" when x"4600",
			x"0000" when x"4601",
			x"0000" when x"4602",
			x"0000" when x"4603",
			x"0000" when x"4604",
			x"0000" when x"4605",
			x"0000" when x"4606",
			x"0000" when x"4607",
			x"0000" when x"4608",
			x"0000" when x"4609",
			x"0000" when x"460A",
			x"0000" when x"460B",
			x"0000" when x"460C",
			x"0000" when x"460D",
			x"0000" when x"460E",
			x"0000" when x"460F",
			x"0000" when x"4610",
			x"0000" when x"4611",
			x"0000" when x"4612",
			x"0000" when x"4613",
			x"0000" when x"4614",
			x"0000" when x"4615",
			x"0000" when x"4616",
			x"0000" when x"4617",
			x"0000" when x"4618",
			x"0000" when x"4619",
			x"0000" when x"461A",
			x"0000" when x"461B",
			x"0000" when x"461C",
			x"0000" when x"461D",
			x"0000" when x"461E",
			x"0000" when x"461F",
			x"0000" when x"4620",
			x"0000" when x"4621",
			x"0000" when x"4622",
			x"0000" when x"4623",
			x"0000" when x"4624",
			x"0000" when x"4625",
			x"0000" when x"4626",
			x"0000" when x"4627",
			x"0000" when x"4628",
			x"0000" when x"4629",
			x"0000" when x"462A",
			x"0000" when x"462B",
			x"0000" when x"462C",
			x"0000" when x"462D",
			x"0000" when x"462E",
			x"0000" when x"462F",
			x"0000" when x"4630",
			x"0000" when x"4631",
			x"0000" when x"4632",
			x"0000" when x"4633",
			x"0000" when x"4634",
			x"0000" when x"4635",
			x"0000" when x"4636",
			x"0000" when x"4637",
			x"0000" when x"4638",
			x"0000" when x"4639",
			x"0000" when x"463A",
			x"0000" when x"463B",
			x"0000" when x"463C",
			x"0000" when x"463D",
			x"0000" when x"463E",
			x"0000" when x"463F",
			x"0000" when x"4640",
			x"0000" when x"4641",
			x"0000" when x"4642",
			x"0000" when x"4643",
			x"0000" when x"4644",
			x"0000" when x"4645",
			x"0000" when x"4646",
			x"0000" when x"4647",
			x"0000" when x"4648",
			x"0000" when x"4649",
			x"0000" when x"464A",
			x"0000" when x"464B",
			x"0000" when x"464C",
			x"0000" when x"464D",
			x"0000" when x"464E",
			x"0000" when x"464F",
			x"0000" when x"4650",
			x"0000" when x"4651",
			x"0000" when x"4652",
			x"0000" when x"4653",
			x"0000" when x"4654",
			x"0000" when x"4655",
			x"0000" when x"4656",
			x"0000" when x"4657",
			x"0000" when x"4658",
			x"0000" when x"4659",
			x"0000" when x"465A",
			x"0000" when x"465B",
			x"0000" when x"465C",
			x"0000" when x"465D",
			x"0000" when x"465E",
			x"0000" when x"465F",
			x"0000" when x"4660",
			x"0000" when x"4661",
			x"0000" when x"4662",
			x"0000" when x"4663",
			x"0000" when x"4664",
			x"0000" when x"4665",
			x"0000" when x"4666",
			x"0000" when x"4667",
			x"0000" when x"4668",
			x"0000" when x"4669",
			x"0000" when x"466A",
			x"0000" when x"466B",
			x"0000" when x"466C",
			x"0000" when x"466D",
			x"0000" when x"466E",
			x"0000" when x"466F",
			x"0000" when x"4670",
			x"0000" when x"4671",
			x"0000" when x"4672",
			x"0000" when x"4673",
			x"0000" when x"4674",
			x"0000" when x"4675",
			x"0000" when x"4676",
			x"0000" when x"4677",
			x"0000" when x"4678",
			x"0000" when x"4679",
			x"0000" when x"467A",
			x"0000" when x"467B",
			x"0000" when x"467C",
			x"0000" when x"467D",
			x"0000" when x"467E",
			x"0000" when x"467F",
			x"0000" when x"4680",
			x"0000" when x"4681",
			x"0000" when x"4682",
			x"0000" when x"4683",
			x"0000" when x"4684",
			x"0000" when x"4685",
			x"0000" when x"4686",
			x"0000" when x"4687",
			x"0000" when x"4688",
			x"0000" when x"4689",
			x"0000" when x"468A",
			x"0000" when x"468B",
			x"0000" when x"468C",
			x"0000" when x"468D",
			x"0000" when x"468E",
			x"0000" when x"468F",
			x"0000" when x"4690",
			x"0000" when x"4691",
			x"0000" when x"4692",
			x"0000" when x"4693",
			x"0000" when x"4694",
			x"0000" when x"4695",
			x"0000" when x"4696",
			x"0000" when x"4697",
			x"0000" when x"4698",
			x"0000" when x"4699",
			x"0000" when x"469A",
			x"0000" when x"469B",
			x"0000" when x"469C",
			x"0000" when x"469D",
			x"0000" when x"469E",
			x"0000" when x"469F",
			x"0000" when x"46A0",
			x"0000" when x"46A1",
			x"0000" when x"46A2",
			x"0000" when x"46A3",
			x"0000" when x"46A4",
			x"0000" when x"46A5",
			x"0000" when x"46A6",
			x"0000" when x"46A7",
			x"0000" when x"46A8",
			x"0000" when x"46A9",
			x"0000" when x"46AA",
			x"0000" when x"46AB",
			x"0000" when x"46AC",
			x"0000" when x"46AD",
			x"0000" when x"46AE",
			x"0000" when x"46AF",
			x"0000" when x"46B0",
			x"0000" when x"46B1",
			x"0000" when x"46B2",
			x"0000" when x"46B3",
			x"0000" when x"46B4",
			x"0000" when x"46B5",
			x"0000" when x"46B6",
			x"0000" when x"46B7",
			x"0000" when x"46B8",
			x"0000" when x"46B9",
			x"0000" when x"46BA",
			x"0000" when x"46BB",
			x"0000" when x"46BC",
			x"0000" when x"46BD",
			x"0000" when x"46BE",
			x"0000" when x"46BF",
			x"0000" when x"46C0",
			x"0000" when x"46C1",
			x"0000" when x"46C2",
			x"0000" when x"46C3",
			x"0000" when x"46C4",
			x"0000" when x"46C5",
			x"0000" when x"46C6",
			x"0000" when x"46C7",
			x"0000" when x"46C8",
			x"0000" when x"46C9",
			x"0000" when x"46CA",
			x"0000" when x"46CB",
			x"0000" when x"46CC",
			x"0000" when x"46CD",
			x"0000" when x"46CE",
			x"0000" when x"46CF",
			x"0000" when x"46D0",
			x"0000" when x"46D1",
			x"0000" when x"46D2",
			x"0000" when x"46D3",
			x"0000" when x"46D4",
			x"0000" when x"46D5",
			x"0000" when x"46D6",
			x"0000" when x"46D7",
			x"0000" when x"46D8",
			x"0000" when x"46D9",
			x"0000" when x"46DA",
			x"0000" when x"46DB",
			x"0000" when x"46DC",
			x"0000" when x"46DD",
			x"0000" when x"46DE",
			x"0000" when x"46DF",
			x"0000" when x"46E0",
			x"0000" when x"46E1",
			x"0000" when x"46E2",
			x"0000" when x"46E3",
			x"0000" when x"46E4",
			x"0000" when x"46E5",
			x"0000" when x"46E6",
			x"0000" when x"46E7",
			x"0000" when x"46E8",
			x"0000" when x"46E9",
			x"0000" when x"46EA",
			x"0000" when x"46EB",
			x"0000" when x"46EC",
			x"0000" when x"46ED",
			x"0000" when x"46EE",
			x"0000" when x"46EF",
			x"0000" when x"46F0",
			x"0000" when x"46F1",
			x"0000" when x"46F2",
			x"0000" when x"46F3",
			x"0000" when x"46F4",
			x"0000" when x"46F5",
			x"0000" when x"46F6",
			x"0000" when x"46F7",
			x"0000" when x"46F8",
			x"0000" when x"46F9",
			x"0000" when x"46FA",
			x"0000" when x"46FB",
			x"0000" when x"46FC",
			x"0000" when x"46FD",
			x"0000" when x"46FE",
			x"0000" when x"46FF",
			x"0000" when x"4700",
			x"0000" when x"4701",
			x"0000" when x"4702",
			x"0000" when x"4703",
			x"0000" when x"4704",
			x"0000" when x"4705",
			x"0000" when x"4706",
			x"0000" when x"4707",
			x"0000" when x"4708",
			x"0000" when x"4709",
			x"0000" when x"470A",
			x"0000" when x"470B",
			x"0000" when x"470C",
			x"0000" when x"470D",
			x"0000" when x"470E",
			x"0000" when x"470F",
			x"0000" when x"4710",
			x"0000" when x"4711",
			x"0000" when x"4712",
			x"0000" when x"4713",
			x"0000" when x"4714",
			x"0000" when x"4715",
			x"0000" when x"4716",
			x"0000" when x"4717",
			x"0000" when x"4718",
			x"0000" when x"4719",
			x"0000" when x"471A",
			x"0000" when x"471B",
			x"0000" when x"471C",
			x"0000" when x"471D",
			x"0000" when x"471E",
			x"0000" when x"471F",
			x"0000" when x"4720",
			x"0000" when x"4721",
			x"0000" when x"4722",
			x"0000" when x"4723",
			x"0000" when x"4724",
			x"0000" when x"4725",
			x"0000" when x"4726",
			x"0000" when x"4727",
			x"0000" when x"4728",
			x"0000" when x"4729",
			x"0000" when x"472A",
			x"0000" when x"472B",
			x"0000" when x"472C",
			x"0000" when x"472D",
			x"0000" when x"472E",
			x"0000" when x"472F",
			x"0000" when x"4730",
			x"0000" when x"4731",
			x"0000" when x"4732",
			x"0000" when x"4733",
			x"0000" when x"4734",
			x"0000" when x"4735",
			x"0000" when x"4736",
			x"0000" when x"4737",
			x"0000" when x"4738",
			x"0000" when x"4739",
			x"0000" when x"473A",
			x"0000" when x"473B",
			x"0000" when x"473C",
			x"0000" when x"473D",
			x"0000" when x"473E",
			x"0000" when x"473F",
			x"0000" when x"4740",
			x"0000" when x"4741",
			x"0000" when x"4742",
			x"0000" when x"4743",
			x"0000" when x"4744",
			x"0000" when x"4745",
			x"0000" when x"4746",
			x"0000" when x"4747",
			x"0000" when x"4748",
			x"0000" when x"4749",
			x"0000" when x"474A",
			x"0000" when x"474B",
			x"0000" when x"474C",
			x"0000" when x"474D",
			x"0000" when x"474E",
			x"0000" when x"474F",
			x"0000" when x"4750",
			x"0000" when x"4751",
			x"0000" when x"4752",
			x"0000" when x"4753",
			x"0000" when x"4754",
			x"0000" when x"4755",
			x"0000" when x"4756",
			x"0000" when x"4757",
			x"0000" when x"4758",
			x"0000" when x"4759",
			x"0000" when x"475A",
			x"0000" when x"475B",
			x"0000" when x"475C",
			x"0000" when x"475D",
			x"0000" when x"475E",
			x"0000" when x"475F",
			x"0000" when x"4760",
			x"0000" when x"4761",
			x"0000" when x"4762",
			x"0000" when x"4763",
			x"0000" when x"4764",
			x"0000" when x"4765",
			x"0000" when x"4766",
			x"0000" when x"4767",
			x"0000" when x"4768",
			x"0000" when x"4769",
			x"0000" when x"476A",
			x"0000" when x"476B",
			x"0000" when x"476C",
			x"0000" when x"476D",
			x"0000" when x"476E",
			x"0000" when x"476F",
			x"0000" when x"4770",
			x"0000" when x"4771",
			x"0000" when x"4772",
			x"0000" when x"4773",
			x"0000" when x"4774",
			x"0000" when x"4775",
			x"0000" when x"4776",
			x"0000" when x"4777",
			x"0000" when x"4778",
			x"0000" when x"4779",
			x"0000" when x"477A",
			x"0000" when x"477B",
			x"0000" when x"477C",
			x"0000" when x"477D",
			x"0000" when x"477E",
			x"0000" when x"477F",
			x"0000" when x"4780",
			x"0000" when x"4781",
			x"0000" when x"4782",
			x"0000" when x"4783",
			x"0000" when x"4784",
			x"0000" when x"4785",
			x"0000" when x"4786",
			x"0000" when x"4787",
			x"0000" when x"4788",
			x"0000" when x"4789",
			x"0000" when x"478A",
			x"0000" when x"478B",
			x"0000" when x"478C",
			x"0000" when x"478D",
			x"0000" when x"478E",
			x"0000" when x"478F",
			x"0000" when x"4790",
			x"0000" when x"4791",
			x"0000" when x"4792",
			x"0000" when x"4793",
			x"0000" when x"4794",
			x"0000" when x"4795",
			x"0000" when x"4796",
			x"0000" when x"4797",
			x"0000" when x"4798",
			x"0000" when x"4799",
			x"0000" when x"479A",
			x"0000" when x"479B",
			x"0000" when x"479C",
			x"0000" when x"479D",
			x"0000" when x"479E",
			x"0000" when x"479F",
			x"0000" when x"47A0",
			x"0000" when x"47A1",
			x"0000" when x"47A2",
			x"0000" when x"47A3",
			x"0000" when x"47A4",
			x"0000" when x"47A5",
			x"0000" when x"47A6",
			x"0000" when x"47A7",
			x"0000" when x"47A8",
			x"0000" when x"47A9",
			x"0000" when x"47AA",
			x"0000" when x"47AB",
			x"0000" when x"47AC",
			x"0000" when x"47AD",
			x"0000" when x"47AE",
			x"0000" when x"47AF",
			x"0000" when x"47B0",
			x"0000" when x"47B1",
			x"0000" when x"47B2",
			x"0000" when x"47B3",
			x"0000" when x"47B4",
			x"0000" when x"47B5",
			x"0000" when x"47B6",
			x"0000" when x"47B7",
			x"0000" when x"47B8",
			x"0000" when x"47B9",
			x"0000" when x"47BA",
			x"0000" when x"47BB",
			x"0000" when x"47BC",
			x"0000" when x"47BD",
			x"0000" when x"47BE",
			x"0000" when x"47BF",
			x"0000" when x"47C0",
			x"0000" when x"47C1",
			x"0000" when x"47C2",
			x"0000" when x"47C3",
			x"0000" when x"47C4",
			x"0000" when x"47C5",
			x"0000" when x"47C6",
			x"0000" when x"47C7",
			x"0000" when x"47C8",
			x"0000" when x"47C9",
			x"0000" when x"47CA",
			x"0000" when x"47CB",
			x"0000" when x"47CC",
			x"0000" when x"47CD",
			x"0000" when x"47CE",
			x"0000" when x"47CF",
			x"0000" when x"47D0",
			x"0000" when x"47D1",
			x"0000" when x"47D2",
			x"0000" when x"47D3",
			x"0000" when x"47D4",
			x"0000" when x"47D5",
			x"0000" when x"47D6",
			x"0000" when x"47D7",
			x"0000" when x"47D8",
			x"0000" when x"47D9",
			x"0000" when x"47DA",
			x"0000" when x"47DB",
			x"0000" when x"47DC",
			x"0000" when x"47DD",
			x"0000" when x"47DE",
			x"0000" when x"47DF",
			x"0000" when x"47E0",
			x"0000" when x"47E1",
			x"0000" when x"47E2",
			x"0000" when x"47E3",
			x"0000" when x"47E4",
			x"0000" when x"47E5",
			x"0000" when x"47E6",
			x"0000" when x"47E7",
			x"0000" when x"47E8",
			x"0000" when x"47E9",
			x"0000" when x"47EA",
			x"0000" when x"47EB",
			x"0000" when x"47EC",
			x"0000" when x"47ED",
			x"0000" when x"47EE",
			x"0000" when x"47EF",
			x"0000" when x"47F0",
			x"0000" when x"47F1",
			x"0000" when x"47F2",
			x"0000" when x"47F3",
			x"0000" when x"47F4",
			x"0000" when x"47F5",
			x"0000" when x"47F6",
			x"0000" when x"47F7",
			x"0000" when x"47F8",
			x"0000" when x"47F9",
			x"0000" when x"47FA",
			x"0000" when x"47FB",
			x"0000" when x"47FC",
			x"0000" when x"47FD",
			x"0000" when x"47FE",
			x"0000" when x"47FF",
			x"0000" when x"4800",
			x"0000" when x"4801",
			x"0000" when x"4802",
			x"0000" when x"4803",
			x"0000" when x"4804",
			x"0000" when x"4805",
			x"0000" when x"4806",
			x"0000" when x"4807",
			x"0000" when x"4808",
			x"0000" when x"4809",
			x"0000" when x"480A",
			x"0000" when x"480B",
			x"0000" when x"480C",
			x"0000" when x"480D",
			x"0000" when x"480E",
			x"0000" when x"480F",
			x"0000" when x"4810",
			x"0000" when x"4811",
			x"0000" when x"4812",
			x"0000" when x"4813",
			x"0000" when x"4814",
			x"0000" when x"4815",
			x"0000" when x"4816",
			x"0000" when x"4817",
			x"0000" when x"4818",
			x"0000" when x"4819",
			x"0000" when x"481A",
			x"0000" when x"481B",
			x"0000" when x"481C",
			x"0000" when x"481D",
			x"0000" when x"481E",
			x"0000" when x"481F",
			x"0000" when x"4820",
			x"0000" when x"4821",
			x"0000" when x"4822",
			x"0000" when x"4823",
			x"0000" when x"4824",
			x"0000" when x"4825",
			x"0000" when x"4826",
			x"0000" when x"4827",
			x"0000" when x"4828",
			x"0000" when x"4829",
			x"0000" when x"482A",
			x"0000" when x"482B",
			x"0000" when x"482C",
			x"0000" when x"482D",
			x"0000" when x"482E",
			x"0000" when x"482F",
			x"0000" when x"4830",
			x"0000" when x"4831",
			x"0000" when x"4832",
			x"0000" when x"4833",
			x"0000" when x"4834",
			x"0000" when x"4835",
			x"0000" when x"4836",
			x"0000" when x"4837",
			x"0000" when x"4838",
			x"0000" when x"4839",
			x"0000" when x"483A",
			x"0000" when x"483B",
			x"0000" when x"483C",
			x"0000" when x"483D",
			x"0000" when x"483E",
			x"0000" when x"483F",
			x"0000" when x"4840",
			x"0000" when x"4841",
			x"0000" when x"4842",
			x"0000" when x"4843",
			x"0000" when x"4844",
			x"0000" when x"4845",
			x"0000" when x"4846",
			x"0000" when x"4847",
			x"0000" when x"4848",
			x"0000" when x"4849",
			x"0000" when x"484A",
			x"0000" when x"484B",
			x"0000" when x"484C",
			x"0000" when x"484D",
			x"0000" when x"484E",
			x"0000" when x"484F",
			x"0000" when x"4850",
			x"0000" when x"4851",
			x"0000" when x"4852",
			x"0000" when x"4853",
			x"0000" when x"4854",
			x"0000" when x"4855",
			x"0000" when x"4856",
			x"0000" when x"4857",
			x"0000" when x"4858",
			x"0000" when x"4859",
			x"0000" when x"485A",
			x"0000" when x"485B",
			x"0000" when x"485C",
			x"0000" when x"485D",
			x"0000" when x"485E",
			x"0000" when x"485F",
			x"0000" when x"4860",
			x"0000" when x"4861",
			x"0000" when x"4862",
			x"0000" when x"4863",
			x"0000" when x"4864",
			x"0000" when x"4865",
			x"0000" when x"4866",
			x"0000" when x"4867",
			x"0000" when x"4868",
			x"0000" when x"4869",
			x"0000" when x"486A",
			x"0000" when x"486B",
			x"0000" when x"486C",
			x"0000" when x"486D",
			x"0000" when x"486E",
			x"0000" when x"486F",
			x"0000" when x"4870",
			x"0000" when x"4871",
			x"0000" when x"4872",
			x"0000" when x"4873",
			x"0000" when x"4874",
			x"0000" when x"4875",
			x"0000" when x"4876",
			x"0000" when x"4877",
			x"0000" when x"4878",
			x"0000" when x"4879",
			x"0000" when x"487A",
			x"0000" when x"487B",
			x"0000" when x"487C",
			x"0000" when x"487D",
			x"0000" when x"487E",
			x"0000" when x"487F",
			x"0000" when x"4880",
			x"0000" when x"4881",
			x"0000" when x"4882",
			x"0000" when x"4883",
			x"0000" when x"4884",
			x"0000" when x"4885",
			x"0000" when x"4886",
			x"0000" when x"4887",
			x"0000" when x"4888",
			x"0000" when x"4889",
			x"0000" when x"488A",
			x"0000" when x"488B",
			x"0000" when x"488C",
			x"0000" when x"488D",
			x"0000" when x"488E",
			x"0000" when x"488F",
			x"0000" when x"4890",
			x"0000" when x"4891",
			x"0000" when x"4892",
			x"0000" when x"4893",
			x"0000" when x"4894",
			x"0000" when x"4895",
			x"0000" when x"4896",
			x"0000" when x"4897",
			x"0000" when x"4898",
			x"0000" when x"4899",
			x"0000" when x"489A",
			x"0000" when x"489B",
			x"0000" when x"489C",
			x"0000" when x"489D",
			x"0000" when x"489E",
			x"0000" when x"489F",
			x"0000" when x"48A0",
			x"0000" when x"48A1",
			x"0000" when x"48A2",
			x"0000" when x"48A3",
			x"0000" when x"48A4",
			x"0000" when x"48A5",
			x"0000" when x"48A6",
			x"0000" when x"48A7",
			x"0000" when x"48A8",
			x"0000" when x"48A9",
			x"0000" when x"48AA",
			x"0000" when x"48AB",
			x"0000" when x"48AC",
			x"0000" when x"48AD",
			x"0000" when x"48AE",
			x"0000" when x"48AF",
			x"0000" when x"48B0",
			x"0000" when x"48B1",
			x"0000" when x"48B2",
			x"0000" when x"48B3",
			x"0000" when x"48B4",
			x"0000" when x"48B5",
			x"0000" when x"48B6",
			x"0000" when x"48B7",
			x"0000" when x"48B8",
			x"0000" when x"48B9",
			x"0000" when x"48BA",
			x"0000" when x"48BB",
			x"0000" when x"48BC",
			x"0000" when x"48BD",
			x"0000" when x"48BE",
			x"0000" when x"48BF",
			x"0000" when x"48C0",
			x"0000" when x"48C1",
			x"0000" when x"48C2",
			x"0000" when x"48C3",
			x"0000" when x"48C4",
			x"0000" when x"48C5",
			x"0000" when x"48C6",
			x"0000" when x"48C7",
			x"0000" when x"48C8",
			x"0000" when x"48C9",
			x"0000" when x"48CA",
			x"0000" when x"48CB",
			x"0000" when x"48CC",
			x"0000" when x"48CD",
			x"0000" when x"48CE",
			x"0000" when x"48CF",
			x"0000" when x"48D0",
			x"0000" when x"48D1",
			x"0000" when x"48D2",
			x"0000" when x"48D3",
			x"0000" when x"48D4",
			x"0000" when x"48D5",
			x"0000" when x"48D6",
			x"0000" when x"48D7",
			x"0000" when x"48D8",
			x"0000" when x"48D9",
			x"0000" when x"48DA",
			x"0000" when x"48DB",
			x"0000" when x"48DC",
			x"0000" when x"48DD",
			x"0000" when x"48DE",
			x"0000" when x"48DF",
			x"0000" when x"48E0",
			x"0000" when x"48E1",
			x"0000" when x"48E2",
			x"0000" when x"48E3",
			x"0000" when x"48E4",
			x"0000" when x"48E5",
			x"0000" when x"48E6",
			x"0000" when x"48E7",
			x"0000" when x"48E8",
			x"0000" when x"48E9",
			x"0000" when x"48EA",
			x"0000" when x"48EB",
			x"0000" when x"48EC",
			x"0000" when x"48ED",
			x"0000" when x"48EE",
			x"0000" when x"48EF",
			x"0000" when x"48F0",
			x"0000" when x"48F1",
			x"0000" when x"48F2",
			x"0000" when x"48F3",
			x"0000" when x"48F4",
			x"0000" when x"48F5",
			x"0000" when x"48F6",
			x"0000" when x"48F7",
			x"0000" when x"48F8",
			x"0000" when x"48F9",
			x"0000" when x"48FA",
			x"0000" when x"48FB",
			x"0000" when x"48FC",
			x"0000" when x"48FD",
			x"0000" when x"48FE",
			x"0000" when x"48FF",
			x"0000" when x"4900",
			x"0000" when x"4901",
			x"0000" when x"4902",
			x"0000" when x"4903",
			x"0000" when x"4904",
			x"0000" when x"4905",
			x"0000" when x"4906",
			x"0000" when x"4907",
			x"0000" when x"4908",
			x"0000" when x"4909",
			x"0000" when x"490A",
			x"0000" when x"490B",
			x"0000" when x"490C",
			x"0000" when x"490D",
			x"0000" when x"490E",
			x"0000" when x"490F",
			x"0000" when x"4910",
			x"0000" when x"4911",
			x"0000" when x"4912",
			x"0000" when x"4913",
			x"0000" when x"4914",
			x"0000" when x"4915",
			x"0000" when x"4916",
			x"0000" when x"4917",
			x"0000" when x"4918",
			x"0000" when x"4919",
			x"0000" when x"491A",
			x"0000" when x"491B",
			x"0000" when x"491C",
			x"0000" when x"491D",
			x"0000" when x"491E",
			x"0000" when x"491F",
			x"0000" when x"4920",
			x"0000" when x"4921",
			x"0000" when x"4922",
			x"0000" when x"4923",
			x"0000" when x"4924",
			x"0000" when x"4925",
			x"0000" when x"4926",
			x"0000" when x"4927",
			x"0000" when x"4928",
			x"0000" when x"4929",
			x"0000" when x"492A",
			x"0000" when x"492B",
			x"0000" when x"492C",
			x"0000" when x"492D",
			x"0000" when x"492E",
			x"0000" when x"492F",
			x"0000" when x"4930",
			x"0000" when x"4931",
			x"0000" when x"4932",
			x"0000" when x"4933",
			x"0000" when x"4934",
			x"0000" when x"4935",
			x"0000" when x"4936",
			x"0000" when x"4937",
			x"0000" when x"4938",
			x"0000" when x"4939",
			x"0000" when x"493A",
			x"0000" when x"493B",
			x"0000" when x"493C",
			x"0000" when x"493D",
			x"0000" when x"493E",
			x"0000" when x"493F",
			x"0000" when x"4940",
			x"0000" when x"4941",
			x"0000" when x"4942",
			x"0000" when x"4943",
			x"0000" when x"4944",
			x"0000" when x"4945",
			x"0000" when x"4946",
			x"0000" when x"4947",
			x"0000" when x"4948",
			x"0000" when x"4949",
			x"0000" when x"494A",
			x"0000" when x"494B",
			x"0000" when x"494C",
			x"0000" when x"494D",
			x"0000" when x"494E",
			x"0000" when x"494F",
			x"0000" when x"4950",
			x"0000" when x"4951",
			x"0000" when x"4952",
			x"0000" when x"4953",
			x"0000" when x"4954",
			x"0000" when x"4955",
			x"0000" when x"4956",
			x"0000" when x"4957",
			x"0000" when x"4958",
			x"0000" when x"4959",
			x"0000" when x"495A",
			x"0000" when x"495B",
			x"0000" when x"495C",
			x"0000" when x"495D",
			x"0000" when x"495E",
			x"0000" when x"495F",
			x"0000" when x"4960",
			x"0000" when x"4961",
			x"0000" when x"4962",
			x"0000" when x"4963",
			x"0000" when x"4964",
			x"0000" when x"4965",
			x"0000" when x"4966",
			x"0000" when x"4967",
			x"0000" when x"4968",
			x"0000" when x"4969",
			x"0000" when x"496A",
			x"0000" when x"496B",
			x"0000" when x"496C",
			x"0000" when x"496D",
			x"0000" when x"496E",
			x"0000" when x"496F",
			x"0000" when x"4970",
			x"0000" when x"4971",
			x"0000" when x"4972",
			x"0000" when x"4973",
			x"0000" when x"4974",
			x"0000" when x"4975",
			x"0000" when x"4976",
			x"0000" when x"4977",
			x"0000" when x"4978",
			x"0000" when x"4979",
			x"0000" when x"497A",
			x"0000" when x"497B",
			x"0000" when x"497C",
			x"0000" when x"497D",
			x"0000" when x"497E",
			x"0000" when x"497F",
			x"0000" when x"4980",
			x"0000" when x"4981",
			x"0000" when x"4982",
			x"0000" when x"4983",
			x"0000" when x"4984",
			x"0000" when x"4985",
			x"0000" when x"4986",
			x"0000" when x"4987",
			x"0000" when x"4988",
			x"0000" when x"4989",
			x"0000" when x"498A",
			x"0000" when x"498B",
			x"0000" when x"498C",
			x"0000" when x"498D",
			x"0000" when x"498E",
			x"0000" when x"498F",
			x"0000" when x"4990",
			x"0000" when x"4991",
			x"0000" when x"4992",
			x"0000" when x"4993",
			x"0000" when x"4994",
			x"0000" when x"4995",
			x"0000" when x"4996",
			x"0000" when x"4997",
			x"0000" when x"4998",
			x"0000" when x"4999",
			x"0000" when x"499A",
			x"0000" when x"499B",
			x"0000" when x"499C",
			x"0000" when x"499D",
			x"0000" when x"499E",
			x"0000" when x"499F",
			x"0000" when x"49A0",
			x"0000" when x"49A1",
			x"0000" when x"49A2",
			x"0000" when x"49A3",
			x"0000" when x"49A4",
			x"0000" when x"49A5",
			x"0000" when x"49A6",
			x"0000" when x"49A7",
			x"0000" when x"49A8",
			x"0000" when x"49A9",
			x"0000" when x"49AA",
			x"0000" when x"49AB",
			x"0000" when x"49AC",
			x"0000" when x"49AD",
			x"0000" when x"49AE",
			x"0000" when x"49AF",
			x"0000" when x"49B0",
			x"0000" when x"49B1",
			x"0000" when x"49B2",
			x"0000" when x"49B3",
			x"0000" when x"49B4",
			x"0000" when x"49B5",
			x"0000" when x"49B6",
			x"0000" when x"49B7",
			x"0000" when x"49B8",
			x"0000" when x"49B9",
			x"0000" when x"49BA",
			x"0000" when x"49BB",
			x"0000" when x"49BC",
			x"0000" when x"49BD",
			x"0000" when x"49BE",
			x"0000" when x"49BF",
			x"0000" when x"49C0",
			x"0000" when x"49C1",
			x"0000" when x"49C2",
			x"0000" when x"49C3",
			x"0000" when x"49C4",
			x"0000" when x"49C5",
			x"0000" when x"49C6",
			x"0000" when x"49C7",
			x"0000" when x"49C8",
			x"0000" when x"49C9",
			x"0000" when x"49CA",
			x"0000" when x"49CB",
			x"0000" when x"49CC",
			x"0000" when x"49CD",
			x"0000" when x"49CE",
			x"0000" when x"49CF",
			x"0000" when x"49D0",
			x"0000" when x"49D1",
			x"0000" when x"49D2",
			x"0000" when x"49D3",
			x"0000" when x"49D4",
			x"0000" when x"49D5",
			x"0000" when x"49D6",
			x"0000" when x"49D7",
			x"0000" when x"49D8",
			x"0000" when x"49D9",
			x"0000" when x"49DA",
			x"0000" when x"49DB",
			x"0000" when x"49DC",
			x"0000" when x"49DD",
			x"0000" when x"49DE",
			x"0000" when x"49DF",
			x"0000" when x"49E0",
			x"0000" when x"49E1",
			x"0000" when x"49E2",
			x"0000" when x"49E3",
			x"0000" when x"49E4",
			x"0000" when x"49E5",
			x"0000" when x"49E6",
			x"0000" when x"49E7",
			x"0000" when x"49E8",
			x"0000" when x"49E9",
			x"0000" when x"49EA",
			x"0000" when x"49EB",
			x"0000" when x"49EC",
			x"0000" when x"49ED",
			x"0000" when x"49EE",
			x"0000" when x"49EF",
			x"0000" when x"49F0",
			x"0000" when x"49F1",
			x"0000" when x"49F2",
			x"0000" when x"49F3",
			x"0000" when x"49F4",
			x"0000" when x"49F5",
			x"0000" when x"49F6",
			x"0000" when x"49F7",
			x"0000" when x"49F8",
			x"0000" when x"49F9",
			x"0000" when x"49FA",
			x"0000" when x"49FB",
			x"0000" when x"49FC",
			x"0000" when x"49FD",
			x"0000" when x"49FE",
			x"0000" when x"49FF",
			x"0000" when x"4A00",
			x"0000" when x"4A01",
			x"0000" when x"4A02",
			x"0000" when x"4A03",
			x"0000" when x"4A04",
			x"0000" when x"4A05",
			x"0000" when x"4A06",
			x"0000" when x"4A07",
			x"0000" when x"4A08",
			x"0000" when x"4A09",
			x"0000" when x"4A0A",
			x"0000" when x"4A0B",
			x"0000" when x"4A0C",
			x"0000" when x"4A0D",
			x"0000" when x"4A0E",
			x"0000" when x"4A0F",
			x"0000" when x"4A10",
			x"0000" when x"4A11",
			x"0000" when x"4A12",
			x"0000" when x"4A13",
			x"0000" when x"4A14",
			x"0000" when x"4A15",
			x"0000" when x"4A16",
			x"0000" when x"4A17",
			x"0000" when x"4A18",
			x"0000" when x"4A19",
			x"0000" when x"4A1A",
			x"0000" when x"4A1B",
			x"0000" when x"4A1C",
			x"0000" when x"4A1D",
			x"0000" when x"4A1E",
			x"0000" when x"4A1F",
			x"0000" when x"4A20",
			x"0000" when x"4A21",
			x"0000" when x"4A22",
			x"0000" when x"4A23",
			x"0000" when x"4A24",
			x"0000" when x"4A25",
			x"0000" when x"4A26",
			x"0000" when x"4A27",
			x"0000" when x"4A28",
			x"0000" when x"4A29",
			x"0000" when x"4A2A",
			x"0000" when x"4A2B",
			x"0000" when x"4A2C",
			x"0000" when x"4A2D",
			x"0000" when x"4A2E",
			x"0000" when x"4A2F",
			x"0000" when x"4A30",
			x"0000" when x"4A31",
			x"0000" when x"4A32",
			x"0000" when x"4A33",
			x"0000" when x"4A34",
			x"0000" when x"4A35",
			x"0000" when x"4A36",
			x"0000" when x"4A37",
			x"0000" when x"4A38",
			x"0000" when x"4A39",
			x"0000" when x"4A3A",
			x"0000" when x"4A3B",
			x"0000" when x"4A3C",
			x"0000" when x"4A3D",
			x"0000" when x"4A3E",
			x"0000" when x"4A3F",
			x"0000" when x"4A40",
			x"0000" when x"4A41",
			x"0000" when x"4A42",
			x"0000" when x"4A43",
			x"0000" when x"4A44",
			x"0000" when x"4A45",
			x"0000" when x"4A46",
			x"0000" when x"4A47",
			x"0000" when x"4A48",
			x"0000" when x"4A49",
			x"0000" when x"4A4A",
			x"0000" when x"4A4B",
			x"0000" when x"4A4C",
			x"0000" when x"4A4D",
			x"0000" when x"4A4E",
			x"0000" when x"4A4F",
			x"0000" when x"4A50",
			x"0000" when x"4A51",
			x"0000" when x"4A52",
			x"0000" when x"4A53",
			x"0000" when x"4A54",
			x"0000" when x"4A55",
			x"0000" when x"4A56",
			x"0000" when x"4A57",
			x"0000" when x"4A58",
			x"0000" when x"4A59",
			x"0000" when x"4A5A",
			x"0000" when x"4A5B",
			x"0000" when x"4A5C",
			x"0000" when x"4A5D",
			x"0000" when x"4A5E",
			x"0000" when x"4A5F",
			x"0000" when x"4A60",
			x"0000" when x"4A61",
			x"0000" when x"4A62",
			x"0000" when x"4A63",
			x"0000" when x"4A64",
			x"0000" when x"4A65",
			x"0000" when x"4A66",
			x"0000" when x"4A67",
			x"0000" when x"4A68",
			x"0000" when x"4A69",
			x"0000" when x"4A6A",
			x"0000" when x"4A6B",
			x"0000" when x"4A6C",
			x"0000" when x"4A6D",
			x"0000" when x"4A6E",
			x"0000" when x"4A6F",
			x"0000" when x"4A70",
			x"0000" when x"4A71",
			x"0000" when x"4A72",
			x"0000" when x"4A73",
			x"0000" when x"4A74",
			x"0000" when x"4A75",
			x"0000" when x"4A76",
			x"0000" when x"4A77",
			x"0000" when x"4A78",
			x"0000" when x"4A79",
			x"0000" when x"4A7A",
			x"0000" when x"4A7B",
			x"0000" when x"4A7C",
			x"0000" when x"4A7D",
			x"0000" when x"4A7E",
			x"0000" when x"4A7F",
			x"0000" when x"4A80",
			x"0000" when x"4A81",
			x"0000" when x"4A82",
			x"0000" when x"4A83",
			x"0000" when x"4A84",
			x"0000" when x"4A85",
			x"0000" when x"4A86",
			x"0000" when x"4A87",
			x"0000" when x"4A88",
			x"0000" when x"4A89",
			x"0000" when x"4A8A",
			x"0000" when x"4A8B",
			x"0000" when x"4A8C",
			x"0000" when x"4A8D",
			x"0000" when x"4A8E",
			x"0000" when x"4A8F",
			x"0000" when x"4A90",
			x"0000" when x"4A91",
			x"0000" when x"4A92",
			x"0000" when x"4A93",
			x"0000" when x"4A94",
			x"0000" when x"4A95",
			x"0000" when x"4A96",
			x"0000" when x"4A97",
			x"0000" when x"4A98",
			x"0000" when x"4A99",
			x"0000" when x"4A9A",
			x"0000" when x"4A9B",
			x"0000" when x"4A9C",
			x"0000" when x"4A9D",
			x"0000" when x"4A9E",
			x"0000" when x"4A9F",
			x"0000" when x"4AA0",
			x"0000" when x"4AA1",
			x"0000" when x"4AA2",
			x"0000" when x"4AA3",
			x"0000" when x"4AA4",
			x"0000" when x"4AA5",
			x"0000" when x"4AA6",
			x"0000" when x"4AA7",
			x"0000" when x"4AA8",
			x"0000" when x"4AA9",
			x"0000" when x"4AAA",
			x"0000" when x"4AAB",
			x"0000" when x"4AAC",
			x"0000" when x"4AAD",
			x"0000" when x"4AAE",
			x"0000" when x"4AAF",
			x"0000" when x"4AB0",
			x"0000" when x"4AB1",
			x"0000" when x"4AB2",
			x"0000" when x"4AB3",
			x"0000" when x"4AB4",
			x"0000" when x"4AB5",
			x"0000" when x"4AB6",
			x"0000" when x"4AB7",
			x"0000" when x"4AB8",
			x"0000" when x"4AB9",
			x"0000" when x"4ABA",
			x"0000" when x"4ABB",
			x"0000" when x"4ABC",
			x"0000" when x"4ABD",
			x"0000" when x"4ABE",
			x"0000" when x"4ABF",
			x"0000" when x"4AC0",
			x"0000" when x"4AC1",
			x"0000" when x"4AC2",
			x"0000" when x"4AC3",
			x"0000" when x"4AC4",
			x"0000" when x"4AC5",
			x"0000" when x"4AC6",
			x"0000" when x"4AC7",
			x"0000" when x"4AC8",
			x"0000" when x"4AC9",
			x"0000" when x"4ACA",
			x"0000" when x"4ACB",
			x"0000" when x"4ACC",
			x"0000" when x"4ACD",
			x"0000" when x"4ACE",
			x"0000" when x"4ACF",
			x"0000" when x"4AD0",
			x"0000" when x"4AD1",
			x"0000" when x"4AD2",
			x"0000" when x"4AD3",
			x"0000" when x"4AD4",
			x"0000" when x"4AD5",
			x"0000" when x"4AD6",
			x"0000" when x"4AD7",
			x"0000" when x"4AD8",
			x"0000" when x"4AD9",
			x"0000" when x"4ADA",
			x"0000" when x"4ADB",
			x"0000" when x"4ADC",
			x"0000" when x"4ADD",
			x"0000" when x"4ADE",
			x"0000" when x"4ADF",
			x"0000" when x"4AE0",
			x"0000" when x"4AE1",
			x"0000" when x"4AE2",
			x"0000" when x"4AE3",
			x"0000" when x"4AE4",
			x"0000" when x"4AE5",
			x"0000" when x"4AE6",
			x"0000" when x"4AE7",
			x"0000" when x"4AE8",
			x"0000" when x"4AE9",
			x"0000" when x"4AEA",
			x"0000" when x"4AEB",
			x"0000" when x"4AEC",
			x"0000" when x"4AED",
			x"0000" when x"4AEE",
			x"0000" when x"4AEF",
			x"0000" when x"4AF0",
			x"0000" when x"4AF1",
			x"0000" when x"4AF2",
			x"0000" when x"4AF3",
			x"0000" when x"4AF4",
			x"0000" when x"4AF5",
			x"0000" when x"4AF6",
			x"0000" when x"4AF7",
			x"0000" when x"4AF8",
			x"0000" when x"4AF9",
			x"0000" when x"4AFA",
			x"0000" when x"4AFB",
			x"0000" when x"4AFC",
			x"0000" when x"4AFD",
			x"0000" when x"4AFE",
			x"0000" when x"4AFF",
			x"0000" when x"4B00",
			x"0000" when x"4B01",
			x"0000" when x"4B02",
			x"0000" when x"4B03",
			x"0000" when x"4B04",
			x"0000" when x"4B05",
			x"0000" when x"4B06",
			x"0000" when x"4B07",
			x"0000" when x"4B08",
			x"0000" when x"4B09",
			x"0000" when x"4B0A",
			x"0000" when x"4B0B",
			x"0000" when x"4B0C",
			x"0000" when x"4B0D",
			x"0000" when x"4B0E",
			x"0000" when x"4B0F",
			x"0000" when x"4B10",
			x"0000" when x"4B11",
			x"0000" when x"4B12",
			x"0000" when x"4B13",
			x"0000" when x"4B14",
			x"0000" when x"4B15",
			x"0000" when x"4B16",
			x"0000" when x"4B17",
			x"0000" when x"4B18",
			x"0000" when x"4B19",
			x"0000" when x"4B1A",
			x"0000" when x"4B1B",
			x"0000" when x"4B1C",
			x"0000" when x"4B1D",
			x"0000" when x"4B1E",
			x"0000" when x"4B1F",
			x"0000" when x"4B20",
			x"0000" when x"4B21",
			x"0000" when x"4B22",
			x"0000" when x"4B23",
			x"0000" when x"4B24",
			x"0000" when x"4B25",
			x"0000" when x"4B26",
			x"0000" when x"4B27",
			x"0000" when x"4B28",
			x"0000" when x"4B29",
			x"0000" when x"4B2A",
			x"0000" when x"4B2B",
			x"0000" when x"4B2C",
			x"0000" when x"4B2D",
			x"0000" when x"4B2E",
			x"0000" when x"4B2F",
			x"0000" when x"4B30",
			x"0000" when x"4B31",
			x"0000" when x"4B32",
			x"0000" when x"4B33",
			x"0000" when x"4B34",
			x"0000" when x"4B35",
			x"0000" when x"4B36",
			x"0000" when x"4B37",
			x"0000" when x"4B38",
			x"0000" when x"4B39",
			x"0000" when x"4B3A",
			x"0000" when x"4B3B",
			x"0000" when x"4B3C",
			x"0000" when x"4B3D",
			x"0000" when x"4B3E",
			x"0000" when x"4B3F",
			x"0000" when x"4B40",
			x"0000" when x"4B41",
			x"0000" when x"4B42",
			x"0000" when x"4B43",
			x"0000" when x"4B44",
			x"0000" when x"4B45",
			x"0000" when x"4B46",
			x"0000" when x"4B47",
			x"0000" when x"4B48",
			x"0000" when x"4B49",
			x"0000" when x"4B4A",
			x"0000" when x"4B4B",
			x"0000" when x"4B4C",
			x"0000" when x"4B4D",
			x"0000" when x"4B4E",
			x"0000" when x"4B4F",
			x"0000" when x"4B50",
			x"0000" when x"4B51",
			x"0000" when x"4B52",
			x"0000" when x"4B53",
			x"0000" when x"4B54",
			x"0000" when x"4B55",
			x"0000" when x"4B56",
			x"0000" when x"4B57",
			x"0000" when x"4B58",
			x"0000" when x"4B59",
			x"0000" when x"4B5A",
			x"0000" when x"4B5B",
			x"0000" when x"4B5C",
			x"0000" when x"4B5D",
			x"0000" when x"4B5E",
			x"0000" when x"4B5F",
			x"0000" when x"4B60",
			x"0000" when x"4B61",
			x"0000" when x"4B62",
			x"0000" when x"4B63",
			x"0000" when x"4B64",
			x"0000" when x"4B65",
			x"0000" when x"4B66",
			x"0000" when x"4B67",
			x"0000" when x"4B68",
			x"0000" when x"4B69",
			x"0000" when x"4B6A",
			x"0000" when x"4B6B",
			x"0000" when x"4B6C",
			x"0000" when x"4B6D",
			x"0000" when x"4B6E",
			x"0000" when x"4B6F",
			x"0000" when x"4B70",
			x"0000" when x"4B71",
			x"0000" when x"4B72",
			x"0000" when x"4B73",
			x"0000" when x"4B74",
			x"0000" when x"4B75",
			x"0000" when x"4B76",
			x"0000" when x"4B77",
			x"0000" when x"4B78",
			x"0000" when x"4B79",
			x"0000" when x"4B7A",
			x"0000" when x"4B7B",
			x"0000" when x"4B7C",
			x"0000" when x"4B7D",
			x"0000" when x"4B7E",
			x"0000" when x"4B7F",
			x"0000" when x"4B80",
			x"0000" when x"4B81",
			x"0000" when x"4B82",
			x"0000" when x"4B83",
			x"0000" when x"4B84",
			x"0000" when x"4B85",
			x"0000" when x"4B86",
			x"0000" when x"4B87",
			x"0000" when x"4B88",
			x"0000" when x"4B89",
			x"0000" when x"4B8A",
			x"0000" when x"4B8B",
			x"0000" when x"4B8C",
			x"0000" when x"4B8D",
			x"0000" when x"4B8E",
			x"0000" when x"4B8F",
			x"0000" when x"4B90",
			x"0000" when x"4B91",
			x"0000" when x"4B92",
			x"0000" when x"4B93",
			x"0000" when x"4B94",
			x"0000" when x"4B95",
			x"0000" when x"4B96",
			x"0000" when x"4B97",
			x"0000" when x"4B98",
			x"0000" when x"4B99",
			x"0000" when x"4B9A",
			x"0000" when x"4B9B",
			x"0000" when x"4B9C",
			x"0000" when x"4B9D",
			x"0000" when x"4B9E",
			x"0000" when x"4B9F",
			x"0000" when x"4BA0",
			x"0000" when x"4BA1",
			x"0000" when x"4BA2",
			x"0000" when x"4BA3",
			x"0000" when x"4BA4",
			x"0000" when x"4BA5",
			x"0000" when x"4BA6",
			x"0000" when x"4BA7",
			x"0000" when x"4BA8",
			x"0000" when x"4BA9",
			x"0000" when x"4BAA",
			x"0000" when x"4BAB",
			x"0000" when x"4BAC",
			x"0000" when x"4BAD",
			x"0000" when x"4BAE",
			x"0000" when x"4BAF",
			x"0000" when x"4BB0",
			x"0000" when x"4BB1",
			x"0000" when x"4BB2",
			x"0000" when x"4BB3",
			x"0000" when x"4BB4",
			x"0000" when x"4BB5",
			x"0000" when x"4BB6",
			x"0000" when x"4BB7",
			x"0000" when x"4BB8",
			x"0000" when x"4BB9",
			x"0000" when x"4BBA",
			x"0000" when x"4BBB",
			x"0000" when x"4BBC",
			x"0000" when x"4BBD",
			x"0000" when x"4BBE",
			x"0000" when x"4BBF",
			x"0000" when x"4BC0",
			x"0000" when x"4BC1",
			x"0000" when x"4BC2",
			x"0000" when x"4BC3",
			x"0000" when x"4BC4",
			x"0000" when x"4BC5",
			x"0000" when x"4BC6",
			x"0000" when x"4BC7",
			x"0000" when x"4BC8",
			x"0000" when x"4BC9",
			x"0000" when x"4BCA",
			x"0000" when x"4BCB",
			x"0000" when x"4BCC",
			x"0000" when x"4BCD",
			x"0000" when x"4BCE",
			x"0000" when x"4BCF",
			x"0000" when x"4BD0",
			x"0000" when x"4BD1",
			x"0000" when x"4BD2",
			x"0000" when x"4BD3",
			x"0000" when x"4BD4",
			x"0000" when x"4BD5",
			x"0000" when x"4BD6",
			x"0000" when x"4BD7",
			x"0000" when x"4BD8",
			x"0000" when x"4BD9",
			x"0000" when x"4BDA",
			x"0000" when x"4BDB",
			x"0000" when x"4BDC",
			x"0000" when x"4BDD",
			x"0000" when x"4BDE",
			x"0000" when x"4BDF",
			x"0000" when x"4BE0",
			x"0000" when x"4BE1",
			x"0000" when x"4BE2",
			x"0000" when x"4BE3",
			x"0000" when x"4BE4",
			x"0000" when x"4BE5",
			x"0000" when x"4BE6",
			x"0000" when x"4BE7",
			x"0000" when x"4BE8",
			x"0000" when x"4BE9",
			x"0000" when x"4BEA",
			x"0000" when x"4BEB",
			x"0000" when x"4BEC",
			x"0000" when x"4BED",
			x"0000" when x"4BEE",
			x"0000" when x"4BEF",
			x"0000" when x"4BF0",
			x"0000" when x"4BF1",
			x"0000" when x"4BF2",
			x"0000" when x"4BF3",
			x"0000" when x"4BF4",
			x"0000" when x"4BF5",
			x"0000" when x"4BF6",
			x"0000" when x"4BF7",
			x"0000" when x"4BF8",
			x"0000" when x"4BF9",
			x"0000" when x"4BFA",
			x"0000" when x"4BFB",
			x"0000" when x"4BFC",
			x"0000" when x"4BFD",
			x"0000" when x"4BFE",
			x"0000" when x"4BFF",
			x"0000" when x"4C00",
			x"0000" when x"4C01",
			x"0000" when x"4C02",
			x"0000" when x"4C03",
			x"0000" when x"4C04",
			x"0000" when x"4C05",
			x"0000" when x"4C06",
			x"0000" when x"4C07",
			x"0000" when x"4C08",
			x"0000" when x"4C09",
			x"0000" when x"4C0A",
			x"0000" when x"4C0B",
			x"0000" when x"4C0C",
			x"0000" when x"4C0D",
			x"0000" when x"4C0E",
			x"0000" when x"4C0F",
			x"0000" when x"4C10",
			x"0000" when x"4C11",
			x"0000" when x"4C12",
			x"0000" when x"4C13",
			x"0000" when x"4C14",
			x"0000" when x"4C15",
			x"0000" when x"4C16",
			x"0000" when x"4C17",
			x"0000" when x"4C18",
			x"0000" when x"4C19",
			x"0000" when x"4C1A",
			x"0000" when x"4C1B",
			x"0000" when x"4C1C",
			x"0000" when x"4C1D",
			x"0000" when x"4C1E",
			x"0000" when x"4C1F",
			x"0000" when x"4C20",
			x"0000" when x"4C21",
			x"0000" when x"4C22",
			x"0000" when x"4C23",
			x"0000" when x"4C24",
			x"0000" when x"4C25",
			x"0000" when x"4C26",
			x"0000" when x"4C27",
			x"0000" when x"4C28",
			x"0000" when x"4C29",
			x"0000" when x"4C2A",
			x"0000" when x"4C2B",
			x"0000" when x"4C2C",
			x"0000" when x"4C2D",
			x"0000" when x"4C2E",
			x"0000" when x"4C2F",
			x"0000" when x"4C30",
			x"0000" when x"4C31",
			x"0000" when x"4C32",
			x"0000" when x"4C33",
			x"0000" when x"4C34",
			x"0000" when x"4C35",
			x"0000" when x"4C36",
			x"0000" when x"4C37",
			x"0000" when x"4C38",
			x"0000" when x"4C39",
			x"0000" when x"4C3A",
			x"0000" when x"4C3B",
			x"0000" when x"4C3C",
			x"0000" when x"4C3D",
			x"0000" when x"4C3E",
			x"0000" when x"4C3F",
			x"0000" when x"4C40",
			x"0000" when x"4C41",
			x"0000" when x"4C42",
			x"0000" when x"4C43",
			x"0000" when x"4C44",
			x"0000" when x"4C45",
			x"0000" when x"4C46",
			x"0000" when x"4C47",
			x"0000" when x"4C48",
			x"0000" when x"4C49",
			x"0000" when x"4C4A",
			x"0000" when x"4C4B",
			x"0000" when x"4C4C",
			x"0000" when x"4C4D",
			x"0000" when x"4C4E",
			x"0000" when x"4C4F",
			x"0000" when x"4C50",
			x"0000" when x"4C51",
			x"0000" when x"4C52",
			x"0000" when x"4C53",
			x"0000" when x"4C54",
			x"0000" when x"4C55",
			x"0000" when x"4C56",
			x"0000" when x"4C57",
			x"0000" when x"4C58",
			x"0000" when x"4C59",
			x"0000" when x"4C5A",
			x"0000" when x"4C5B",
			x"0000" when x"4C5C",
			x"0000" when x"4C5D",
			x"0000" when x"4C5E",
			x"0000" when x"4C5F",
			x"0000" when x"4C60",
			x"0000" when x"4C61",
			x"0000" when x"4C62",
			x"0000" when x"4C63",
			x"0000" when x"4C64",
			x"0000" when x"4C65",
			x"0000" when x"4C66",
			x"0000" when x"4C67",
			x"0000" when x"4C68",
			x"0000" when x"4C69",
			x"0000" when x"4C6A",
			x"0000" when x"4C6B",
			x"0000" when x"4C6C",
			x"0000" when x"4C6D",
			x"0000" when x"4C6E",
			x"0000" when x"4C6F",
			x"0000" when x"4C70",
			x"0000" when x"4C71",
			x"0000" when x"4C72",
			x"0000" when x"4C73",
			x"0000" when x"4C74",
			x"0000" when x"4C75",
			x"0000" when x"4C76",
			x"0000" when x"4C77",
			x"0000" when x"4C78",
			x"0000" when x"4C79",
			x"0000" when x"4C7A",
			x"0000" when x"4C7B",
			x"0000" when x"4C7C",
			x"0000" when x"4C7D",
			x"0000" when x"4C7E",
			x"0000" when x"4C7F",
			x"0000" when x"4C80",
			x"0000" when x"4C81",
			x"0000" when x"4C82",
			x"0000" when x"4C83",
			x"0000" when x"4C84",
			x"0000" when x"4C85",
			x"0000" when x"4C86",
			x"0000" when x"4C87",
			x"0000" when x"4C88",
			x"0000" when x"4C89",
			x"0000" when x"4C8A",
			x"0000" when x"4C8B",
			x"0000" when x"4C8C",
			x"0000" when x"4C8D",
			x"0000" when x"4C8E",
			x"0000" when x"4C8F",
			x"0000" when x"4C90",
			x"0000" when x"4C91",
			x"0000" when x"4C92",
			x"0000" when x"4C93",
			x"0000" when x"4C94",
			x"0000" when x"4C95",
			x"0000" when x"4C96",
			x"0000" when x"4C97",
			x"0000" when x"4C98",
			x"0000" when x"4C99",
			x"0000" when x"4C9A",
			x"0000" when x"4C9B",
			x"0000" when x"4C9C",
			x"0000" when x"4C9D",
			x"0000" when x"4C9E",
			x"0000" when x"4C9F",
			x"0000" when x"4CA0",
			x"0000" when x"4CA1",
			x"0000" when x"4CA2",
			x"0000" when x"4CA3",
			x"0000" when x"4CA4",
			x"0000" when x"4CA5",
			x"0000" when x"4CA6",
			x"0000" when x"4CA7",
			x"0000" when x"4CA8",
			x"0000" when x"4CA9",
			x"0000" when x"4CAA",
			x"0000" when x"4CAB",
			x"0000" when x"4CAC",
			x"0000" when x"4CAD",
			x"0000" when x"4CAE",
			x"0000" when x"4CAF",
			x"0000" when x"4CB0",
			x"0000" when x"4CB1",
			x"0000" when x"4CB2",
			x"0000" when x"4CB3",
			x"0000" when x"4CB4",
			x"0000" when x"4CB5",
			x"0000" when x"4CB6",
			x"0000" when x"4CB7",
			x"0000" when x"4CB8",
			x"0000" when x"4CB9",
			x"0000" when x"4CBA",
			x"0000" when x"4CBB",
			x"0000" when x"4CBC",
			x"0000" when x"4CBD",
			x"0000" when x"4CBE",
			x"0000" when x"4CBF",
			x"0000" when x"4CC0",
			x"0000" when x"4CC1",
			x"0000" when x"4CC2",
			x"0000" when x"4CC3",
			x"0000" when x"4CC4",
			x"0000" when x"4CC5",
			x"0000" when x"4CC6",
			x"0000" when x"4CC7",
			x"0000" when x"4CC8",
			x"0000" when x"4CC9",
			x"0000" when x"4CCA",
			x"0000" when x"4CCB",
			x"0000" when x"4CCC",
			x"0000" when x"4CCD",
			x"0000" when x"4CCE",
			x"0000" when x"4CCF",
			x"0000" when x"4CD0",
			x"0000" when x"4CD1",
			x"0000" when x"4CD2",
			x"0000" when x"4CD3",
			x"0000" when x"4CD4",
			x"0000" when x"4CD5",
			x"0000" when x"4CD6",
			x"0000" when x"4CD7",
			x"0000" when x"4CD8",
			x"0000" when x"4CD9",
			x"0000" when x"4CDA",
			x"0000" when x"4CDB",
			x"0000" when x"4CDC",
			x"0000" when x"4CDD",
			x"0000" when x"4CDE",
			x"0000" when x"4CDF",
			x"0000" when x"4CE0",
			x"0000" when x"4CE1",
			x"0000" when x"4CE2",
			x"0000" when x"4CE3",
			x"0000" when x"4CE4",
			x"0000" when x"4CE5",
			x"0000" when x"4CE6",
			x"0000" when x"4CE7",
			x"0000" when x"4CE8",
			x"0000" when x"4CE9",
			x"0000" when x"4CEA",
			x"0000" when x"4CEB",
			x"0000" when x"4CEC",
			x"0000" when x"4CED",
			x"0000" when x"4CEE",
			x"0000" when x"4CEF",
			x"0000" when x"4CF0",
			x"0000" when x"4CF1",
			x"0000" when x"4CF2",
			x"0000" when x"4CF3",
			x"0000" when x"4CF4",
			x"0000" when x"4CF5",
			x"0000" when x"4CF6",
			x"0000" when x"4CF7",
			x"0000" when x"4CF8",
			x"0000" when x"4CF9",
			x"0000" when x"4CFA",
			x"0000" when x"4CFB",
			x"0000" when x"4CFC",
			x"0000" when x"4CFD",
			x"0000" when x"4CFE",
			x"0000" when x"4CFF",
			x"0000" when x"4D00",
			x"0000" when x"4D01",
			x"0000" when x"4D02",
			x"0000" when x"4D03",
			x"0000" when x"4D04",
			x"0000" when x"4D05",
			x"0000" when x"4D06",
			x"0000" when x"4D07",
			x"0000" when x"4D08",
			x"0000" when x"4D09",
			x"0000" when x"4D0A",
			x"0000" when x"4D0B",
			x"0000" when x"4D0C",
			x"0000" when x"4D0D",
			x"0000" when x"4D0E",
			x"0000" when x"4D0F",
			x"0000" when x"4D10",
			x"0000" when x"4D11",
			x"0000" when x"4D12",
			x"0000" when x"4D13",
			x"0000" when x"4D14",
			x"0000" when x"4D15",
			x"0000" when x"4D16",
			x"0000" when x"4D17",
			x"0000" when x"4D18",
			x"0000" when x"4D19",
			x"0000" when x"4D1A",
			x"0000" when x"4D1B",
			x"0000" when x"4D1C",
			x"0000" when x"4D1D",
			x"0000" when x"4D1E",
			x"0000" when x"4D1F",
			x"0000" when x"4D20",
			x"0000" when x"4D21",
			x"0000" when x"4D22",
			x"0000" when x"4D23",
			x"0000" when x"4D24",
			x"0000" when x"4D25",
			x"0000" when x"4D26",
			x"0000" when x"4D27",
			x"0000" when x"4D28",
			x"0000" when x"4D29",
			x"0000" when x"4D2A",
			x"0000" when x"4D2B",
			x"0000" when x"4D2C",
			x"0000" when x"4D2D",
			x"0000" when x"4D2E",
			x"0000" when x"4D2F",
			x"0000" when x"4D30",
			x"0000" when x"4D31",
			x"0000" when x"4D32",
			x"0000" when x"4D33",
			x"0000" when x"4D34",
			x"0000" when x"4D35",
			x"0000" when x"4D36",
			x"0000" when x"4D37",
			x"0000" when x"4D38",
			x"0000" when x"4D39",
			x"0000" when x"4D3A",
			x"0000" when x"4D3B",
			x"0000" when x"4D3C",
			x"0000" when x"4D3D",
			x"0000" when x"4D3E",
			x"0000" when x"4D3F",
			x"0000" when x"4D40",
			x"0000" when x"4D41",
			x"0000" when x"4D42",
			x"0000" when x"4D43",
			x"0000" when x"4D44",
			x"0000" when x"4D45",
			x"0000" when x"4D46",
			x"0000" when x"4D47",
			x"0000" when x"4D48",
			x"0000" when x"4D49",
			x"0000" when x"4D4A",
			x"0000" when x"4D4B",
			x"0000" when x"4D4C",
			x"0000" when x"4D4D",
			x"0000" when x"4D4E",
			x"0000" when x"4D4F",
			x"0000" when x"4D50",
			x"0000" when x"4D51",
			x"0000" when x"4D52",
			x"0000" when x"4D53",
			x"0000" when x"4D54",
			x"0000" when x"4D55",
			x"0000" when x"4D56",
			x"0000" when x"4D57",
			x"0000" when x"4D58",
			x"0000" when x"4D59",
			x"0000" when x"4D5A",
			x"0000" when x"4D5B",
			x"0000" when x"4D5C",
			x"0000" when x"4D5D",
			x"0000" when x"4D5E",
			x"0000" when x"4D5F",
			x"0000" when x"4D60",
			x"0000" when x"4D61",
			x"0000" when x"4D62",
			x"0000" when x"4D63",
			x"0000" when x"4D64",
			x"0000" when x"4D65",
			x"0000" when x"4D66",
			x"0000" when x"4D67",
			x"0000" when x"4D68",
			x"0000" when x"4D69",
			x"0000" when x"4D6A",
			x"0000" when x"4D6B",
			x"0000" when x"4D6C",
			x"0000" when x"4D6D",
			x"0000" when x"4D6E",
			x"0000" when x"4D6F",
			x"0000" when x"4D70",
			x"0000" when x"4D71",
			x"0000" when x"4D72",
			x"0000" when x"4D73",
			x"0000" when x"4D74",
			x"0000" when x"4D75",
			x"0000" when x"4D76",
			x"0000" when x"4D77",
			x"0000" when x"4D78",
			x"0000" when x"4D79",
			x"0000" when x"4D7A",
			x"0000" when x"4D7B",
			x"0000" when x"4D7C",
			x"0000" when x"4D7D",
			x"0000" when x"4D7E",
			x"0000" when x"4D7F",
			x"0000" when x"4D80",
			x"0000" when x"4D81",
			x"0000" when x"4D82",
			x"0000" when x"4D83",
			x"0000" when x"4D84",
			x"0000" when x"4D85",
			x"0000" when x"4D86",
			x"0000" when x"4D87",
			x"0000" when x"4D88",
			x"0000" when x"4D89",
			x"0000" when x"4D8A",
			x"0000" when x"4D8B",
			x"0000" when x"4D8C",
			x"0000" when x"4D8D",
			x"0000" when x"4D8E",
			x"0000" when x"4D8F",
			x"0000" when x"4D90",
			x"0000" when x"4D91",
			x"0000" when x"4D92",
			x"0000" when x"4D93",
			x"0000" when x"4D94",
			x"0000" when x"4D95",
			x"0000" when x"4D96",
			x"0000" when x"4D97",
			x"0000" when x"4D98",
			x"0000" when x"4D99",
			x"0000" when x"4D9A",
			x"0000" when x"4D9B",
			x"0000" when x"4D9C",
			x"0000" when x"4D9D",
			x"0000" when x"4D9E",
			x"0000" when x"4D9F",
			x"0000" when x"4DA0",
			x"0000" when x"4DA1",
			x"0000" when x"4DA2",
			x"0000" when x"4DA3",
			x"0000" when x"4DA4",
			x"0000" when x"4DA5",
			x"0000" when x"4DA6",
			x"0000" when x"4DA7",
			x"0000" when x"4DA8",
			x"0000" when x"4DA9",
			x"0000" when x"4DAA",
			x"0000" when x"4DAB",
			x"0000" when x"4DAC",
			x"0000" when x"4DAD",
			x"0000" when x"4DAE",
			x"0000" when x"4DAF",
			x"0000" when x"4DB0",
			x"0000" when x"4DB1",
			x"0000" when x"4DB2",
			x"0000" when x"4DB3",
			x"0000" when x"4DB4",
			x"0000" when x"4DB5",
			x"0000" when x"4DB6",
			x"0000" when x"4DB7",
			x"0000" when x"4DB8",
			x"0000" when x"4DB9",
			x"0000" when x"4DBA",
			x"0000" when x"4DBB",
			x"0000" when x"4DBC",
			x"0000" when x"4DBD",
			x"0000" when x"4DBE",
			x"0000" when x"4DBF",
			x"0000" when x"4DC0",
			x"0000" when x"4DC1",
			x"0000" when x"4DC2",
			x"0000" when x"4DC3",
			x"0000" when x"4DC4",
			x"0000" when x"4DC5",
			x"0000" when x"4DC6",
			x"0000" when x"4DC7",
			x"0000" when x"4DC8",
			x"0000" when x"4DC9",
			x"0000" when x"4DCA",
			x"0000" when x"4DCB",
			x"0000" when x"4DCC",
			x"0000" when x"4DCD",
			x"0000" when x"4DCE",
			x"0000" when x"4DCF",
			x"0000" when x"4DD0",
			x"0000" when x"4DD1",
			x"0000" when x"4DD2",
			x"0000" when x"4DD3",
			x"0000" when x"4DD4",
			x"0000" when x"4DD5",
			x"0000" when x"4DD6",
			x"0000" when x"4DD7",
			x"0000" when x"4DD8",
			x"0000" when x"4DD9",
			x"0000" when x"4DDA",
			x"0000" when x"4DDB",
			x"0000" when x"4DDC",
			x"0000" when x"4DDD",
			x"0000" when x"4DDE",
			x"0000" when x"4DDF",
			x"0000" when x"4DE0",
			x"0000" when x"4DE1",
			x"0000" when x"4DE2",
			x"0000" when x"4DE3",
			x"0000" when x"4DE4",
			x"0000" when x"4DE5",
			x"0000" when x"4DE6",
			x"0000" when x"4DE7",
			x"0000" when x"4DE8",
			x"0000" when x"4DE9",
			x"0000" when x"4DEA",
			x"0000" when x"4DEB",
			x"0000" when x"4DEC",
			x"0000" when x"4DED",
			x"0000" when x"4DEE",
			x"0000" when x"4DEF",
			x"0000" when x"4DF0",
			x"0000" when x"4DF1",
			x"0000" when x"4DF2",
			x"0000" when x"4DF3",
			x"0000" when x"4DF4",
			x"0000" when x"4DF5",
			x"0000" when x"4DF6",
			x"0000" when x"4DF7",
			x"0000" when x"4DF8",
			x"0000" when x"4DF9",
			x"0000" when x"4DFA",
			x"0000" when x"4DFB",
			x"0000" when x"4DFC",
			x"0000" when x"4DFD",
			x"0000" when x"4DFE",
			x"0000" when x"4DFF",
			x"0000" when x"4E00",
			x"0000" when x"4E01",
			x"0000" when x"4E02",
			x"0000" when x"4E03",
			x"0000" when x"4E04",
			x"0000" when x"4E05",
			x"0000" when x"4E06",
			x"0000" when x"4E07",
			x"0000" when x"4E08",
			x"0000" when x"4E09",
			x"0000" when x"4E0A",
			x"0000" when x"4E0B",
			x"0000" when x"4E0C",
			x"0000" when x"4E0D",
			x"0000" when x"4E0E",
			x"0000" when x"4E0F",
			x"0000" when x"4E10",
			x"0000" when x"4E11",
			x"0000" when x"4E12",
			x"0000" when x"4E13",
			x"0000" when x"4E14",
			x"0000" when x"4E15",
			x"0000" when x"4E16",
			x"0000" when x"4E17",
			x"0000" when x"4E18",
			x"0000" when x"4E19",
			x"0000" when x"4E1A",
			x"0000" when x"4E1B",
			x"0000" when x"4E1C",
			x"0000" when x"4E1D",
			x"0000" when x"4E1E",
			x"0000" when x"4E1F",
			x"0000" when x"4E20",
			x"0000" when x"4E21",
			x"0000" when x"4E22",
			x"0000" when x"4E23",
			x"0000" when x"4E24",
			x"0000" when x"4E25",
			x"0000" when x"4E26",
			x"0000" when x"4E27",
			x"0000" when x"4E28",
			x"0000" when x"4E29",
			x"0000" when x"4E2A",
			x"0000" when x"4E2B",
			x"0000" when x"4E2C",
			x"0000" when x"4E2D",
			x"0000" when x"4E2E",
			x"0000" when x"4E2F",
			x"0000" when x"4E30",
			x"0000" when x"4E31",
			x"0000" when x"4E32",
			x"0000" when x"4E33",
			x"0000" when x"4E34",
			x"0000" when x"4E35",
			x"0000" when x"4E36",
			x"0000" when x"4E37",
			x"0000" when x"4E38",
			x"0000" when x"4E39",
			x"0000" when x"4E3A",
			x"0000" when x"4E3B",
			x"0000" when x"4E3C",
			x"0000" when x"4E3D",
			x"0000" when x"4E3E",
			x"0000" when x"4E3F",
			x"0000" when x"4E40",
			x"0000" when x"4E41",
			x"0000" when x"4E42",
			x"0000" when x"4E43",
			x"0000" when x"4E44",
			x"0000" when x"4E45",
			x"0000" when x"4E46",
			x"0000" when x"4E47",
			x"0000" when x"4E48",
			x"0000" when x"4E49",
			x"0000" when x"4E4A",
			x"0000" when x"4E4B",
			x"0000" when x"4E4C",
			x"0000" when x"4E4D",
			x"0000" when x"4E4E",
			x"0000" when x"4E4F",
			x"0000" when x"4E50",
			x"0000" when x"4E51",
			x"0000" when x"4E52",
			x"0000" when x"4E53",
			x"0000" when x"4E54",
			x"0000" when x"4E55",
			x"0000" when x"4E56",
			x"0000" when x"4E57",
			x"0000" when x"4E58",
			x"0000" when x"4E59",
			x"0000" when x"4E5A",
			x"0000" when x"4E5B",
			x"0000" when x"4E5C",
			x"0000" when x"4E5D",
			x"0000" when x"4E5E",
			x"0000" when x"4E5F",
			x"0000" when x"4E60",
			x"0000" when x"4E61",
			x"0000" when x"4E62",
			x"0000" when x"4E63",
			x"0000" when x"4E64",
			x"0000" when x"4E65",
			x"0000" when x"4E66",
			x"0000" when x"4E67",
			x"0000" when x"4E68",
			x"0000" when x"4E69",
			x"0000" when x"4E6A",
			x"0000" when x"4E6B",
			x"0000" when x"4E6C",
			x"0000" when x"4E6D",
			x"0000" when x"4E6E",
			x"0000" when x"4E6F",
			x"0000" when x"4E70",
			x"0000" when x"4E71",
			x"0000" when x"4E72",
			x"0000" when x"4E73",
			x"0000" when x"4E74",
			x"0000" when x"4E75",
			x"0000" when x"4E76",
			x"0000" when x"4E77",
			x"0000" when x"4E78",
			x"0000" when x"4E79",
			x"0000" when x"4E7A",
			x"0000" when x"4E7B",
			x"0000" when x"4E7C",
			x"0000" when x"4E7D",
			x"0000" when x"4E7E",
			x"0000" when x"4E7F",
			x"0000" when x"4E80",
			x"0000" when x"4E81",
			x"0000" when x"4E82",
			x"0000" when x"4E83",
			x"0000" when x"4E84",
			x"0000" when x"4E85",
			x"0000" when x"4E86",
			x"0000" when x"4E87",
			x"0000" when x"4E88",
			x"0000" when x"4E89",
			x"0000" when x"4E8A",
			x"0000" when x"4E8B",
			x"0000" when x"4E8C",
			x"0000" when x"4E8D",
			x"0000" when x"4E8E",
			x"0000" when x"4E8F",
			x"0000" when x"4E90",
			x"0000" when x"4E91",
			x"0000" when x"4E92",
			x"0000" when x"4E93",
			x"0000" when x"4E94",
			x"0000" when x"4E95",
			x"0000" when x"4E96",
			x"0000" when x"4E97",
			x"0000" when x"4E98",
			x"0000" when x"4E99",
			x"0000" when x"4E9A",
			x"0000" when x"4E9B",
			x"0000" when x"4E9C",
			x"0000" when x"4E9D",
			x"0000" when x"4E9E",
			x"0000" when x"4E9F",
			x"0000" when x"4EA0",
			x"0000" when x"4EA1",
			x"0000" when x"4EA2",
			x"0000" when x"4EA3",
			x"0000" when x"4EA4",
			x"0000" when x"4EA5",
			x"0000" when x"4EA6",
			x"0000" when x"4EA7",
			x"0000" when x"4EA8",
			x"0000" when x"4EA9",
			x"0000" when x"4EAA",
			x"0000" when x"4EAB",
			x"0000" when x"4EAC",
			x"0000" when x"4EAD",
			x"0000" when x"4EAE",
			x"0000" when x"4EAF",
			x"0000" when x"4EB0",
			x"0000" when x"4EB1",
			x"0000" when x"4EB2",
			x"0000" when x"4EB3",
			x"0000" when x"4EB4",
			x"0000" when x"4EB5",
			x"0000" when x"4EB6",
			x"0000" when x"4EB7",
			x"0000" when x"4EB8",
			x"0000" when x"4EB9",
			x"0000" when x"4EBA",
			x"0000" when x"4EBB",
			x"0000" when x"4EBC",
			x"0000" when x"4EBD",
			x"0000" when x"4EBE",
			x"0000" when x"4EBF",
			x"0000" when x"4EC0",
			x"0000" when x"4EC1",
			x"0000" when x"4EC2",
			x"0000" when x"4EC3",
			x"0000" when x"4EC4",
			x"0000" when x"4EC5",
			x"0000" when x"4EC6",
			x"0000" when x"4EC7",
			x"0000" when x"4EC8",
			x"0000" when x"4EC9",
			x"0000" when x"4ECA",
			x"0000" when x"4ECB",
			x"0000" when x"4ECC",
			x"0000" when x"4ECD",
			x"0000" when x"4ECE",
			x"0000" when x"4ECF",
			x"0000" when x"4ED0",
			x"0000" when x"4ED1",
			x"0000" when x"4ED2",
			x"0000" when x"4ED3",
			x"0000" when x"4ED4",
			x"0000" when x"4ED5",
			x"0000" when x"4ED6",
			x"0000" when x"4ED7",
			x"0000" when x"4ED8",
			x"0000" when x"4ED9",
			x"0000" when x"4EDA",
			x"0000" when x"4EDB",
			x"0000" when x"4EDC",
			x"0000" when x"4EDD",
			x"0000" when x"4EDE",
			x"0000" when x"4EDF",
			x"0000" when x"4EE0",
			x"0000" when x"4EE1",
			x"0000" when x"4EE2",
			x"0000" when x"4EE3",
			x"0000" when x"4EE4",
			x"0000" when x"4EE5",
			x"0000" when x"4EE6",
			x"0000" when x"4EE7",
			x"0000" when x"4EE8",
			x"0000" when x"4EE9",
			x"0000" when x"4EEA",
			x"0000" when x"4EEB",
			x"0000" when x"4EEC",
			x"0000" when x"4EED",
			x"0000" when x"4EEE",
			x"0000" when x"4EEF",
			x"0000" when x"4EF0",
			x"0000" when x"4EF1",
			x"0000" when x"4EF2",
			x"0000" when x"4EF3",
			x"0000" when x"4EF4",
			x"0000" when x"4EF5",
			x"0000" when x"4EF6",
			x"0000" when x"4EF7",
			x"0000" when x"4EF8",
			x"0000" when x"4EF9",
			x"0000" when x"4EFA",
			x"0000" when x"4EFB",
			x"0000" when x"4EFC",
			x"0000" when x"4EFD",
			x"0000" when x"4EFE",
			x"0000" when x"4EFF",
			x"0000" when x"4F00",
			x"0000" when x"4F01",
			x"0000" when x"4F02",
			x"0000" when x"4F03",
			x"0000" when x"4F04",
			x"0000" when x"4F05",
			x"0000" when x"4F06",
			x"0000" when x"4F07",
			x"0000" when x"4F08",
			x"0000" when x"4F09",
			x"0000" when x"4F0A",
			x"0000" when x"4F0B",
			x"0000" when x"4F0C",
			x"0000" when x"4F0D",
			x"0000" when x"4F0E",
			x"0000" when x"4F0F",
			x"0000" when x"4F10",
			x"0000" when x"4F11",
			x"0000" when x"4F12",
			x"0000" when x"4F13",
			x"0000" when x"4F14",
			x"0000" when x"4F15",
			x"0000" when x"4F16",
			x"0000" when x"4F17",
			x"0000" when x"4F18",
			x"0000" when x"4F19",
			x"0000" when x"4F1A",
			x"0000" when x"4F1B",
			x"0000" when x"4F1C",
			x"0000" when x"4F1D",
			x"0000" when x"4F1E",
			x"0000" when x"4F1F",
			x"0000" when x"4F20",
			x"0000" when x"4F21",
			x"0000" when x"4F22",
			x"0000" when x"4F23",
			x"0000" when x"4F24",
			x"0000" when x"4F25",
			x"0000" when x"4F26",
			x"0000" when x"4F27",
			x"0000" when x"4F28",
			x"0000" when x"4F29",
			x"0000" when x"4F2A",
			x"0000" when x"4F2B",
			x"0000" when x"4F2C",
			x"0000" when x"4F2D",
			x"0000" when x"4F2E",
			x"0000" when x"4F2F",
			x"0000" when x"4F30",
			x"0000" when x"4F31",
			x"0000" when x"4F32",
			x"0000" when x"4F33",
			x"0000" when x"4F34",
			x"0000" when x"4F35",
			x"0000" when x"4F36",
			x"0000" when x"4F37",
			x"0000" when x"4F38",
			x"0000" when x"4F39",
			x"0000" when x"4F3A",
			x"0000" when x"4F3B",
			x"0000" when x"4F3C",
			x"0000" when x"4F3D",
			x"0000" when x"4F3E",
			x"0000" when x"4F3F",
			x"0000" when x"4F40",
			x"0000" when x"4F41",
			x"0000" when x"4F42",
			x"0000" when x"4F43",
			x"0000" when x"4F44",
			x"0000" when x"4F45",
			x"0000" when x"4F46",
			x"0000" when x"4F47",
			x"0000" when x"4F48",
			x"0000" when x"4F49",
			x"0000" when x"4F4A",
			x"0000" when x"4F4B",
			x"0000" when x"4F4C",
			x"0000" when x"4F4D",
			x"0000" when x"4F4E",
			x"0000" when x"4F4F",
			x"0000" when x"4F50",
			x"0000" when x"4F51",
			x"0000" when x"4F52",
			x"0000" when x"4F53",
			x"0000" when x"4F54",
			x"0000" when x"4F55",
			x"0000" when x"4F56",
			x"0000" when x"4F57",
			x"0000" when x"4F58",
			x"0000" when x"4F59",
			x"0000" when x"4F5A",
			x"0000" when x"4F5B",
			x"0000" when x"4F5C",
			x"0000" when x"4F5D",
			x"0000" when x"4F5E",
			x"0000" when x"4F5F",
			x"0000" when x"4F60",
			x"0000" when x"4F61",
			x"0000" when x"4F62",
			x"0000" when x"4F63",
			x"0000" when x"4F64",
			x"0000" when x"4F65",
			x"0000" when x"4F66",
			x"0000" when x"4F67",
			x"0000" when x"4F68",
			x"0000" when x"4F69",
			x"0000" when x"4F6A",
			x"0000" when x"4F6B",
			x"0000" when x"4F6C",
			x"0000" when x"4F6D",
			x"0000" when x"4F6E",
			x"0000" when x"4F6F",
			x"0000" when x"4F70",
			x"0000" when x"4F71",
			x"0000" when x"4F72",
			x"0000" when x"4F73",
			x"0000" when x"4F74",
			x"0000" when x"4F75",
			x"0000" when x"4F76",
			x"0000" when x"4F77",
			x"0000" when x"4F78",
			x"0000" when x"4F79",
			x"0000" when x"4F7A",
			x"0000" when x"4F7B",
			x"0000" when x"4F7C",
			x"0000" when x"4F7D",
			x"0000" when x"4F7E",
			x"0000" when x"4F7F",
			x"0000" when x"4F80",
			x"0000" when x"4F81",
			x"0000" when x"4F82",
			x"0000" when x"4F83",
			x"0000" when x"4F84",
			x"0000" when x"4F85",
			x"0000" when x"4F86",
			x"0000" when x"4F87",
			x"0000" when x"4F88",
			x"0000" when x"4F89",
			x"0000" when x"4F8A",
			x"0000" when x"4F8B",
			x"0000" when x"4F8C",
			x"0000" when x"4F8D",
			x"0000" when x"4F8E",
			x"0000" when x"4F8F",
			x"0000" when x"4F90",
			x"0000" when x"4F91",
			x"0000" when x"4F92",
			x"0000" when x"4F93",
			x"0000" when x"4F94",
			x"0000" when x"4F95",
			x"0000" when x"4F96",
			x"0000" when x"4F97",
			x"0000" when x"4F98",
			x"0000" when x"4F99",
			x"0000" when x"4F9A",
			x"0000" when x"4F9B",
			x"0000" when x"4F9C",
			x"0000" when x"4F9D",
			x"0000" when x"4F9E",
			x"0000" when x"4F9F",
			x"0000" when x"4FA0",
			x"0000" when x"4FA1",
			x"0000" when x"4FA2",
			x"0000" when x"4FA3",
			x"0000" when x"4FA4",
			x"0000" when x"4FA5",
			x"0000" when x"4FA6",
			x"0000" when x"4FA7",
			x"0000" when x"4FA8",
			x"0000" when x"4FA9",
			x"0000" when x"4FAA",
			x"0000" when x"4FAB",
			x"0000" when x"4FAC",
			x"0000" when x"4FAD",
			x"0000" when x"4FAE",
			x"0000" when x"4FAF",
			x"0000" when x"4FB0",
			x"0000" when x"4FB1",
			x"0000" when x"4FB2",
			x"0000" when x"4FB3",
			x"0000" when x"4FB4",
			x"0000" when x"4FB5",
			x"0000" when x"4FB6",
			x"0000" when x"4FB7",
			x"0000" when x"4FB8",
			x"0000" when x"4FB9",
			x"0000" when x"4FBA",
			x"0000" when x"4FBB",
			x"0000" when x"4FBC",
			x"0000" when x"4FBD",
			x"0000" when x"4FBE",
			x"0000" when x"4FBF",
			x"0000" when x"4FC0",
			x"0000" when x"4FC1",
			x"0000" when x"4FC2",
			x"0000" when x"4FC3",
			x"0000" when x"4FC4",
			x"0000" when x"4FC5",
			x"0000" when x"4FC6",
			x"0000" when x"4FC7",
			x"0000" when x"4FC8",
			x"0000" when x"4FC9",
			x"0000" when x"4FCA",
			x"0000" when x"4FCB",
			x"0000" when x"4FCC",
			x"0000" when x"4FCD",
			x"0000" when x"4FCE",
			x"0000" when x"4FCF",
			x"0000" when x"4FD0",
			x"0000" when x"4FD1",
			x"0000" when x"4FD2",
			x"0000" when x"4FD3",
			x"0000" when x"4FD4",
			x"0000" when x"4FD5",
			x"0000" when x"4FD6",
			x"0000" when x"4FD7",
			x"0000" when x"4FD8",
			x"0000" when x"4FD9",
			x"0000" when x"4FDA",
			x"0000" when x"4FDB",
			x"0000" when x"4FDC",
			x"0000" when x"4FDD",
			x"0000" when x"4FDE",
			x"0000" when x"4FDF",
			x"0000" when x"4FE0",
			x"0000" when x"4FE1",
			x"0000" when x"4FE2",
			x"0000" when x"4FE3",
			x"0000" when x"4FE4",
			x"0000" when x"4FE5",
			x"0000" when x"4FE6",
			x"0000" when x"4FE7",
			x"0000" when x"4FE8",
			x"0000" when x"4FE9",
			x"0000" when x"4FEA",
			x"0000" when x"4FEB",
			x"0000" when x"4FEC",
			x"0000" when x"4FED",
			x"0000" when x"4FEE",
			x"0000" when x"4FEF",
			x"0000" when x"4FF0",
			x"0000" when x"4FF1",
			x"0000" when x"4FF2",
			x"0000" when x"4FF3",
			x"0000" when x"4FF4",
			x"0000" when x"4FF5",
			x"0000" when x"4FF6",
			x"0000" when x"4FF7",
			x"0000" when x"4FF8",
			x"0000" when x"4FF9",
			x"0000" when x"4FFA",
			x"0000" when x"4FFB",
			x"0000" when x"4FFC",
			x"0000" when x"4FFD",
			x"0000" when x"4FFE",
			x"0000" when x"4FFF",
			x"0000" when x"5000",
			x"0000" when x"5001",
			x"0000" when x"5002",
			x"0000" when x"5003",
			x"0000" when x"5004",
			x"0000" when x"5005",
			x"0000" when x"5006",
			x"0000" when x"5007",
			x"0000" when x"5008",
			x"0000" when x"5009",
			x"0000" when x"500A",
			x"0000" when x"500B",
			x"0000" when x"500C",
			x"0000" when x"500D",
			x"0000" when x"500E",
			x"0000" when x"500F",
			x"0000" when x"5010",
			x"0000" when x"5011",
			x"0000" when x"5012",
			x"0000" when x"5013",
			x"0000" when x"5014",
			x"0000" when x"5015",
			x"0000" when x"5016",
			x"0000" when x"5017",
			x"0000" when x"5018",
			x"0000" when x"5019",
			x"0000" when x"501A",
			x"0000" when x"501B",
			x"0000" when x"501C",
			x"0000" when x"501D",
			x"0000" when x"501E",
			x"0000" when x"501F",
			x"0000" when x"5020",
			x"0000" when x"5021",
			x"0000" when x"5022",
			x"0000" when x"5023",
			x"0000" when x"5024",
			x"0000" when x"5025",
			x"0000" when x"5026",
			x"0000" when x"5027",
			x"0000" when x"5028",
			x"0000" when x"5029",
			x"0000" when x"502A",
			x"0000" when x"502B",
			x"0000" when x"502C",
			x"0000" when x"502D",
			x"0000" when x"502E",
			x"0000" when x"502F",
			x"0000" when x"5030",
			x"0000" when x"5031",
			x"0000" when x"5032",
			x"0000" when x"5033",
			x"0000" when x"5034",
			x"0000" when x"5035",
			x"0000" when x"5036",
			x"0000" when x"5037",
			x"0000" when x"5038",
			x"0000" when x"5039",
			x"0000" when x"503A",
			x"0000" when x"503B",
			x"0000" when x"503C",
			x"0000" when x"503D",
			x"0000" when x"503E",
			x"0000" when x"503F",
			x"0000" when x"5040",
			x"0000" when x"5041",
			x"0000" when x"5042",
			x"0000" when x"5043",
			x"0000" when x"5044",
			x"0000" when x"5045",
			x"0000" when x"5046",
			x"0000" when x"5047",
			x"0000" when x"5048",
			x"0000" when x"5049",
			x"0000" when x"504A",
			x"0000" when x"504B",
			x"0000" when x"504C",
			x"0000" when x"504D",
			x"0000" when x"504E",
			x"0000" when x"504F",
			x"0000" when x"5050",
			x"0000" when x"5051",
			x"0000" when x"5052",
			x"0000" when x"5053",
			x"0000" when x"5054",
			x"0000" when x"5055",
			x"0000" when x"5056",
			x"0000" when x"5057",
			x"0000" when x"5058",
			x"0000" when x"5059",
			x"0000" when x"505A",
			x"0000" when x"505B",
			x"0000" when x"505C",
			x"0000" when x"505D",
			x"0000" when x"505E",
			x"0000" when x"505F",
			x"0000" when x"5060",
			x"0000" when x"5061",
			x"0000" when x"5062",
			x"0000" when x"5063",
			x"0000" when x"5064",
			x"0000" when x"5065",
			x"0000" when x"5066",
			x"0000" when x"5067",
			x"0000" when x"5068",
			x"0000" when x"5069",
			x"0000" when x"506A",
			x"0000" when x"506B",
			x"0000" when x"506C",
			x"0000" when x"506D",
			x"0000" when x"506E",
			x"0000" when x"506F",
			x"0000" when x"5070",
			x"0000" when x"5071",
			x"0000" when x"5072",
			x"0000" when x"5073",
			x"0000" when x"5074",
			x"0000" when x"5075",
			x"0000" when x"5076",
			x"0000" when x"5077",
			x"0000" when x"5078",
			x"0000" when x"5079",
			x"0000" when x"507A",
			x"0000" when x"507B",
			x"0000" when x"507C",
			x"0000" when x"507D",
			x"0000" when x"507E",
			x"0000" when x"507F",
			x"0000" when x"5080",
			x"0000" when x"5081",
			x"0000" when x"5082",
			x"0000" when x"5083",
			x"0000" when x"5084",
			x"0000" when x"5085",
			x"0000" when x"5086",
			x"0000" when x"5087",
			x"0000" when x"5088",
			x"0000" when x"5089",
			x"0000" when x"508A",
			x"0000" when x"508B",
			x"0000" when x"508C",
			x"0000" when x"508D",
			x"0000" when x"508E",
			x"0000" when x"508F",
			x"0000" when x"5090",
			x"0000" when x"5091",
			x"0000" when x"5092",
			x"0000" when x"5093",
			x"0000" when x"5094",
			x"0000" when x"5095",
			x"0000" when x"5096",
			x"0000" when x"5097",
			x"0000" when x"5098",
			x"0000" when x"5099",
			x"0000" when x"509A",
			x"0000" when x"509B",
			x"0000" when x"509C",
			x"0000" when x"509D",
			x"0000" when x"509E",
			x"0000" when x"509F",
			x"0000" when x"50A0",
			x"0000" when x"50A1",
			x"0000" when x"50A2",
			x"0000" when x"50A3",
			x"0000" when x"50A4",
			x"0000" when x"50A5",
			x"0000" when x"50A6",
			x"0000" when x"50A7",
			x"0000" when x"50A8",
			x"0000" when x"50A9",
			x"0000" when x"50AA",
			x"0000" when x"50AB",
			x"0000" when x"50AC",
			x"0000" when x"50AD",
			x"0000" when x"50AE",
			x"0000" when x"50AF",
			x"0000" when x"50B0",
			x"0000" when x"50B1",
			x"0000" when x"50B2",
			x"0000" when x"50B3",
			x"0000" when x"50B4",
			x"0000" when x"50B5",
			x"0000" when x"50B6",
			x"0000" when x"50B7",
			x"0000" when x"50B8",
			x"0000" when x"50B9",
			x"0000" when x"50BA",
			x"0000" when x"50BB",
			x"0000" when x"50BC",
			x"0000" when x"50BD",
			x"0000" when x"50BE",
			x"0000" when x"50BF",
			x"0000" when x"50C0",
			x"0000" when x"50C1",
			x"0000" when x"50C2",
			x"0000" when x"50C3",
			x"0000" when x"50C4",
			x"0000" when x"50C5",
			x"0000" when x"50C6",
			x"0000" when x"50C7",
			x"0000" when x"50C8",
			x"0000" when x"50C9",
			x"0000" when x"50CA",
			x"0000" when x"50CB",
			x"0000" when x"50CC",
			x"0000" when x"50CD",
			x"0000" when x"50CE",
			x"0000" when x"50CF",
			x"0000" when x"50D0",
			x"0000" when x"50D1",
			x"0000" when x"50D2",
			x"0000" when x"50D3",
			x"0000" when x"50D4",
			x"0000" when x"50D5",
			x"0000" when x"50D6",
			x"0000" when x"50D7",
			x"0000" when x"50D8",
			x"0000" when x"50D9",
			x"0000" when x"50DA",
			x"0000" when x"50DB",
			x"0000" when x"50DC",
			x"0000" when x"50DD",
			x"0000" when x"50DE",
			x"0000" when x"50DF",
			x"0000" when x"50E0",
			x"0000" when x"50E1",
			x"0000" when x"50E2",
			x"0000" when x"50E3",
			x"0000" when x"50E4",
			x"0000" when x"50E5",
			x"0000" when x"50E6",
			x"0000" when x"50E7",
			x"0000" when x"50E8",
			x"0000" when x"50E9",
			x"0000" when x"50EA",
			x"0000" when x"50EB",
			x"0000" when x"50EC",
			x"0000" when x"50ED",
			x"0000" when x"50EE",
			x"0000" when x"50EF",
			x"0000" when x"50F0",
			x"0000" when x"50F1",
			x"0000" when x"50F2",
			x"0000" when x"50F3",
			x"0000" when x"50F4",
			x"0000" when x"50F5",
			x"0000" when x"50F6",
			x"0000" when x"50F7",
			x"0000" when x"50F8",
			x"0000" when x"50F9",
			x"0000" when x"50FA",
			x"0000" when x"50FB",
			x"0000" when x"50FC",
			x"0000" when x"50FD",
			x"0000" when x"50FE",
			x"0000" when x"50FF",
			x"0000" when x"5100",
			x"0000" when x"5101",
			x"0000" when x"5102",
			x"0000" when x"5103",
			x"0000" when x"5104",
			x"0000" when x"5105",
			x"0000" when x"5106",
			x"0000" when x"5107",
			x"0000" when x"5108",
			x"0000" when x"5109",
			x"0000" when x"510A",
			x"0000" when x"510B",
			x"0000" when x"510C",
			x"0000" when x"510D",
			x"0000" when x"510E",
			x"0000" when x"510F",
			x"0000" when x"5110",
			x"0000" when x"5111",
			x"0000" when x"5112",
			x"0000" when x"5113",
			x"0000" when x"5114",
			x"0000" when x"5115",
			x"0000" when x"5116",
			x"0000" when x"5117",
			x"0000" when x"5118",
			x"0000" when x"5119",
			x"0000" when x"511A",
			x"0000" when x"511B",
			x"0000" when x"511C",
			x"0000" when x"511D",
			x"0000" when x"511E",
			x"0000" when x"511F",
			x"0000" when x"5120",
			x"0000" when x"5121",
			x"0000" when x"5122",
			x"0000" when x"5123",
			x"0000" when x"5124",
			x"0000" when x"5125",
			x"0000" when x"5126",
			x"0000" when x"5127",
			x"0000" when x"5128",
			x"0000" when x"5129",
			x"0000" when x"512A",
			x"0000" when x"512B",
			x"0000" when x"512C",
			x"0000" when x"512D",
			x"0000" when x"512E",
			x"0000" when x"512F",
			x"0000" when x"5130",
			x"0000" when x"5131",
			x"0000" when x"5132",
			x"0000" when x"5133",
			x"0000" when x"5134",
			x"0000" when x"5135",
			x"0000" when x"5136",
			x"0000" when x"5137",
			x"0000" when x"5138",
			x"0000" when x"5139",
			x"0000" when x"513A",
			x"0000" when x"513B",
			x"0000" when x"513C",
			x"0000" when x"513D",
			x"0000" when x"513E",
			x"0000" when x"513F",
			x"0000" when x"5140",
			x"0000" when x"5141",
			x"0000" when x"5142",
			x"0000" when x"5143",
			x"0000" when x"5144",
			x"0000" when x"5145",
			x"0000" when x"5146",
			x"0000" when x"5147",
			x"0000" when x"5148",
			x"0000" when x"5149",
			x"0000" when x"514A",
			x"0000" when x"514B",
			x"0000" when x"514C",
			x"0000" when x"514D",
			x"0000" when x"514E",
			x"0000" when x"514F",
			x"0000" when x"5150",
			x"0000" when x"5151",
			x"0000" when x"5152",
			x"0000" when x"5153",
			x"0000" when x"5154",
			x"0000" when x"5155",
			x"0000" when x"5156",
			x"0000" when x"5157",
			x"0000" when x"5158",
			x"0000" when x"5159",
			x"0000" when x"515A",
			x"0000" when x"515B",
			x"0000" when x"515C",
			x"0000" when x"515D",
			x"0000" when x"515E",
			x"0000" when x"515F",
			x"0000" when x"5160",
			x"0000" when x"5161",
			x"0000" when x"5162",
			x"0000" when x"5163",
			x"0000" when x"5164",
			x"0000" when x"5165",
			x"0000" when x"5166",
			x"0000" when x"5167",
			x"0000" when x"5168",
			x"0000" when x"5169",
			x"0000" when x"516A",
			x"0000" when x"516B",
			x"0000" when x"516C",
			x"0000" when x"516D",
			x"0000" when x"516E",
			x"0000" when x"516F",
			x"0000" when x"5170",
			x"0000" when x"5171",
			x"0000" when x"5172",
			x"0000" when x"5173",
			x"0000" when x"5174",
			x"0000" when x"5175",
			x"0000" when x"5176",
			x"0000" when x"5177",
			x"0000" when x"5178",
			x"0000" when x"5179",
			x"0000" when x"517A",
			x"0000" when x"517B",
			x"0000" when x"517C",
			x"0000" when x"517D",
			x"0000" when x"517E",
			x"0000" when x"517F",
			x"0000" when x"5180",
			x"0000" when x"5181",
			x"0000" when x"5182",
			x"0000" when x"5183",
			x"0000" when x"5184",
			x"0000" when x"5185",
			x"0000" when x"5186",
			x"0000" when x"5187",
			x"0000" when x"5188",
			x"0000" when x"5189",
			x"0000" when x"518A",
			x"0000" when x"518B",
			x"0000" when x"518C",
			x"0000" when x"518D",
			x"0000" when x"518E",
			x"0000" when x"518F",
			x"0000" when x"5190",
			x"0000" when x"5191",
			x"0000" when x"5192",
			x"0000" when x"5193",
			x"0000" when x"5194",
			x"0000" when x"5195",
			x"0000" when x"5196",
			x"0000" when x"5197",
			x"0000" when x"5198",
			x"0000" when x"5199",
			x"0000" when x"519A",
			x"0000" when x"519B",
			x"0000" when x"519C",
			x"0000" when x"519D",
			x"0000" when x"519E",
			x"0000" when x"519F",
			x"0000" when x"51A0",
			x"0000" when x"51A1",
			x"0000" when x"51A2",
			x"0000" when x"51A3",
			x"0000" when x"51A4",
			x"0000" when x"51A5",
			x"0000" when x"51A6",
			x"0000" when x"51A7",
			x"0000" when x"51A8",
			x"0000" when x"51A9",
			x"0000" when x"51AA",
			x"0000" when x"51AB",
			x"0000" when x"51AC",
			x"0000" when x"51AD",
			x"0000" when x"51AE",
			x"0000" when x"51AF",
			x"0000" when x"51B0",
			x"0000" when x"51B1",
			x"0000" when x"51B2",
			x"0000" when x"51B3",
			x"0000" when x"51B4",
			x"0000" when x"51B5",
			x"0000" when x"51B6",
			x"0000" when x"51B7",
			x"0000" when x"51B8",
			x"0000" when x"51B9",
			x"0000" when x"51BA",
			x"0000" when x"51BB",
			x"0000" when x"51BC",
			x"0000" when x"51BD",
			x"0000" when x"51BE",
			x"0000" when x"51BF",
			x"0000" when x"51C0",
			x"0000" when x"51C1",
			x"0000" when x"51C2",
			x"0000" when x"51C3",
			x"0000" when x"51C4",
			x"0000" when x"51C5",
			x"0000" when x"51C6",
			x"0000" when x"51C7",
			x"0000" when x"51C8",
			x"0000" when x"51C9",
			x"0000" when x"51CA",
			x"0000" when x"51CB",
			x"0000" when x"51CC",
			x"0000" when x"51CD",
			x"0000" when x"51CE",
			x"0000" when x"51CF",
			x"0000" when x"51D0",
			x"0000" when x"51D1",
			x"0000" when x"51D2",
			x"0000" when x"51D3",
			x"0000" when x"51D4",
			x"0000" when x"51D5",
			x"0000" when x"51D6",
			x"0000" when x"51D7",
			x"0000" when x"51D8",
			x"0000" when x"51D9",
			x"0000" when x"51DA",
			x"0000" when x"51DB",
			x"0000" when x"51DC",
			x"0000" when x"51DD",
			x"0000" when x"51DE",
			x"0000" when x"51DF",
			x"0000" when x"51E0",
			x"0000" when x"51E1",
			x"0000" when x"51E2",
			x"0000" when x"51E3",
			x"0000" when x"51E4",
			x"0000" when x"51E5",
			x"0000" when x"51E6",
			x"0000" when x"51E7",
			x"0000" when x"51E8",
			x"0000" when x"51E9",
			x"0000" when x"51EA",
			x"0000" when x"51EB",
			x"0000" when x"51EC",
			x"0000" when x"51ED",
			x"0000" when x"51EE",
			x"0000" when x"51EF",
			x"0000" when x"51F0",
			x"0000" when x"51F1",
			x"0000" when x"51F2",
			x"0000" when x"51F3",
			x"0000" when x"51F4",
			x"0000" when x"51F5",
			x"0000" when x"51F6",
			x"0000" when x"51F7",
			x"0000" when x"51F8",
			x"0000" when x"51F9",
			x"0000" when x"51FA",
			x"0000" when x"51FB",
			x"0000" when x"51FC",
			x"0000" when x"51FD",
			x"0000" when x"51FE",
			x"0000" when x"51FF",
			x"0000" when x"5200",
			x"0000" when x"5201",
			x"0000" when x"5202",
			x"0000" when x"5203",
			x"0000" when x"5204",
			x"0000" when x"5205",
			x"0000" when x"5206",
			x"0000" when x"5207",
			x"0000" when x"5208",
			x"0000" when x"5209",
			x"0000" when x"520A",
			x"0000" when x"520B",
			x"0000" when x"520C",
			x"0000" when x"520D",
			x"0000" when x"520E",
			x"0000" when x"520F",
			x"0000" when x"5210",
			x"0000" when x"5211",
			x"0000" when x"5212",
			x"0000" when x"5213",
			x"0000" when x"5214",
			x"0000" when x"5215",
			x"0000" when x"5216",
			x"0000" when x"5217",
			x"0000" when x"5218",
			x"0000" when x"5219",
			x"0000" when x"521A",
			x"0000" when x"521B",
			x"0000" when x"521C",
			x"0000" when x"521D",
			x"0000" when x"521E",
			x"0000" when x"521F",
			x"0000" when x"5220",
			x"0000" when x"5221",
			x"0000" when x"5222",
			x"0000" when x"5223",
			x"0000" when x"5224",
			x"0000" when x"5225",
			x"0000" when x"5226",
			x"0000" when x"5227",
			x"0000" when x"5228",
			x"0000" when x"5229",
			x"0000" when x"522A",
			x"0000" when x"522B",
			x"0000" when x"522C",
			x"0000" when x"522D",
			x"0000" when x"522E",
			x"0000" when x"522F",
			x"0000" when x"5230",
			x"0000" when x"5231",
			x"0000" when x"5232",
			x"0000" when x"5233",
			x"0000" when x"5234",
			x"0000" when x"5235",
			x"0000" when x"5236",
			x"0000" when x"5237",
			x"0000" when x"5238",
			x"0000" when x"5239",
			x"0000" when x"523A",
			x"0000" when x"523B",
			x"0000" when x"523C",
			x"0000" when x"523D",
			x"0000" when x"523E",
			x"0000" when x"523F",
			x"0000" when x"5240",
			x"0000" when x"5241",
			x"0000" when x"5242",
			x"0000" when x"5243",
			x"0000" when x"5244",
			x"0000" when x"5245",
			x"0000" when x"5246",
			x"0000" when x"5247",
			x"0000" when x"5248",
			x"0000" when x"5249",
			x"0000" when x"524A",
			x"0000" when x"524B",
			x"0000" when x"524C",
			x"0000" when x"524D",
			x"0000" when x"524E",
			x"0000" when x"524F",
			x"0000" when x"5250",
			x"0000" when x"5251",
			x"0000" when x"5252",
			x"0000" when x"5253",
			x"0000" when x"5254",
			x"0000" when x"5255",
			x"0000" when x"5256",
			x"0000" when x"5257",
			x"0000" when x"5258",
			x"0000" when x"5259",
			x"0000" when x"525A",
			x"0000" when x"525B",
			x"0000" when x"525C",
			x"0000" when x"525D",
			x"0000" when x"525E",
			x"0000" when x"525F",
			x"0000" when x"5260",
			x"0000" when x"5261",
			x"0000" when x"5262",
			x"0000" when x"5263",
			x"0000" when x"5264",
			x"0000" when x"5265",
			x"0000" when x"5266",
			x"0000" when x"5267",
			x"0000" when x"5268",
			x"0000" when x"5269",
			x"0000" when x"526A",
			x"0000" when x"526B",
			x"0000" when x"526C",
			x"0000" when x"526D",
			x"0000" when x"526E",
			x"0000" when x"526F",
			x"0000" when x"5270",
			x"0000" when x"5271",
			x"0000" when x"5272",
			x"0000" when x"5273",
			x"0000" when x"5274",
			x"0000" when x"5275",
			x"0000" when x"5276",
			x"0000" when x"5277",
			x"0000" when x"5278",
			x"0000" when x"5279",
			x"0000" when x"527A",
			x"0000" when x"527B",
			x"0000" when x"527C",
			x"0000" when x"527D",
			x"0000" when x"527E",
			x"0000" when x"527F",
			x"0000" when x"5280",
			x"0000" when x"5281",
			x"0000" when x"5282",
			x"0000" when x"5283",
			x"0000" when x"5284",
			x"0000" when x"5285",
			x"0000" when x"5286",
			x"0000" when x"5287",
			x"0000" when x"5288",
			x"0000" when x"5289",
			x"0000" when x"528A",
			x"0000" when x"528B",
			x"0000" when x"528C",
			x"0000" when x"528D",
			x"0000" when x"528E",
			x"0000" when x"528F",
			x"0000" when x"5290",
			x"0000" when x"5291",
			x"0000" when x"5292",
			x"0000" when x"5293",
			x"0000" when x"5294",
			x"0000" when x"5295",
			x"0000" when x"5296",
			x"0000" when x"5297",
			x"0000" when x"5298",
			x"0000" when x"5299",
			x"0000" when x"529A",
			x"0000" when x"529B",
			x"0000" when x"529C",
			x"0000" when x"529D",
			x"0000" when x"529E",
			x"0000" when x"529F",
			x"0000" when x"52A0",
			x"0000" when x"52A1",
			x"0000" when x"52A2",
			x"0000" when x"52A3",
			x"0000" when x"52A4",
			x"0000" when x"52A5",
			x"0000" when x"52A6",
			x"0000" when x"52A7",
			x"0000" when x"52A8",
			x"0000" when x"52A9",
			x"0000" when x"52AA",
			x"0000" when x"52AB",
			x"0000" when x"52AC",
			x"0000" when x"52AD",
			x"0000" when x"52AE",
			x"0000" when x"52AF",
			x"0000" when x"52B0",
			x"0000" when x"52B1",
			x"0000" when x"52B2",
			x"0000" when x"52B3",
			x"0000" when x"52B4",
			x"0000" when x"52B5",
			x"0000" when x"52B6",
			x"0000" when x"52B7",
			x"0000" when x"52B8",
			x"0000" when x"52B9",
			x"0000" when x"52BA",
			x"0000" when x"52BB",
			x"0000" when x"52BC",
			x"0000" when x"52BD",
			x"0000" when x"52BE",
			x"0000" when x"52BF",
			x"0000" when x"52C0",
			x"0000" when x"52C1",
			x"0000" when x"52C2",
			x"0000" when x"52C3",
			x"0000" when x"52C4",
			x"0000" when x"52C5",
			x"0000" when x"52C6",
			x"0000" when x"52C7",
			x"0000" when x"52C8",
			x"0000" when x"52C9",
			x"0000" when x"52CA",
			x"0000" when x"52CB",
			x"0000" when x"52CC",
			x"0000" when x"52CD",
			x"0000" when x"52CE",
			x"0000" when x"52CF",
			x"0000" when x"52D0",
			x"0000" when x"52D1",
			x"0000" when x"52D2",
			x"0000" when x"52D3",
			x"0000" when x"52D4",
			x"0000" when x"52D5",
			x"0000" when x"52D6",
			x"0000" when x"52D7",
			x"0000" when x"52D8",
			x"0000" when x"52D9",
			x"0000" when x"52DA",
			x"0000" when x"52DB",
			x"0000" when x"52DC",
			x"0000" when x"52DD",
			x"0000" when x"52DE",
			x"0000" when x"52DF",
			x"0000" when x"52E0",
			x"0000" when x"52E1",
			x"0000" when x"52E2",
			x"0000" when x"52E3",
			x"0000" when x"52E4",
			x"0000" when x"52E5",
			x"0000" when x"52E6",
			x"0000" when x"52E7",
			x"0000" when x"52E8",
			x"0000" when x"52E9",
			x"0000" when x"52EA",
			x"0000" when x"52EB",
			x"0000" when x"52EC",
			x"0000" when x"52ED",
			x"0000" when x"52EE",
			x"0000" when x"52EF",
			x"0000" when x"52F0",
			x"0000" when x"52F1",
			x"0000" when x"52F2",
			x"0000" when x"52F3",
			x"0000" when x"52F4",
			x"0000" when x"52F5",
			x"0000" when x"52F6",
			x"0000" when x"52F7",
			x"0000" when x"52F8",
			x"0000" when x"52F9",
			x"0000" when x"52FA",
			x"0000" when x"52FB",
			x"0000" when x"52FC",
			x"0000" when x"52FD",
			x"0000" when x"52FE",
			x"0000" when x"52FF",
			x"0000" when x"5300",
			x"0000" when x"5301",
			x"0000" when x"5302",
			x"0000" when x"5303",
			x"0000" when x"5304",
			x"0000" when x"5305",
			x"0000" when x"5306",
			x"0000" when x"5307",
			x"0000" when x"5308",
			x"0000" when x"5309",
			x"0000" when x"530A",
			x"0000" when x"530B",
			x"0000" when x"530C",
			x"0000" when x"530D",
			x"0000" when x"530E",
			x"0000" when x"530F",
			x"0000" when x"5310",
			x"0000" when x"5311",
			x"0000" when x"5312",
			x"0000" when x"5313",
			x"0000" when x"5314",
			x"0000" when x"5315",
			x"0000" when x"5316",
			x"0000" when x"5317",
			x"0000" when x"5318",
			x"0000" when x"5319",
			x"0000" when x"531A",
			x"0000" when x"531B",
			x"0000" when x"531C",
			x"0000" when x"531D",
			x"0000" when x"531E",
			x"0000" when x"531F",
			x"0000" when x"5320",
			x"0000" when x"5321",
			x"0000" when x"5322",
			x"0000" when x"5323",
			x"0000" when x"5324",
			x"0000" when x"5325",
			x"0000" when x"5326",
			x"0000" when x"5327",
			x"0000" when x"5328",
			x"0000" when x"5329",
			x"0000" when x"532A",
			x"0000" when x"532B",
			x"0000" when x"532C",
			x"0000" when x"532D",
			x"0000" when x"532E",
			x"0000" when x"532F",
			x"0000" when x"5330",
			x"0000" when x"5331",
			x"0000" when x"5332",
			x"0000" when x"5333",
			x"0000" when x"5334",
			x"0000" when x"5335",
			x"0000" when x"5336",
			x"0000" when x"5337",
			x"0000" when x"5338",
			x"0000" when x"5339",
			x"0000" when x"533A",
			x"0000" when x"533B",
			x"0000" when x"533C",
			x"0000" when x"533D",
			x"0000" when x"533E",
			x"0000" when x"533F",
			x"0000" when x"5340",
			x"0000" when x"5341",
			x"0000" when x"5342",
			x"0000" when x"5343",
			x"0000" when x"5344",
			x"0000" when x"5345",
			x"0000" when x"5346",
			x"0000" when x"5347",
			x"0000" when x"5348",
			x"0000" when x"5349",
			x"0000" when x"534A",
			x"0000" when x"534B",
			x"0000" when x"534C",
			x"0000" when x"534D",
			x"0000" when x"534E",
			x"0000" when x"534F",
			x"0000" when x"5350",
			x"0000" when x"5351",
			x"0000" when x"5352",
			x"0000" when x"5353",
			x"0000" when x"5354",
			x"0000" when x"5355",
			x"0000" when x"5356",
			x"0000" when x"5357",
			x"0000" when x"5358",
			x"0000" when x"5359",
			x"0000" when x"535A",
			x"0000" when x"535B",
			x"0000" when x"535C",
			x"0000" when x"535D",
			x"0000" when x"535E",
			x"0000" when x"535F",
			x"0000" when x"5360",
			x"0000" when x"5361",
			x"0000" when x"5362",
			x"0000" when x"5363",
			x"0000" when x"5364",
			x"0000" when x"5365",
			x"0000" when x"5366",
			x"0000" when x"5367",
			x"0000" when x"5368",
			x"0000" when x"5369",
			x"0000" when x"536A",
			x"0000" when x"536B",
			x"0000" when x"536C",
			x"0000" when x"536D",
			x"0000" when x"536E",
			x"0000" when x"536F",
			x"0000" when x"5370",
			x"0000" when x"5371",
			x"0000" when x"5372",
			x"0000" when x"5373",
			x"0000" when x"5374",
			x"0000" when x"5375",
			x"0000" when x"5376",
			x"0000" when x"5377",
			x"0000" when x"5378",
			x"0000" when x"5379",
			x"0000" when x"537A",
			x"0000" when x"537B",
			x"0000" when x"537C",
			x"0000" when x"537D",
			x"0000" when x"537E",
			x"0000" when x"537F",
			x"0000" when x"5380",
			x"0000" when x"5381",
			x"0000" when x"5382",
			x"0000" when x"5383",
			x"0000" when x"5384",
			x"0000" when x"5385",
			x"0000" when x"5386",
			x"0000" when x"5387",
			x"0000" when x"5388",
			x"0000" when x"5389",
			x"0000" when x"538A",
			x"0000" when x"538B",
			x"0000" when x"538C",
			x"0000" when x"538D",
			x"0000" when x"538E",
			x"0000" when x"538F",
			x"0000" when x"5390",
			x"0000" when x"5391",
			x"0000" when x"5392",
			x"0000" when x"5393",
			x"0000" when x"5394",
			x"0000" when x"5395",
			x"0000" when x"5396",
			x"0000" when x"5397",
			x"0000" when x"5398",
			x"0000" when x"5399",
			x"0000" when x"539A",
			x"0000" when x"539B",
			x"0000" when x"539C",
			x"0000" when x"539D",
			x"0000" when x"539E",
			x"0000" when x"539F",
			x"0000" when x"53A0",
			x"0000" when x"53A1",
			x"0000" when x"53A2",
			x"0000" when x"53A3",
			x"0000" when x"53A4",
			x"0000" when x"53A5",
			x"0000" when x"53A6",
			x"0000" when x"53A7",
			x"0000" when x"53A8",
			x"0000" when x"53A9",
			x"0000" when x"53AA",
			x"0000" when x"53AB",
			x"0000" when x"53AC",
			x"0000" when x"53AD",
			x"0000" when x"53AE",
			x"0000" when x"53AF",
			x"0000" when x"53B0",
			x"0000" when x"53B1",
			x"0000" when x"53B2",
			x"0000" when x"53B3",
			x"0000" when x"53B4",
			x"0000" when x"53B5",
			x"0000" when x"53B6",
			x"0000" when x"53B7",
			x"0000" when x"53B8",
			x"0000" when x"53B9",
			x"0000" when x"53BA",
			x"0000" when x"53BB",
			x"0000" when x"53BC",
			x"0000" when x"53BD",
			x"0000" when x"53BE",
			x"0000" when x"53BF",
			x"0000" when x"53C0",
			x"0000" when x"53C1",
			x"0000" when x"53C2",
			x"0000" when x"53C3",
			x"0000" when x"53C4",
			x"0000" when x"53C5",
			x"0000" when x"53C6",
			x"0000" when x"53C7",
			x"0000" when x"53C8",
			x"0000" when x"53C9",
			x"0000" when x"53CA",
			x"0000" when x"53CB",
			x"0000" when x"53CC",
			x"0000" when x"53CD",
			x"0000" when x"53CE",
			x"0000" when x"53CF",
			x"0000" when x"53D0",
			x"0000" when x"53D1",
			x"0000" when x"53D2",
			x"0000" when x"53D3",
			x"0000" when x"53D4",
			x"0000" when x"53D5",
			x"0000" when x"53D6",
			x"0000" when x"53D7",
			x"0000" when x"53D8",
			x"0000" when x"53D9",
			x"0000" when x"53DA",
			x"0000" when x"53DB",
			x"0000" when x"53DC",
			x"0000" when x"53DD",
			x"0000" when x"53DE",
			x"0000" when x"53DF",
			x"0000" when x"53E0",
			x"0000" when x"53E1",
			x"0000" when x"53E2",
			x"0000" when x"53E3",
			x"0000" when x"53E4",
			x"0000" when x"53E5",
			x"0000" when x"53E6",
			x"0000" when x"53E7",
			x"0000" when x"53E8",
			x"0000" when x"53E9",
			x"0000" when x"53EA",
			x"0000" when x"53EB",
			x"0000" when x"53EC",
			x"0000" when x"53ED",
			x"0000" when x"53EE",
			x"0000" when x"53EF",
			x"0000" when x"53F0",
			x"0000" when x"53F1",
			x"0000" when x"53F2",
			x"0000" when x"53F3",
			x"0000" when x"53F4",
			x"0000" when x"53F5",
			x"0000" when x"53F6",
			x"0000" when x"53F7",
			x"0000" when x"53F8",
			x"0000" when x"53F9",
			x"0000" when x"53FA",
			x"0000" when x"53FB",
			x"0000" when x"53FC",
			x"0000" when x"53FD",
			x"0000" when x"53FE",
			x"0000" when x"53FF",
			x"0000" when x"5400",
			x"0000" when x"5401",
			x"0000" when x"5402",
			x"0000" when x"5403",
			x"0000" when x"5404",
			x"0000" when x"5405",
			x"0000" when x"5406",
			x"0000" when x"5407",
			x"0000" when x"5408",
			x"0000" when x"5409",
			x"0000" when x"540A",
			x"0000" when x"540B",
			x"0000" when x"540C",
			x"0000" when x"540D",
			x"0000" when x"540E",
			x"0000" when x"540F",
			x"0000" when x"5410",
			x"0000" when x"5411",
			x"0000" when x"5412",
			x"0000" when x"5413",
			x"0000" when x"5414",
			x"0000" when x"5415",
			x"0000" when x"5416",
			x"0000" when x"5417",
			x"0000" when x"5418",
			x"0000" when x"5419",
			x"0000" when x"541A",
			x"0000" when x"541B",
			x"0000" when x"541C",
			x"0000" when x"541D",
			x"0000" when x"541E",
			x"0000" when x"541F",
			x"0000" when x"5420",
			x"0000" when x"5421",
			x"0000" when x"5422",
			x"0000" when x"5423",
			x"0000" when x"5424",
			x"0000" when x"5425",
			x"0000" when x"5426",
			x"0000" when x"5427",
			x"0000" when x"5428",
			x"0000" when x"5429",
			x"0000" when x"542A",
			x"0000" when x"542B",
			x"0000" when x"542C",
			x"0000" when x"542D",
			x"0000" when x"542E",
			x"0000" when x"542F",
			x"0000" when x"5430",
			x"0000" when x"5431",
			x"0000" when x"5432",
			x"0000" when x"5433",
			x"0000" when x"5434",
			x"0000" when x"5435",
			x"0000" when x"5436",
			x"0000" when x"5437",
			x"0000" when x"5438",
			x"0000" when x"5439",
			x"0000" when x"543A",
			x"0000" when x"543B",
			x"0000" when x"543C",
			x"0000" when x"543D",
			x"0000" when x"543E",
			x"0000" when x"543F",
			x"0000" when x"5440",
			x"0000" when x"5441",
			x"0000" when x"5442",
			x"0000" when x"5443",
			x"0000" when x"5444",
			x"0000" when x"5445",
			x"0000" when x"5446",
			x"0000" when x"5447",
			x"0000" when x"5448",
			x"0000" when x"5449",
			x"0000" when x"544A",
			x"0000" when x"544B",
			x"0000" when x"544C",
			x"0000" when x"544D",
			x"0000" when x"544E",
			x"0000" when x"544F",
			x"0000" when x"5450",
			x"0000" when x"5451",
			x"0000" when x"5452",
			x"0000" when x"5453",
			x"0000" when x"5454",
			x"0000" when x"5455",
			x"0000" when x"5456",
			x"0000" when x"5457",
			x"0000" when x"5458",
			x"0000" when x"5459",
			x"0000" when x"545A",
			x"0000" when x"545B",
			x"0000" when x"545C",
			x"0000" when x"545D",
			x"0000" when x"545E",
			x"0000" when x"545F",
			x"0000" when x"5460",
			x"0000" when x"5461",
			x"0000" when x"5462",
			x"0000" when x"5463",
			x"0000" when x"5464",
			x"0000" when x"5465",
			x"0000" when x"5466",
			x"0000" when x"5467",
			x"0000" when x"5468",
			x"0000" when x"5469",
			x"0000" when x"546A",
			x"0000" when x"546B",
			x"0000" when x"546C",
			x"0000" when x"546D",
			x"0000" when x"546E",
			x"0000" when x"546F",
			x"0000" when x"5470",
			x"0000" when x"5471",
			x"0000" when x"5472",
			x"0000" when x"5473",
			x"0000" when x"5474",
			x"0000" when x"5475",
			x"0000" when x"5476",
			x"0000" when x"5477",
			x"0000" when x"5478",
			x"0000" when x"5479",
			x"0000" when x"547A",
			x"0000" when x"547B",
			x"0000" when x"547C",
			x"0000" when x"547D",
			x"0000" when x"547E",
			x"0000" when x"547F",
			x"0000" when x"5480",
			x"0000" when x"5481",
			x"0000" when x"5482",
			x"0000" when x"5483",
			x"0000" when x"5484",
			x"0000" when x"5485",
			x"0000" when x"5486",
			x"0000" when x"5487",
			x"0000" when x"5488",
			x"0000" when x"5489",
			x"0000" when x"548A",
			x"0000" when x"548B",
			x"0000" when x"548C",
			x"0000" when x"548D",
			x"0000" when x"548E",
			x"0000" when x"548F",
			x"0000" when x"5490",
			x"0000" when x"5491",
			x"0000" when x"5492",
			x"0000" when x"5493",
			x"0000" when x"5494",
			x"0000" when x"5495",
			x"0000" when x"5496",
			x"0000" when x"5497",
			x"0000" when x"5498",
			x"0000" when x"5499",
			x"0000" when x"549A",
			x"0000" when x"549B",
			x"0000" when x"549C",
			x"0000" when x"549D",
			x"0000" when x"549E",
			x"0000" when x"549F",
			x"0000" when x"54A0",
			x"0000" when x"54A1",
			x"0000" when x"54A2",
			x"0000" when x"54A3",
			x"0000" when x"54A4",
			x"0000" when x"54A5",
			x"0000" when x"54A6",
			x"0000" when x"54A7",
			x"0000" when x"54A8",
			x"0000" when x"54A9",
			x"0000" when x"54AA",
			x"0000" when x"54AB",
			x"0000" when x"54AC",
			x"0000" when x"54AD",
			x"0000" when x"54AE",
			x"0000" when x"54AF",
			x"0000" when x"54B0",
			x"0000" when x"54B1",
			x"0000" when x"54B2",
			x"0000" when x"54B3",
			x"0000" when x"54B4",
			x"0000" when x"54B5",
			x"0000" when x"54B6",
			x"0000" when x"54B7",
			x"0000" when x"54B8",
			x"0000" when x"54B9",
			x"0000" when x"54BA",
			x"0000" when x"54BB",
			x"0000" when x"54BC",
			x"0000" when x"54BD",
			x"0000" when x"54BE",
			x"0000" when x"54BF",
			x"0000" when x"54C0",
			x"0000" when x"54C1",
			x"0000" when x"54C2",
			x"0000" when x"54C3",
			x"0000" when x"54C4",
			x"0000" when x"54C5",
			x"0000" when x"54C6",
			x"0000" when x"54C7",
			x"0000" when x"54C8",
			x"0000" when x"54C9",
			x"0000" when x"54CA",
			x"0000" when x"54CB",
			x"0000" when x"54CC",
			x"0000" when x"54CD",
			x"0000" when x"54CE",
			x"0000" when x"54CF",
			x"0000" when x"54D0",
			x"0000" when x"54D1",
			x"0000" when x"54D2",
			x"0000" when x"54D3",
			x"0000" when x"54D4",
			x"0000" when x"54D5",
			x"0000" when x"54D6",
			x"0000" when x"54D7",
			x"0000" when x"54D8",
			x"0000" when x"54D9",
			x"0000" when x"54DA",
			x"0000" when x"54DB",
			x"0000" when x"54DC",
			x"0000" when x"54DD",
			x"0000" when x"54DE",
			x"0000" when x"54DF",
			x"0000" when x"54E0",
			x"0000" when x"54E1",
			x"0000" when x"54E2",
			x"0000" when x"54E3",
			x"0000" when x"54E4",
			x"0000" when x"54E5",
			x"0000" when x"54E6",
			x"0000" when x"54E7",
			x"0000" when x"54E8",
			x"0000" when x"54E9",
			x"0000" when x"54EA",
			x"0000" when x"54EB",
			x"0000" when x"54EC",
			x"0000" when x"54ED",
			x"0000" when x"54EE",
			x"0000" when x"54EF",
			x"0000" when x"54F0",
			x"0000" when x"54F1",
			x"0000" when x"54F2",
			x"0000" when x"54F3",
			x"0000" when x"54F4",
			x"0000" when x"54F5",
			x"0000" when x"54F6",
			x"0000" when x"54F7",
			x"0000" when x"54F8",
			x"0000" when x"54F9",
			x"0000" when x"54FA",
			x"0000" when x"54FB",
			x"0000" when x"54FC",
			x"0000" when x"54FD",
			x"0000" when x"54FE",
			x"0000" when x"54FF",
			x"0000" when x"5500",
			x"0000" when x"5501",
			x"0000" when x"5502",
			x"0000" when x"5503",
			x"0000" when x"5504",
			x"0000" when x"5505",
			x"0000" when x"5506",
			x"0000" when x"5507",
			x"0000" when x"5508",
			x"0000" when x"5509",
			x"0000" when x"550A",
			x"0000" when x"550B",
			x"0000" when x"550C",
			x"0000" when x"550D",
			x"0000" when x"550E",
			x"0000" when x"550F",
			x"0000" when x"5510",
			x"0000" when x"5511",
			x"0000" when x"5512",
			x"0000" when x"5513",
			x"0000" when x"5514",
			x"0000" when x"5515",
			x"0000" when x"5516",
			x"0000" when x"5517",
			x"0000" when x"5518",
			x"0000" when x"5519",
			x"0000" when x"551A",
			x"0000" when x"551B",
			x"0000" when x"551C",
			x"0000" when x"551D",
			x"0000" when x"551E",
			x"0000" when x"551F",
			x"0000" when x"5520",
			x"0000" when x"5521",
			x"0000" when x"5522",
			x"0000" when x"5523",
			x"0000" when x"5524",
			x"0000" when x"5525",
			x"0000" when x"5526",
			x"0000" when x"5527",
			x"0000" when x"5528",
			x"0000" when x"5529",
			x"0000" when x"552A",
			x"0000" when x"552B",
			x"0000" when x"552C",
			x"0000" when x"552D",
			x"0000" when x"552E",
			x"0000" when x"552F",
			x"0000" when x"5530",
			x"0000" when x"5531",
			x"0000" when x"5532",
			x"0000" when x"5533",
			x"0000" when x"5534",
			x"0000" when x"5535",
			x"0000" when x"5536",
			x"0000" when x"5537",
			x"0000" when x"5538",
			x"0000" when x"5539",
			x"0000" when x"553A",
			x"0000" when x"553B",
			x"0000" when x"553C",
			x"0000" when x"553D",
			x"0000" when x"553E",
			x"0000" when x"553F",
			x"0000" when x"5540",
			x"0000" when x"5541",
			x"0000" when x"5542",
			x"0000" when x"5543",
			x"0000" when x"5544",
			x"0000" when x"5545",
			x"0000" when x"5546",
			x"0000" when x"5547",
			x"0000" when x"5548",
			x"0000" when x"5549",
			x"0000" when x"554A",
			x"0000" when x"554B",
			x"0000" when x"554C",
			x"0000" when x"554D",
			x"0000" when x"554E",
			x"0000" when x"554F",
			x"0000" when x"5550",
			x"0000" when x"5551",
			x"0000" when x"5552",
			x"0000" when x"5553",
			x"0000" when x"5554",
			x"0000" when x"5555",
			x"0000" when x"5556",
			x"0000" when x"5557",
			x"0000" when x"5558",
			x"0000" when x"5559",
			x"0000" when x"555A",
			x"0000" when x"555B",
			x"0000" when x"555C",
			x"0000" when x"555D",
			x"0000" when x"555E",
			x"0000" when x"555F",
			x"0000" when x"5560",
			x"0000" when x"5561",
			x"0000" when x"5562",
			x"0000" when x"5563",
			x"0000" when x"5564",
			x"0000" when x"5565",
			x"0000" when x"5566",
			x"0000" when x"5567",
			x"0000" when x"5568",
			x"0000" when x"5569",
			x"0000" when x"556A",
			x"0000" when x"556B",
			x"0000" when x"556C",
			x"0000" when x"556D",
			x"0000" when x"556E",
			x"0000" when x"556F",
			x"0000" when x"5570",
			x"0000" when x"5571",
			x"0000" when x"5572",
			x"0000" when x"5573",
			x"0000" when x"5574",
			x"0000" when x"5575",
			x"0000" when x"5576",
			x"0000" when x"5577",
			x"0000" when x"5578",
			x"0000" when x"5579",
			x"0000" when x"557A",
			x"0000" when x"557B",
			x"0000" when x"557C",
			x"0000" when x"557D",
			x"0000" when x"557E",
			x"0000" when x"557F",
			x"0000" when x"5580",
			x"0000" when x"5581",
			x"0000" when x"5582",
			x"0000" when x"5583",
			x"0000" when x"5584",
			x"0000" when x"5585",
			x"0000" when x"5586",
			x"0000" when x"5587",
			x"0000" when x"5588",
			x"0000" when x"5589",
			x"0000" when x"558A",
			x"0000" when x"558B",
			x"0000" when x"558C",
			x"0000" when x"558D",
			x"0000" when x"558E",
			x"0000" when x"558F",
			x"0000" when x"5590",
			x"0000" when x"5591",
			x"0000" when x"5592",
			x"0000" when x"5593",
			x"0000" when x"5594",
			x"0000" when x"5595",
			x"0000" when x"5596",
			x"0000" when x"5597",
			x"0000" when x"5598",
			x"0000" when x"5599",
			x"0000" when x"559A",
			x"0000" when x"559B",
			x"0000" when x"559C",
			x"0000" when x"559D",
			x"0000" when x"559E",
			x"0000" when x"559F",
			x"0000" when x"55A0",
			x"0000" when x"55A1",
			x"0000" when x"55A2",
			x"0000" when x"55A3",
			x"0000" when x"55A4",
			x"0000" when x"55A5",
			x"0000" when x"55A6",
			x"0000" when x"55A7",
			x"0000" when x"55A8",
			x"0000" when x"55A9",
			x"0000" when x"55AA",
			x"0000" when x"55AB",
			x"0000" when x"55AC",
			x"0000" when x"55AD",
			x"0000" when x"55AE",
			x"0000" when x"55AF",
			x"0000" when x"55B0",
			x"0000" when x"55B1",
			x"0000" when x"55B2",
			x"0000" when x"55B3",
			x"0000" when x"55B4",
			x"0000" when x"55B5",
			x"0000" when x"55B6",
			x"0000" when x"55B7",
			x"0000" when x"55B8",
			x"0000" when x"55B9",
			x"0000" when x"55BA",
			x"0000" when x"55BB",
			x"0000" when x"55BC",
			x"0000" when x"55BD",
			x"0000" when x"55BE",
			x"0000" when x"55BF",
			x"0000" when x"55C0",
			x"0000" when x"55C1",
			x"0000" when x"55C2",
			x"0000" when x"55C3",
			x"0000" when x"55C4",
			x"0000" when x"55C5",
			x"0000" when x"55C6",
			x"0000" when x"55C7",
			x"0000" when x"55C8",
			x"0000" when x"55C9",
			x"0000" when x"55CA",
			x"0000" when x"55CB",
			x"0000" when x"55CC",
			x"0000" when x"55CD",
			x"0000" when x"55CE",
			x"0000" when x"55CF",
			x"0000" when x"55D0",
			x"0000" when x"55D1",
			x"0000" when x"55D2",
			x"0000" when x"55D3",
			x"0000" when x"55D4",
			x"0000" when x"55D5",
			x"0000" when x"55D6",
			x"0000" when x"55D7",
			x"0000" when x"55D8",
			x"0000" when x"55D9",
			x"0000" when x"55DA",
			x"0000" when x"55DB",
			x"0000" when x"55DC",
			x"0000" when x"55DD",
			x"0000" when x"55DE",
			x"0000" when x"55DF",
			x"0000" when x"55E0",
			x"0000" when x"55E1",
			x"0000" when x"55E2",
			x"0000" when x"55E3",
			x"0000" when x"55E4",
			x"0000" when x"55E5",
			x"0000" when x"55E6",
			x"0000" when x"55E7",
			x"0000" when x"55E8",
			x"0000" when x"55E9",
			x"0000" when x"55EA",
			x"0000" when x"55EB",
			x"0000" when x"55EC",
			x"0000" when x"55ED",
			x"0000" when x"55EE",
			x"0000" when x"55EF",
			x"0000" when x"55F0",
			x"0000" when x"55F1",
			x"0000" when x"55F2",
			x"0000" when x"55F3",
			x"0000" when x"55F4",
			x"0000" when x"55F5",
			x"0000" when x"55F6",
			x"0000" when x"55F7",
			x"0000" when x"55F8",
			x"0000" when x"55F9",
			x"0000" when x"55FA",
			x"0000" when x"55FB",
			x"0000" when x"55FC",
			x"0000" when x"55FD",
			x"0000" when x"55FE",
			x"0000" when x"55FF",
			x"0000" when x"5600",
			x"0000" when x"5601",
			x"0000" when x"5602",
			x"0000" when x"5603",
			x"0000" when x"5604",
			x"0000" when x"5605",
			x"0000" when x"5606",
			x"0000" when x"5607",
			x"0000" when x"5608",
			x"0000" when x"5609",
			x"0000" when x"560A",
			x"0000" when x"560B",
			x"0000" when x"560C",
			x"0000" when x"560D",
			x"0000" when x"560E",
			x"0000" when x"560F",
			x"0000" when x"5610",
			x"0000" when x"5611",
			x"0000" when x"5612",
			x"0000" when x"5613",
			x"0000" when x"5614",
			x"0000" when x"5615",
			x"0000" when x"5616",
			x"0000" when x"5617",
			x"0000" when x"5618",
			x"0000" when x"5619",
			x"0000" when x"561A",
			x"0000" when x"561B",
			x"0000" when x"561C",
			x"0000" when x"561D",
			x"0000" when x"561E",
			x"0000" when x"561F",
			x"0000" when x"5620",
			x"0000" when x"5621",
			x"0000" when x"5622",
			x"0000" when x"5623",
			x"0000" when x"5624",
			x"0000" when x"5625",
			x"0000" when x"5626",
			x"0000" when x"5627",
			x"0000" when x"5628",
			x"0000" when x"5629",
			x"0000" when x"562A",
			x"0000" when x"562B",
			x"0000" when x"562C",
			x"0000" when x"562D",
			x"0000" when x"562E",
			x"0000" when x"562F",
			x"0000" when x"5630",
			x"0000" when x"5631",
			x"0000" when x"5632",
			x"0000" when x"5633",
			x"0000" when x"5634",
			x"0000" when x"5635",
			x"0000" when x"5636",
			x"0000" when x"5637",
			x"0000" when x"5638",
			x"0000" when x"5639",
			x"0000" when x"563A",
			x"0000" when x"563B",
			x"0000" when x"563C",
			x"0000" when x"563D",
			x"0000" when x"563E",
			x"0000" when x"563F",
			x"0000" when x"5640",
			x"0000" when x"5641",
			x"0000" when x"5642",
			x"0000" when x"5643",
			x"0000" when x"5644",
			x"0000" when x"5645",
			x"0000" when x"5646",
			x"0000" when x"5647",
			x"0000" when x"5648",
			x"0000" when x"5649",
			x"0000" when x"564A",
			x"0000" when x"564B",
			x"0000" when x"564C",
			x"0000" when x"564D",
			x"0000" when x"564E",
			x"0000" when x"564F",
			x"0000" when x"5650",
			x"0000" when x"5651",
			x"0000" when x"5652",
			x"0000" when x"5653",
			x"0000" when x"5654",
			x"0000" when x"5655",
			x"0000" when x"5656",
			x"0000" when x"5657",
			x"0000" when x"5658",
			x"0000" when x"5659",
			x"0000" when x"565A",
			x"0000" when x"565B",
			x"0000" when x"565C",
			x"0000" when x"565D",
			x"0000" when x"565E",
			x"0000" when x"565F",
			x"0000" when x"5660",
			x"0000" when x"5661",
			x"0000" when x"5662",
			x"0000" when x"5663",
			x"0000" when x"5664",
			x"0000" when x"5665",
			x"0000" when x"5666",
			x"0000" when x"5667",
			x"0000" when x"5668",
			x"0000" when x"5669",
			x"0000" when x"566A",
			x"0000" when x"566B",
			x"0000" when x"566C",
			x"0000" when x"566D",
			x"0000" when x"566E",
			x"0000" when x"566F",
			x"0000" when x"5670",
			x"0000" when x"5671",
			x"0000" when x"5672",
			x"0000" when x"5673",
			x"0000" when x"5674",
			x"0000" when x"5675",
			x"0000" when x"5676",
			x"0000" when x"5677",
			x"0000" when x"5678",
			x"0000" when x"5679",
			x"0000" when x"567A",
			x"0000" when x"567B",
			x"0000" when x"567C",
			x"0000" when x"567D",
			x"0000" when x"567E",
			x"0000" when x"567F",
			x"0000" when x"5680",
			x"0000" when x"5681",
			x"0000" when x"5682",
			x"0000" when x"5683",
			x"0000" when x"5684",
			x"0000" when x"5685",
			x"0000" when x"5686",
			x"0000" when x"5687",
			x"0000" when x"5688",
			x"0000" when x"5689",
			x"0000" when x"568A",
			x"0000" when x"568B",
			x"0000" when x"568C",
			x"0000" when x"568D",
			x"0000" when x"568E",
			x"0000" when x"568F",
			x"0000" when x"5690",
			x"0000" when x"5691",
			x"0000" when x"5692",
			x"0000" when x"5693",
			x"0000" when x"5694",
			x"0000" when x"5695",
			x"0000" when x"5696",
			x"0000" when x"5697",
			x"0000" when x"5698",
			x"0000" when x"5699",
			x"0000" when x"569A",
			x"0000" when x"569B",
			x"0000" when x"569C",
			x"0000" when x"569D",
			x"0000" when x"569E",
			x"0000" when x"569F",
			x"0000" when x"56A0",
			x"0000" when x"56A1",
			x"0000" when x"56A2",
			x"0000" when x"56A3",
			x"0000" when x"56A4",
			x"0000" when x"56A5",
			x"0000" when x"56A6",
			x"0000" when x"56A7",
			x"0000" when x"56A8",
			x"0000" when x"56A9",
			x"0000" when x"56AA",
			x"0000" when x"56AB",
			x"0000" when x"56AC",
			x"0000" when x"56AD",
			x"0000" when x"56AE",
			x"0000" when x"56AF",
			x"0000" when x"56B0",
			x"0000" when x"56B1",
			x"0000" when x"56B2",
			x"0000" when x"56B3",
			x"0000" when x"56B4",
			x"0000" when x"56B5",
			x"0000" when x"56B6",
			x"0000" when x"56B7",
			x"0000" when x"56B8",
			x"0000" when x"56B9",
			x"0000" when x"56BA",
			x"0000" when x"56BB",
			x"0000" when x"56BC",
			x"0000" when x"56BD",
			x"0000" when x"56BE",
			x"0000" when x"56BF",
			x"0000" when x"56C0",
			x"0000" when x"56C1",
			x"0000" when x"56C2",
			x"0000" when x"56C3",
			x"0000" when x"56C4",
			x"0000" when x"56C5",
			x"0000" when x"56C6",
			x"0000" when x"56C7",
			x"0000" when x"56C8",
			x"0000" when x"56C9",
			x"0000" when x"56CA",
			x"0000" when x"56CB",
			x"0000" when x"56CC",
			x"0000" when x"56CD",
			x"0000" when x"56CE",
			x"0000" when x"56CF",
			x"0000" when x"56D0",
			x"0000" when x"56D1",
			x"0000" when x"56D2",
			x"0000" when x"56D3",
			x"0000" when x"56D4",
			x"0000" when x"56D5",
			x"0000" when x"56D6",
			x"0000" when x"56D7",
			x"0000" when x"56D8",
			x"0000" when x"56D9",
			x"0000" when x"56DA",
			x"0000" when x"56DB",
			x"0000" when x"56DC",
			x"0000" when x"56DD",
			x"0000" when x"56DE",
			x"0000" when x"56DF",
			x"0000" when x"56E0",
			x"0000" when x"56E1",
			x"0000" when x"56E2",
			x"0000" when x"56E3",
			x"0000" when x"56E4",
			x"0000" when x"56E5",
			x"0000" when x"56E6",
			x"0000" when x"56E7",
			x"0000" when x"56E8",
			x"0000" when x"56E9",
			x"0000" when x"56EA",
			x"0000" when x"56EB",
			x"0000" when x"56EC",
			x"0000" when x"56ED",
			x"0000" when x"56EE",
			x"0000" when x"56EF",
			x"0000" when x"56F0",
			x"0000" when x"56F1",
			x"0000" when x"56F2",
			x"0000" when x"56F3",
			x"0000" when x"56F4",
			x"0000" when x"56F5",
			x"0000" when x"56F6",
			x"0000" when x"56F7",
			x"0000" when x"56F8",
			x"0000" when x"56F9",
			x"0000" when x"56FA",
			x"0000" when x"56FB",
			x"0000" when x"56FC",
			x"0000" when x"56FD",
			x"0000" when x"56FE",
			x"0000" when x"56FF",
			x"0000" when x"5700",
			x"0000" when x"5701",
			x"0000" when x"5702",
			x"0000" when x"5703",
			x"0000" when x"5704",
			x"0000" when x"5705",
			x"0000" when x"5706",
			x"0000" when x"5707",
			x"0000" when x"5708",
			x"0000" when x"5709",
			x"0000" when x"570A",
			x"0000" when x"570B",
			x"0000" when x"570C",
			x"0000" when x"570D",
			x"0000" when x"570E",
			x"0000" when x"570F",
			x"0000" when x"5710",
			x"0000" when x"5711",
			x"0000" when x"5712",
			x"0000" when x"5713",
			x"0000" when x"5714",
			x"0000" when x"5715",
			x"0000" when x"5716",
			x"0000" when x"5717",
			x"0000" when x"5718",
			x"0000" when x"5719",
			x"0000" when x"571A",
			x"0000" when x"571B",
			x"0000" when x"571C",
			x"0000" when x"571D",
			x"0000" when x"571E",
			x"0000" when x"571F",
			x"0000" when x"5720",
			x"0000" when x"5721",
			x"0000" when x"5722",
			x"0000" when x"5723",
			x"0000" when x"5724",
			x"0000" when x"5725",
			x"0000" when x"5726",
			x"0000" when x"5727",
			x"0000" when x"5728",
			x"0000" when x"5729",
			x"0000" when x"572A",
			x"0000" when x"572B",
			x"0000" when x"572C",
			x"0000" when x"572D",
			x"0000" when x"572E",
			x"0000" when x"572F",
			x"0000" when x"5730",
			x"0000" when x"5731",
			x"0000" when x"5732",
			x"0000" when x"5733",
			x"0000" when x"5734",
			x"0000" when x"5735",
			x"0000" when x"5736",
			x"0000" when x"5737",
			x"0000" when x"5738",
			x"0000" when x"5739",
			x"0000" when x"573A",
			x"0000" when x"573B",
			x"0000" when x"573C",
			x"0000" when x"573D",
			x"0000" when x"573E",
			x"0000" when x"573F",
			x"0000" when x"5740",
			x"0000" when x"5741",
			x"0000" when x"5742",
			x"0000" when x"5743",
			x"0000" when x"5744",
			x"0000" when x"5745",
			x"0000" when x"5746",
			x"0000" when x"5747",
			x"0000" when x"5748",
			x"0000" when x"5749",
			x"0000" when x"574A",
			x"0000" when x"574B",
			x"0000" when x"574C",
			x"0000" when x"574D",
			x"0000" when x"574E",
			x"0000" when x"574F",
			x"0000" when x"5750",
			x"0000" when x"5751",
			x"0000" when x"5752",
			x"0000" when x"5753",
			x"0000" when x"5754",
			x"0000" when x"5755",
			x"0000" when x"5756",
			x"0000" when x"5757",
			x"0000" when x"5758",
			x"0000" when x"5759",
			x"0000" when x"575A",
			x"0000" when x"575B",
			x"0000" when x"575C",
			x"0000" when x"575D",
			x"0000" when x"575E",
			x"0000" when x"575F",
			x"0000" when x"5760",
			x"0000" when x"5761",
			x"0000" when x"5762",
			x"0000" when x"5763",
			x"0000" when x"5764",
			x"0000" when x"5765",
			x"0000" when x"5766",
			x"0000" when x"5767",
			x"0000" when x"5768",
			x"0000" when x"5769",
			x"0000" when x"576A",
			x"0000" when x"576B",
			x"0000" when x"576C",
			x"0000" when x"576D",
			x"0000" when x"576E",
			x"0000" when x"576F",
			x"0000" when x"5770",
			x"0000" when x"5771",
			x"0000" when x"5772",
			x"0000" when x"5773",
			x"0000" when x"5774",
			x"0000" when x"5775",
			x"0000" when x"5776",
			x"0000" when x"5777",
			x"0000" when x"5778",
			x"0000" when x"5779",
			x"0000" when x"577A",
			x"0000" when x"577B",
			x"0000" when x"577C",
			x"0000" when x"577D",
			x"0000" when x"577E",
			x"0000" when x"577F",
			x"0000" when x"5780",
			x"0000" when x"5781",
			x"0000" when x"5782",
			x"0000" when x"5783",
			x"0000" when x"5784",
			x"0000" when x"5785",
			x"0000" when x"5786",
			x"0000" when x"5787",
			x"0000" when x"5788",
			x"0000" when x"5789",
			x"0000" when x"578A",
			x"0000" when x"578B",
			x"0000" when x"578C",
			x"0000" when x"578D",
			x"0000" when x"578E",
			x"0000" when x"578F",
			x"0000" when x"5790",
			x"0000" when x"5791",
			x"0000" when x"5792",
			x"0000" when x"5793",
			x"0000" when x"5794",
			x"0000" when x"5795",
			x"0000" when x"5796",
			x"0000" when x"5797",
			x"0000" when x"5798",
			x"0000" when x"5799",
			x"0000" when x"579A",
			x"0000" when x"579B",
			x"0000" when x"579C",
			x"0000" when x"579D",
			x"0000" when x"579E",
			x"0000" when x"579F",
			x"0000" when x"57A0",
			x"0000" when x"57A1",
			x"0000" when x"57A2",
			x"0000" when x"57A3",
			x"0000" when x"57A4",
			x"0000" when x"57A5",
			x"0000" when x"57A6",
			x"0000" when x"57A7",
			x"0000" when x"57A8",
			x"0000" when x"57A9",
			x"0000" when x"57AA",
			x"0000" when x"57AB",
			x"0000" when x"57AC",
			x"0000" when x"57AD",
			x"0000" when x"57AE",
			x"0000" when x"57AF",
			x"0000" when x"57B0",
			x"0000" when x"57B1",
			x"0000" when x"57B2",
			x"0000" when x"57B3",
			x"0000" when x"57B4",
			x"0000" when x"57B5",
			x"0000" when x"57B6",
			x"0000" when x"57B7",
			x"0000" when x"57B8",
			x"0000" when x"57B9",
			x"0000" when x"57BA",
			x"0000" when x"57BB",
			x"0000" when x"57BC",
			x"0000" when x"57BD",
			x"0000" when x"57BE",
			x"0000" when x"57BF",
			x"0000" when x"57C0",
			x"0000" when x"57C1",
			x"0000" when x"57C2",
			x"0000" when x"57C3",
			x"0000" when x"57C4",
			x"0000" when x"57C5",
			x"0000" when x"57C6",
			x"0000" when x"57C7",
			x"0000" when x"57C8",
			x"0000" when x"57C9",
			x"0000" when x"57CA",
			x"0000" when x"57CB",
			x"0000" when x"57CC",
			x"0000" when x"57CD",
			x"0000" when x"57CE",
			x"0000" when x"57CF",
			x"0000" when x"57D0",
			x"0000" when x"57D1",
			x"0000" when x"57D2",
			x"0000" when x"57D3",
			x"0000" when x"57D4",
			x"0000" when x"57D5",
			x"0000" when x"57D6",
			x"0000" when x"57D7",
			x"0000" when x"57D8",
			x"0000" when x"57D9",
			x"0000" when x"57DA",
			x"0000" when x"57DB",
			x"0000" when x"57DC",
			x"0000" when x"57DD",
			x"0000" when x"57DE",
			x"0000" when x"57DF",
			x"0000" when x"57E0",
			x"0000" when x"57E1",
			x"0000" when x"57E2",
			x"0000" when x"57E3",
			x"0000" when x"57E4",
			x"0000" when x"57E5",
			x"0000" when x"57E6",
			x"0000" when x"57E7",
			x"0000" when x"57E8",
			x"0000" when x"57E9",
			x"0000" when x"57EA",
			x"0000" when x"57EB",
			x"0000" when x"57EC",
			x"0000" when x"57ED",
			x"0000" when x"57EE",
			x"0000" when x"57EF",
			x"0000" when x"57F0",
			x"0000" when x"57F1",
			x"0000" when x"57F2",
			x"0000" when x"57F3",
			x"0000" when x"57F4",
			x"0000" when x"57F5",
			x"0000" when x"57F6",
			x"0000" when x"57F7",
			x"0000" when x"57F8",
			x"0000" when x"57F9",
			x"0000" when x"57FA",
			x"0000" when x"57FB",
			x"0000" when x"57FC",
			x"0000" when x"57FD",
			x"0000" when x"57FE",
			x"0000" when x"57FF",
			x"0000" when x"5800",
			x"0000" when x"5801",
			x"0000" when x"5802",
			x"0000" when x"5803",
			x"0000" when x"5804",
			x"0000" when x"5805",
			x"0000" when x"5806",
			x"0000" when x"5807",
			x"0000" when x"5808",
			x"0000" when x"5809",
			x"0000" when x"580A",
			x"0000" when x"580B",
			x"0000" when x"580C",
			x"0000" when x"580D",
			x"0000" when x"580E",
			x"0000" when x"580F",
			x"0000" when x"5810",
			x"0000" when x"5811",
			x"0000" when x"5812",
			x"0000" when x"5813",
			x"0000" when x"5814",
			x"0000" when x"5815",
			x"0000" when x"5816",
			x"0000" when x"5817",
			x"0000" when x"5818",
			x"0000" when x"5819",
			x"0000" when x"581A",
			x"0000" when x"581B",
			x"0000" when x"581C",
			x"0000" when x"581D",
			x"0000" when x"581E",
			x"0000" when x"581F",
			x"0000" when x"5820",
			x"0000" when x"5821",
			x"0000" when x"5822",
			x"0000" when x"5823",
			x"0000" when x"5824",
			x"0000" when x"5825",
			x"0000" when x"5826",
			x"0000" when x"5827",
			x"0000" when x"5828",
			x"0000" when x"5829",
			x"0000" when x"582A",
			x"0000" when x"582B",
			x"0000" when x"582C",
			x"0000" when x"582D",
			x"0000" when x"582E",
			x"0000" when x"582F",
			x"0000" when x"5830",
			x"0000" when x"5831",
			x"0000" when x"5832",
			x"0000" when x"5833",
			x"0000" when x"5834",
			x"0000" when x"5835",
			x"0000" when x"5836",
			x"0000" when x"5837",
			x"0000" when x"5838",
			x"0000" when x"5839",
			x"0000" when x"583A",
			x"0000" when x"583B",
			x"0000" when x"583C",
			x"0000" when x"583D",
			x"0000" when x"583E",
			x"0000" when x"583F",
			x"0000" when x"5840",
			x"0000" when x"5841",
			x"0000" when x"5842",
			x"0000" when x"5843",
			x"0000" when x"5844",
			x"0000" when x"5845",
			x"0000" when x"5846",
			x"0000" when x"5847",
			x"0000" when x"5848",
			x"0000" when x"5849",
			x"0000" when x"584A",
			x"0000" when x"584B",
			x"0000" when x"584C",
			x"0000" when x"584D",
			x"0000" when x"584E",
			x"0000" when x"584F",
			x"0000" when x"5850",
			x"0000" when x"5851",
			x"0000" when x"5852",
			x"0000" when x"5853",
			x"0000" when x"5854",
			x"0000" when x"5855",
			x"0000" when x"5856",
			x"0000" when x"5857",
			x"0000" when x"5858",
			x"0000" when x"5859",
			x"0000" when x"585A",
			x"0000" when x"585B",
			x"0000" when x"585C",
			x"0000" when x"585D",
			x"0000" when x"585E",
			x"0000" when x"585F",
			x"0000" when x"5860",
			x"0000" when x"5861",
			x"0000" when x"5862",
			x"0000" when x"5863",
			x"0000" when x"5864",
			x"0000" when x"5865",
			x"0000" when x"5866",
			x"0000" when x"5867",
			x"0000" when x"5868",
			x"0000" when x"5869",
			x"0000" when x"586A",
			x"0000" when x"586B",
			x"0000" when x"586C",
			x"0000" when x"586D",
			x"0000" when x"586E",
			x"0000" when x"586F",
			x"0000" when x"5870",
			x"0000" when x"5871",
			x"0000" when x"5872",
			x"0000" when x"5873",
			x"0000" when x"5874",
			x"0000" when x"5875",
			x"0000" when x"5876",
			x"0000" when x"5877",
			x"0000" when x"5878",
			x"0000" when x"5879",
			x"0000" when x"587A",
			x"0000" when x"587B",
			x"0000" when x"587C",
			x"0000" when x"587D",
			x"0000" when x"587E",
			x"0000" when x"587F",
			x"0000" when x"5880",
			x"0000" when x"5881",
			x"0000" when x"5882",
			x"0000" when x"5883",
			x"0000" when x"5884",
			x"0000" when x"5885",
			x"0000" when x"5886",
			x"0000" when x"5887",
			x"0000" when x"5888",
			x"0000" when x"5889",
			x"0000" when x"588A",
			x"0000" when x"588B",
			x"0000" when x"588C",
			x"0000" when x"588D",
			x"0000" when x"588E",
			x"0000" when x"588F",
			x"0000" when x"5890",
			x"0000" when x"5891",
			x"0000" when x"5892",
			x"0000" when x"5893",
			x"0000" when x"5894",
			x"0000" when x"5895",
			x"0000" when x"5896",
			x"0000" when x"5897",
			x"0000" when x"5898",
			x"0000" when x"5899",
			x"0000" when x"589A",
			x"0000" when x"589B",
			x"0000" when x"589C",
			x"0000" when x"589D",
			x"0000" when x"589E",
			x"0000" when x"589F",
			x"0000" when x"58A0",
			x"0000" when x"58A1",
			x"0000" when x"58A2",
			x"0000" when x"58A3",
			x"0000" when x"58A4",
			x"0000" when x"58A5",
			x"0000" when x"58A6",
			x"0000" when x"58A7",
			x"0000" when x"58A8",
			x"0000" when x"58A9",
			x"0000" when x"58AA",
			x"0000" when x"58AB",
			x"0000" when x"58AC",
			x"0000" when x"58AD",
			x"0000" when x"58AE",
			x"0000" when x"58AF",
			x"0000" when x"58B0",
			x"0000" when x"58B1",
			x"0000" when x"58B2",
			x"0000" when x"58B3",
			x"0000" when x"58B4",
			x"0000" when x"58B5",
			x"0000" when x"58B6",
			x"0000" when x"58B7",
			x"0000" when x"58B8",
			x"0000" when x"58B9",
			x"0000" when x"58BA",
			x"0000" when x"58BB",
			x"0000" when x"58BC",
			x"0000" when x"58BD",
			x"0000" when x"58BE",
			x"0000" when x"58BF",
			x"0000" when x"58C0",
			x"0000" when x"58C1",
			x"0000" when x"58C2",
			x"0000" when x"58C3",
			x"0000" when x"58C4",
			x"0000" when x"58C5",
			x"0000" when x"58C6",
			x"0000" when x"58C7",
			x"0000" when x"58C8",
			x"0000" when x"58C9",
			x"0000" when x"58CA",
			x"0000" when x"58CB",
			x"0000" when x"58CC",
			x"0000" when x"58CD",
			x"0000" when x"58CE",
			x"0000" when x"58CF",
			x"0000" when x"58D0",
			x"0000" when x"58D1",
			x"0000" when x"58D2",
			x"0000" when x"58D3",
			x"0000" when x"58D4",
			x"0000" when x"58D5",
			x"0000" when x"58D6",
			x"0000" when x"58D7",
			x"0000" when x"58D8",
			x"0000" when x"58D9",
			x"0000" when x"58DA",
			x"0000" when x"58DB",
			x"0000" when x"58DC",
			x"0000" when x"58DD",
			x"0000" when x"58DE",
			x"0000" when x"58DF",
			x"0000" when x"58E0",
			x"0000" when x"58E1",
			x"0000" when x"58E2",
			x"0000" when x"58E3",
			x"0000" when x"58E4",
			x"0000" when x"58E5",
			x"0000" when x"58E6",
			x"0000" when x"58E7",
			x"0000" when x"58E8",
			x"0000" when x"58E9",
			x"0000" when x"58EA",
			x"0000" when x"58EB",
			x"0000" when x"58EC",
			x"0000" when x"58ED",
			x"0000" when x"58EE",
			x"0000" when x"58EF",
			x"0000" when x"58F0",
			x"0000" when x"58F1",
			x"0000" when x"58F2",
			x"0000" when x"58F3",
			x"0000" when x"58F4",
			x"0000" when x"58F5",
			x"0000" when x"58F6",
			x"0000" when x"58F7",
			x"0000" when x"58F8",
			x"0000" when x"58F9",
			x"0000" when x"58FA",
			x"0000" when x"58FB",
			x"0000" when x"58FC",
			x"0000" when x"58FD",
			x"0000" when x"58FE",
			x"0000" when x"58FF",
			x"0000" when x"5900",
			x"0000" when x"5901",
			x"0000" when x"5902",
			x"0000" when x"5903",
			x"0000" when x"5904",
			x"0000" when x"5905",
			x"0000" when x"5906",
			x"0000" when x"5907",
			x"0000" when x"5908",
			x"0000" when x"5909",
			x"0000" when x"590A",
			x"0000" when x"590B",
			x"0000" when x"590C",
			x"0000" when x"590D",
			x"0000" when x"590E",
			x"0000" when x"590F",
			x"0000" when x"5910",
			x"0000" when x"5911",
			x"0000" when x"5912",
			x"0000" when x"5913",
			x"0000" when x"5914",
			x"0000" when x"5915",
			x"0000" when x"5916",
			x"0000" when x"5917",
			x"0000" when x"5918",
			x"0000" when x"5919",
			x"0000" when x"591A",
			x"0000" when x"591B",
			x"0000" when x"591C",
			x"0000" when x"591D",
			x"0000" when x"591E",
			x"0000" when x"591F",
			x"0000" when x"5920",
			x"0000" when x"5921",
			x"0000" when x"5922",
			x"0000" when x"5923",
			x"0000" when x"5924",
			x"0000" when x"5925",
			x"0000" when x"5926",
			x"0000" when x"5927",
			x"0000" when x"5928",
			x"0000" when x"5929",
			x"0000" when x"592A",
			x"0000" when x"592B",
			x"0000" when x"592C",
			x"0000" when x"592D",
			x"0000" when x"592E",
			x"0000" when x"592F",
			x"0000" when x"5930",
			x"0000" when x"5931",
			x"0000" when x"5932",
			x"0000" when x"5933",
			x"0000" when x"5934",
			x"0000" when x"5935",
			x"0000" when x"5936",
			x"0000" when x"5937",
			x"0000" when x"5938",
			x"0000" when x"5939",
			x"0000" when x"593A",
			x"0000" when x"593B",
			x"0000" when x"593C",
			x"0000" when x"593D",
			x"0000" when x"593E",
			x"0000" when x"593F",
			x"0000" when x"5940",
			x"0000" when x"5941",
			x"0000" when x"5942",
			x"0000" when x"5943",
			x"0000" when x"5944",
			x"0000" when x"5945",
			x"0000" when x"5946",
			x"0000" when x"5947",
			x"0000" when x"5948",
			x"0000" when x"5949",
			x"0000" when x"594A",
			x"0000" when x"594B",
			x"0000" when x"594C",
			x"0000" when x"594D",
			x"0000" when x"594E",
			x"0000" when x"594F",
			x"0000" when x"5950",
			x"0000" when x"5951",
			x"0000" when x"5952",
			x"0000" when x"5953",
			x"0000" when x"5954",
			x"0000" when x"5955",
			x"0000" when x"5956",
			x"0000" when x"5957",
			x"0000" when x"5958",
			x"0000" when x"5959",
			x"0000" when x"595A",
			x"0000" when x"595B",
			x"0000" when x"595C",
			x"0000" when x"595D",
			x"0000" when x"595E",
			x"0000" when x"595F",
			x"0000" when x"5960",
			x"0000" when x"5961",
			x"0000" when x"5962",
			x"0000" when x"5963",
			x"0000" when x"5964",
			x"0000" when x"5965",
			x"0000" when x"5966",
			x"0000" when x"5967",
			x"0000" when x"5968",
			x"0000" when x"5969",
			x"0000" when x"596A",
			x"0000" when x"596B",
			x"0000" when x"596C",
			x"0000" when x"596D",
			x"0000" when x"596E",
			x"0000" when x"596F",
			x"0000" when x"5970",
			x"0000" when x"5971",
			x"0000" when x"5972",
			x"0000" when x"5973",
			x"0000" when x"5974",
			x"0000" when x"5975",
			x"0000" when x"5976",
			x"0000" when x"5977",
			x"0000" when x"5978",
			x"0000" when x"5979",
			x"0000" when x"597A",
			x"0000" when x"597B",
			x"0000" when x"597C",
			x"0000" when x"597D",
			x"0000" when x"597E",
			x"0000" when x"597F",
			x"0000" when x"5980",
			x"0000" when x"5981",
			x"0000" when x"5982",
			x"0000" when x"5983",
			x"0000" when x"5984",
			x"0000" when x"5985",
			x"0000" when x"5986",
			x"0000" when x"5987",
			x"0000" when x"5988",
			x"0000" when x"5989",
			x"0000" when x"598A",
			x"0000" when x"598B",
			x"0000" when x"598C",
			x"0000" when x"598D",
			x"0000" when x"598E",
			x"0000" when x"598F",
			x"0000" when x"5990",
			x"0000" when x"5991",
			x"0000" when x"5992",
			x"0000" when x"5993",
			x"0000" when x"5994",
			x"0000" when x"5995",
			x"0000" when x"5996",
			x"0000" when x"5997",
			x"0000" when x"5998",
			x"0000" when x"5999",
			x"0000" when x"599A",
			x"0000" when x"599B",
			x"0000" when x"599C",
			x"0000" when x"599D",
			x"0000" when x"599E",
			x"0000" when x"599F",
			x"0000" when x"59A0",
			x"0000" when x"59A1",
			x"0000" when x"59A2",
			x"0000" when x"59A3",
			x"0000" when x"59A4",
			x"0000" when x"59A5",
			x"0000" when x"59A6",
			x"0000" when x"59A7",
			x"0000" when x"59A8",
			x"0000" when x"59A9",
			x"0000" when x"59AA",
			x"0000" when x"59AB",
			x"0000" when x"59AC",
			x"0000" when x"59AD",
			x"0000" when x"59AE",
			x"0000" when x"59AF",
			x"0000" when x"59B0",
			x"0000" when x"59B1",
			x"0000" when x"59B2",
			x"0000" when x"59B3",
			x"0000" when x"59B4",
			x"0000" when x"59B5",
			x"0000" when x"59B6",
			x"0000" when x"59B7",
			x"0000" when x"59B8",
			x"0000" when x"59B9",
			x"0000" when x"59BA",
			x"0000" when x"59BB",
			x"0000" when x"59BC",
			x"0000" when x"59BD",
			x"0000" when x"59BE",
			x"0000" when x"59BF",
			x"0000" when x"59C0",
			x"0000" when x"59C1",
			x"0000" when x"59C2",
			x"0000" when x"59C3",
			x"0000" when x"59C4",
			x"0000" when x"59C5",
			x"0000" when x"59C6",
			x"0000" when x"59C7",
			x"0000" when x"59C8",
			x"0000" when x"59C9",
			x"0000" when x"59CA",
			x"0000" when x"59CB",
			x"0000" when x"59CC",
			x"0000" when x"59CD",
			x"0000" when x"59CE",
			x"0000" when x"59CF",
			x"0000" when x"59D0",
			x"0000" when x"59D1",
			x"0000" when x"59D2",
			x"0000" when x"59D3",
			x"0000" when x"59D4",
			x"0000" when x"59D5",
			x"0000" when x"59D6",
			x"0000" when x"59D7",
			x"0000" when x"59D8",
			x"0000" when x"59D9",
			x"0000" when x"59DA",
			x"0000" when x"59DB",
			x"0000" when x"59DC",
			x"0000" when x"59DD",
			x"0000" when x"59DE",
			x"0000" when x"59DF",
			x"0000" when x"59E0",
			x"0000" when x"59E1",
			x"0000" when x"59E2",
			x"0000" when x"59E3",
			x"0000" when x"59E4",
			x"0000" when x"59E5",
			x"0000" when x"59E6",
			x"0000" when x"59E7",
			x"0000" when x"59E8",
			x"0000" when x"59E9",
			x"0000" when x"59EA",
			x"0000" when x"59EB",
			x"0000" when x"59EC",
			x"0000" when x"59ED",
			x"0000" when x"59EE",
			x"0000" when x"59EF",
			x"0000" when x"59F0",
			x"0000" when x"59F1",
			x"0000" when x"59F2",
			x"0000" when x"59F3",
			x"0000" when x"59F4",
			x"0000" when x"59F5",
			x"0000" when x"59F6",
			x"0000" when x"59F7",
			x"0000" when x"59F8",
			x"0000" when x"59F9",
			x"0000" when x"59FA",
			x"0000" when x"59FB",
			x"0000" when x"59FC",
			x"0000" when x"59FD",
			x"0000" when x"59FE",
			x"0000" when x"59FF",
			x"0000" when x"5A00",
			x"0000" when x"5A01",
			x"0000" when x"5A02",
			x"0000" when x"5A03",
			x"0000" when x"5A04",
			x"0000" when x"5A05",
			x"0000" when x"5A06",
			x"0000" when x"5A07",
			x"0000" when x"5A08",
			x"0000" when x"5A09",
			x"0000" when x"5A0A",
			x"0000" when x"5A0B",
			x"0000" when x"5A0C",
			x"0000" when x"5A0D",
			x"0000" when x"5A0E",
			x"0000" when x"5A0F",
			x"0000" when x"5A10",
			x"0000" when x"5A11",
			x"0000" when x"5A12",
			x"0000" when x"5A13",
			x"0000" when x"5A14",
			x"0000" when x"5A15",
			x"0000" when x"5A16",
			x"0000" when x"5A17",
			x"0000" when x"5A18",
			x"0000" when x"5A19",
			x"0000" when x"5A1A",
			x"0000" when x"5A1B",
			x"0000" when x"5A1C",
			x"0000" when x"5A1D",
			x"0000" when x"5A1E",
			x"0000" when x"5A1F",
			x"0000" when x"5A20",
			x"0000" when x"5A21",
			x"0000" when x"5A22",
			x"0000" when x"5A23",
			x"0000" when x"5A24",
			x"0000" when x"5A25",
			x"0000" when x"5A26",
			x"0000" when x"5A27",
			x"0000" when x"5A28",
			x"0000" when x"5A29",
			x"0000" when x"5A2A",
			x"0000" when x"5A2B",
			x"0000" when x"5A2C",
			x"0000" when x"5A2D",
			x"0000" when x"5A2E",
			x"0000" when x"5A2F",
			x"0000" when x"5A30",
			x"0000" when x"5A31",
			x"0000" when x"5A32",
			x"0000" when x"5A33",
			x"0000" when x"5A34",
			x"0000" when x"5A35",
			x"0000" when x"5A36",
			x"0000" when x"5A37",
			x"0000" when x"5A38",
			x"0000" when x"5A39",
			x"0000" when x"5A3A",
			x"0000" when x"5A3B",
			x"0000" when x"5A3C",
			x"0000" when x"5A3D",
			x"0000" when x"5A3E",
			x"0000" when x"5A3F",
			x"0000" when x"5A40",
			x"0000" when x"5A41",
			x"0000" when x"5A42",
			x"0000" when x"5A43",
			x"0000" when x"5A44",
			x"0000" when x"5A45",
			x"0000" when x"5A46",
			x"0000" when x"5A47",
			x"0000" when x"5A48",
			x"0000" when x"5A49",
			x"0000" when x"5A4A",
			x"0000" when x"5A4B",
			x"0000" when x"5A4C",
			x"0000" when x"5A4D",
			x"0000" when x"5A4E",
			x"0000" when x"5A4F",
			x"0000" when x"5A50",
			x"0000" when x"5A51",
			x"0000" when x"5A52",
			x"0000" when x"5A53",
			x"0000" when x"5A54",
			x"0000" when x"5A55",
			x"0000" when x"5A56",
			x"0000" when x"5A57",
			x"0000" when x"5A58",
			x"0000" when x"5A59",
			x"0000" when x"5A5A",
			x"0000" when x"5A5B",
			x"0000" when x"5A5C",
			x"0000" when x"5A5D",
			x"0000" when x"5A5E",
			x"0000" when x"5A5F",
			x"0000" when x"5A60",
			x"0000" when x"5A61",
			x"0000" when x"5A62",
			x"0000" when x"5A63",
			x"0000" when x"5A64",
			x"0000" when x"5A65",
			x"0000" when x"5A66",
			x"0000" when x"5A67",
			x"0000" when x"5A68",
			x"0000" when x"5A69",
			x"0000" when x"5A6A",
			x"0000" when x"5A6B",
			x"0000" when x"5A6C",
			x"0000" when x"5A6D",
			x"0000" when x"5A6E",
			x"0000" when x"5A6F",
			x"0000" when x"5A70",
			x"0000" when x"5A71",
			x"0000" when x"5A72",
			x"0000" when x"5A73",
			x"0000" when x"5A74",
			x"0000" when x"5A75",
			x"0000" when x"5A76",
			x"0000" when x"5A77",
			x"0000" when x"5A78",
			x"0000" when x"5A79",
			x"0000" when x"5A7A",
			x"0000" when x"5A7B",
			x"0000" when x"5A7C",
			x"0000" when x"5A7D",
			x"0000" when x"5A7E",
			x"0000" when x"5A7F",
			x"0000" when x"5A80",
			x"0000" when x"5A81",
			x"0000" when x"5A82",
			x"0000" when x"5A83",
			x"0000" when x"5A84",
			x"0000" when x"5A85",
			x"0000" when x"5A86",
			x"0000" when x"5A87",
			x"0000" when x"5A88",
			x"0000" when x"5A89",
			x"0000" when x"5A8A",
			x"0000" when x"5A8B",
			x"0000" when x"5A8C",
			x"0000" when x"5A8D",
			x"0000" when x"5A8E",
			x"0000" when x"5A8F",
			x"0000" when x"5A90",
			x"0000" when x"5A91",
			x"0000" when x"5A92",
			x"0000" when x"5A93",
			x"0000" when x"5A94",
			x"0000" when x"5A95",
			x"0000" when x"5A96",
			x"0000" when x"5A97",
			x"0000" when x"5A98",
			x"0000" when x"5A99",
			x"0000" when x"5A9A",
			x"0000" when x"5A9B",
			x"0000" when x"5A9C",
			x"0000" when x"5A9D",
			x"0000" when x"5A9E",
			x"0000" when x"5A9F",
			x"0000" when x"5AA0",
			x"0000" when x"5AA1",
			x"0000" when x"5AA2",
			x"0000" when x"5AA3",
			x"0000" when x"5AA4",
			x"0000" when x"5AA5",
			x"0000" when x"5AA6",
			x"0000" when x"5AA7",
			x"0000" when x"5AA8",
			x"0000" when x"5AA9",
			x"0000" when x"5AAA",
			x"0000" when x"5AAB",
			x"0000" when x"5AAC",
			x"0000" when x"5AAD",
			x"0000" when x"5AAE",
			x"0000" when x"5AAF",
			x"0000" when x"5AB0",
			x"0000" when x"5AB1",
			x"0000" when x"5AB2",
			x"0000" when x"5AB3",
			x"0000" when x"5AB4",
			x"0000" when x"5AB5",
			x"0000" when x"5AB6",
			x"0000" when x"5AB7",
			x"0000" when x"5AB8",
			x"0000" when x"5AB9",
			x"0000" when x"5ABA",
			x"0000" when x"5ABB",
			x"0000" when x"5ABC",
			x"0000" when x"5ABD",
			x"0000" when x"5ABE",
			x"0000" when x"5ABF",
			x"0000" when x"5AC0",
			x"0000" when x"5AC1",
			x"0000" when x"5AC2",
			x"0000" when x"5AC3",
			x"0000" when x"5AC4",
			x"0000" when x"5AC5",
			x"0000" when x"5AC6",
			x"0000" when x"5AC7",
			x"0000" when x"5AC8",
			x"0000" when x"5AC9",
			x"0000" when x"5ACA",
			x"0000" when x"5ACB",
			x"0000" when x"5ACC",
			x"0000" when x"5ACD",
			x"0000" when x"5ACE",
			x"0000" when x"5ACF",
			x"0000" when x"5AD0",
			x"0000" when x"5AD1",
			x"0000" when x"5AD2",
			x"0000" when x"5AD3",
			x"0000" when x"5AD4",
			x"0000" when x"5AD5",
			x"0000" when x"5AD6",
			x"0000" when x"5AD7",
			x"0000" when x"5AD8",
			x"0000" when x"5AD9",
			x"0000" when x"5ADA",
			x"0000" when x"5ADB",
			x"0000" when x"5ADC",
			x"0000" when x"5ADD",
			x"0000" when x"5ADE",
			x"0000" when x"5ADF",
			x"0000" when x"5AE0",
			x"0000" when x"5AE1",
			x"0000" when x"5AE2",
			x"0000" when x"5AE3",
			x"0000" when x"5AE4",
			x"0000" when x"5AE5",
			x"0000" when x"5AE6",
			x"0000" when x"5AE7",
			x"0000" when x"5AE8",
			x"0000" when x"5AE9",
			x"0000" when x"5AEA",
			x"0000" when x"5AEB",
			x"0000" when x"5AEC",
			x"0000" when x"5AED",
			x"0000" when x"5AEE",
			x"0000" when x"5AEF",
			x"0000" when x"5AF0",
			x"0000" when x"5AF1",
			x"0000" when x"5AF2",
			x"0000" when x"5AF3",
			x"0000" when x"5AF4",
			x"0000" when x"5AF5",
			x"0000" when x"5AF6",
			x"0000" when x"5AF7",
			x"0000" when x"5AF8",
			x"0000" when x"5AF9",
			x"0000" when x"5AFA",
			x"0000" when x"5AFB",
			x"0000" when x"5AFC",
			x"0000" when x"5AFD",
			x"0000" when x"5AFE",
			x"0000" when x"5AFF",
			x"0000" when x"5B00",
			x"0000" when x"5B01",
			x"0000" when x"5B02",
			x"0000" when x"5B03",
			x"0000" when x"5B04",
			x"0000" when x"5B05",
			x"0000" when x"5B06",
			x"0000" when x"5B07",
			x"0000" when x"5B08",
			x"0000" when x"5B09",
			x"0000" when x"5B0A",
			x"0000" when x"5B0B",
			x"0000" when x"5B0C",
			x"0000" when x"5B0D",
			x"0000" when x"5B0E",
			x"0000" when x"5B0F",
			x"0000" when x"5B10",
			x"0000" when x"5B11",
			x"0000" when x"5B12",
			x"0000" when x"5B13",
			x"0000" when x"5B14",
			x"0000" when x"5B15",
			x"0000" when x"5B16",
			x"0000" when x"5B17",
			x"0000" when x"5B18",
			x"0000" when x"5B19",
			x"0000" when x"5B1A",
			x"0000" when x"5B1B",
			x"0000" when x"5B1C",
			x"0000" when x"5B1D",
			x"0000" when x"5B1E",
			x"0000" when x"5B1F",
			x"0000" when x"5B20",
			x"0000" when x"5B21",
			x"0000" when x"5B22",
			x"0000" when x"5B23",
			x"0000" when x"5B24",
			x"0000" when x"5B25",
			x"0000" when x"5B26",
			x"0000" when x"5B27",
			x"0000" when x"5B28",
			x"0000" when x"5B29",
			x"0000" when x"5B2A",
			x"0000" when x"5B2B",
			x"0000" when x"5B2C",
			x"0000" when x"5B2D",
			x"0000" when x"5B2E",
			x"0000" when x"5B2F",
			x"0000" when x"5B30",
			x"0000" when x"5B31",
			x"0000" when x"5B32",
			x"0000" when x"5B33",
			x"0000" when x"5B34",
			x"0000" when x"5B35",
			x"0000" when x"5B36",
			x"0000" when x"5B37",
			x"0000" when x"5B38",
			x"0000" when x"5B39",
			x"0000" when x"5B3A",
			x"0000" when x"5B3B",
			x"0000" when x"5B3C",
			x"0000" when x"5B3D",
			x"0000" when x"5B3E",
			x"0000" when x"5B3F",
			x"0000" when x"5B40",
			x"0000" when x"5B41",
			x"0000" when x"5B42",
			x"0000" when x"5B43",
			x"0000" when x"5B44",
			x"0000" when x"5B45",
			x"0000" when x"5B46",
			x"0000" when x"5B47",
			x"0000" when x"5B48",
			x"0000" when x"5B49",
			x"0000" when x"5B4A",
			x"0000" when x"5B4B",
			x"0000" when x"5B4C",
			x"0000" when x"5B4D",
			x"0000" when x"5B4E",
			x"0000" when x"5B4F",
			x"0000" when x"5B50",
			x"0000" when x"5B51",
			x"0000" when x"5B52",
			x"0000" when x"5B53",
			x"0000" when x"5B54",
			x"0000" when x"5B55",
			x"0000" when x"5B56",
			x"0000" when x"5B57",
			x"0000" when x"5B58",
			x"0000" when x"5B59",
			x"0000" when x"5B5A",
			x"0000" when x"5B5B",
			x"0000" when x"5B5C",
			x"0000" when x"5B5D",
			x"0000" when x"5B5E",
			x"0000" when x"5B5F",
			x"0000" when x"5B60",
			x"0000" when x"5B61",
			x"0000" when x"5B62",
			x"0000" when x"5B63",
			x"0000" when x"5B64",
			x"0000" when x"5B65",
			x"0000" when x"5B66",
			x"0000" when x"5B67",
			x"0000" when x"5B68",
			x"0000" when x"5B69",
			x"0000" when x"5B6A",
			x"0000" when x"5B6B",
			x"0000" when x"5B6C",
			x"0000" when x"5B6D",
			x"0000" when x"5B6E",
			x"0000" when x"5B6F",
			x"0000" when x"5B70",
			x"0000" when x"5B71",
			x"0000" when x"5B72",
			x"0000" when x"5B73",
			x"0000" when x"5B74",
			x"0000" when x"5B75",
			x"0000" when x"5B76",
			x"0000" when x"5B77",
			x"0000" when x"5B78",
			x"0000" when x"5B79",
			x"0000" when x"5B7A",
			x"0000" when x"5B7B",
			x"0000" when x"5B7C",
			x"0000" when x"5B7D",
			x"0000" when x"5B7E",
			x"0000" when x"5B7F",
			x"0000" when x"5B80",
			x"0000" when x"5B81",
			x"0000" when x"5B82",
			x"0000" when x"5B83",
			x"0000" when x"5B84",
			x"0000" when x"5B85",
			x"0000" when x"5B86",
			x"0000" when x"5B87",
			x"0000" when x"5B88",
			x"0000" when x"5B89",
			x"0000" when x"5B8A",
			x"0000" when x"5B8B",
			x"0000" when x"5B8C",
			x"0000" when x"5B8D",
			x"0000" when x"5B8E",
			x"0000" when x"5B8F",
			x"0000" when x"5B90",
			x"0000" when x"5B91",
			x"0000" when x"5B92",
			x"0000" when x"5B93",
			x"0000" when x"5B94",
			x"0000" when x"5B95",
			x"0000" when x"5B96",
			x"0000" when x"5B97",
			x"0000" when x"5B98",
			x"0000" when x"5B99",
			x"0000" when x"5B9A",
			x"0000" when x"5B9B",
			x"0000" when x"5B9C",
			x"0000" when x"5B9D",
			x"0000" when x"5B9E",
			x"0000" when x"5B9F",
			x"0000" when x"5BA0",
			x"0000" when x"5BA1",
			x"0000" when x"5BA2",
			x"0000" when x"5BA3",
			x"0000" when x"5BA4",
			x"0000" when x"5BA5",
			x"0000" when x"5BA6",
			x"0000" when x"5BA7",
			x"0000" when x"5BA8",
			x"0000" when x"5BA9",
			x"0000" when x"5BAA",
			x"0000" when x"5BAB",
			x"0000" when x"5BAC",
			x"0000" when x"5BAD",
			x"0000" when x"5BAE",
			x"0000" when x"5BAF",
			x"0000" when x"5BB0",
			x"0000" when x"5BB1",
			x"0000" when x"5BB2",
			x"0000" when x"5BB3",
			x"0000" when x"5BB4",
			x"0000" when x"5BB5",
			x"0000" when x"5BB6",
			x"0000" when x"5BB7",
			x"0000" when x"5BB8",
			x"0000" when x"5BB9",
			x"0000" when x"5BBA",
			x"0000" when x"5BBB",
			x"0000" when x"5BBC",
			x"0000" when x"5BBD",
			x"0000" when x"5BBE",
			x"0000" when x"5BBF",
			x"0000" when x"5BC0",
			x"0000" when x"5BC1",
			x"0000" when x"5BC2",
			x"0000" when x"5BC3",
			x"0000" when x"5BC4",
			x"0000" when x"5BC5",
			x"0000" when x"5BC6",
			x"0000" when x"5BC7",
			x"0000" when x"5BC8",
			x"0000" when x"5BC9",
			x"0000" when x"5BCA",
			x"0000" when x"5BCB",
			x"0000" when x"5BCC",
			x"0000" when x"5BCD",
			x"0000" when x"5BCE",
			x"0000" when x"5BCF",
			x"0000" when x"5BD0",
			x"0000" when x"5BD1",
			x"0000" when x"5BD2",
			x"0000" when x"5BD3",
			x"0000" when x"5BD4",
			x"0000" when x"5BD5",
			x"0000" when x"5BD6",
			x"0000" when x"5BD7",
			x"0000" when x"5BD8",
			x"0000" when x"5BD9",
			x"0000" when x"5BDA",
			x"0000" when x"5BDB",
			x"0000" when x"5BDC",
			x"0000" when x"5BDD",
			x"0000" when x"5BDE",
			x"0000" when x"5BDF",
			x"0000" when x"5BE0",
			x"0000" when x"5BE1",
			x"0000" when x"5BE2",
			x"0000" when x"5BE3",
			x"0000" when x"5BE4",
			x"0000" when x"5BE5",
			x"0000" when x"5BE6",
			x"0000" when x"5BE7",
			x"0000" when x"5BE8",
			x"0000" when x"5BE9",
			x"0000" when x"5BEA",
			x"0000" when x"5BEB",
			x"0000" when x"5BEC",
			x"0000" when x"5BED",
			x"0000" when x"5BEE",
			x"0000" when x"5BEF",
			x"0000" when x"5BF0",
			x"0000" when x"5BF1",
			x"0000" when x"5BF2",
			x"0000" when x"5BF3",
			x"0000" when x"5BF4",
			x"0000" when x"5BF5",
			x"0000" when x"5BF6",
			x"0000" when x"5BF7",
			x"0000" when x"5BF8",
			x"0000" when x"5BF9",
			x"0000" when x"5BFA",
			x"0000" when x"5BFB",
			x"0000" when x"5BFC",
			x"0000" when x"5BFD",
			x"0000" when x"5BFE",
			x"0000" when x"5BFF",
			x"0000" when x"5C00",
			x"0000" when x"5C01",
			x"0000" when x"5C02",
			x"0000" when x"5C03",
			x"0000" when x"5C04",
			x"0000" when x"5C05",
			x"0000" when x"5C06",
			x"0000" when x"5C07",
			x"0000" when x"5C08",
			x"0000" when x"5C09",
			x"0000" when x"5C0A",
			x"0000" when x"5C0B",
			x"0000" when x"5C0C",
			x"0000" when x"5C0D",
			x"0000" when x"5C0E",
			x"0000" when x"5C0F",
			x"0000" when x"5C10",
			x"0000" when x"5C11",
			x"0000" when x"5C12",
			x"0000" when x"5C13",
			x"0000" when x"5C14",
			x"0000" when x"5C15",
			x"0000" when x"5C16",
			x"0000" when x"5C17",
			x"0000" when x"5C18",
			x"0000" when x"5C19",
			x"0000" when x"5C1A",
			x"0000" when x"5C1B",
			x"0000" when x"5C1C",
			x"0000" when x"5C1D",
			x"0000" when x"5C1E",
			x"0000" when x"5C1F",
			x"0000" when x"5C20",
			x"0000" when x"5C21",
			x"0000" when x"5C22",
			x"0000" when x"5C23",
			x"0000" when x"5C24",
			x"0000" when x"5C25",
			x"0000" when x"5C26",
			x"0000" when x"5C27",
			x"0000" when x"5C28",
			x"0000" when x"5C29",
			x"0000" when x"5C2A",
			x"0000" when x"5C2B",
			x"0000" when x"5C2C",
			x"0000" when x"5C2D",
			x"0000" when x"5C2E",
			x"0000" when x"5C2F",
			x"0000" when x"5C30",
			x"0000" when x"5C31",
			x"0000" when x"5C32",
			x"0000" when x"5C33",
			x"0000" when x"5C34",
			x"0000" when x"5C35",
			x"0000" when x"5C36",
			x"0000" when x"5C37",
			x"0000" when x"5C38",
			x"0000" when x"5C39",
			x"0000" when x"5C3A",
			x"0000" when x"5C3B",
			x"0000" when x"5C3C",
			x"0000" when x"5C3D",
			x"0000" when x"5C3E",
			x"0000" when x"5C3F",
			x"0000" when x"5C40",
			x"0000" when x"5C41",
			x"0000" when x"5C42",
			x"0000" when x"5C43",
			x"0000" when x"5C44",
			x"0000" when x"5C45",
			x"0000" when x"5C46",
			x"0000" when x"5C47",
			x"0000" when x"5C48",
			x"0000" when x"5C49",
			x"0000" when x"5C4A",
			x"0000" when x"5C4B",
			x"0000" when x"5C4C",
			x"0000" when x"5C4D",
			x"0000" when x"5C4E",
			x"0000" when x"5C4F",
			x"0000" when x"5C50",
			x"0000" when x"5C51",
			x"0000" when x"5C52",
			x"0000" when x"5C53",
			x"0000" when x"5C54",
			x"0000" when x"5C55",
			x"0000" when x"5C56",
			x"0000" when x"5C57",
			x"0000" when x"5C58",
			x"0000" when x"5C59",
			x"0000" when x"5C5A",
			x"0000" when x"5C5B",
			x"0000" when x"5C5C",
			x"0000" when x"5C5D",
			x"0000" when x"5C5E",
			x"0000" when x"5C5F",
			x"0000" when x"5C60",
			x"0000" when x"5C61",
			x"0000" when x"5C62",
			x"0000" when x"5C63",
			x"0000" when x"5C64",
			x"0000" when x"5C65",
			x"0000" when x"5C66",
			x"0000" when x"5C67",
			x"0000" when x"5C68",
			x"0000" when x"5C69",
			x"0000" when x"5C6A",
			x"0000" when x"5C6B",
			x"0000" when x"5C6C",
			x"0000" when x"5C6D",
			x"0000" when x"5C6E",
			x"0000" when x"5C6F",
			x"0000" when x"5C70",
			x"0000" when x"5C71",
			x"0000" when x"5C72",
			x"0000" when x"5C73",
			x"0000" when x"5C74",
			x"0000" when x"5C75",
			x"0000" when x"5C76",
			x"0000" when x"5C77",
			x"0000" when x"5C78",
			x"0000" when x"5C79",
			x"0000" when x"5C7A",
			x"0000" when x"5C7B",
			x"0000" when x"5C7C",
			x"0000" when x"5C7D",
			x"0000" when x"5C7E",
			x"0000" when x"5C7F",
			x"0000" when x"5C80",
			x"0000" when x"5C81",
			x"0000" when x"5C82",
			x"0000" when x"5C83",
			x"0000" when x"5C84",
			x"0000" when x"5C85",
			x"0000" when x"5C86",
			x"0000" when x"5C87",
			x"0000" when x"5C88",
			x"0000" when x"5C89",
			x"0000" when x"5C8A",
			x"0000" when x"5C8B",
			x"0000" when x"5C8C",
			x"0000" when x"5C8D",
			x"0000" when x"5C8E",
			x"0000" when x"5C8F",
			x"0000" when x"5C90",
			x"0000" when x"5C91",
			x"0000" when x"5C92",
			x"0000" when x"5C93",
			x"0000" when x"5C94",
			x"0000" when x"5C95",
			x"0000" when x"5C96",
			x"0000" when x"5C97",
			x"0000" when x"5C98",
			x"0000" when x"5C99",
			x"0000" when x"5C9A",
			x"0000" when x"5C9B",
			x"0000" when x"5C9C",
			x"0000" when x"5C9D",
			x"0000" when x"5C9E",
			x"0000" when x"5C9F",
			x"0000" when x"5CA0",
			x"0000" when x"5CA1",
			x"0000" when x"5CA2",
			x"0000" when x"5CA3",
			x"0000" when x"5CA4",
			x"0000" when x"5CA5",
			x"0000" when x"5CA6",
			x"0000" when x"5CA7",
			x"0000" when x"5CA8",
			x"0000" when x"5CA9",
			x"0000" when x"5CAA",
			x"0000" when x"5CAB",
			x"0000" when x"5CAC",
			x"0000" when x"5CAD",
			x"0000" when x"5CAE",
			x"0000" when x"5CAF",
			x"0000" when x"5CB0",
			x"0000" when x"5CB1",
			x"0000" when x"5CB2",
			x"0000" when x"5CB3",
			x"0000" when x"5CB4",
			x"0000" when x"5CB5",
			x"0000" when x"5CB6",
			x"0000" when x"5CB7",
			x"0000" when x"5CB8",
			x"0000" when x"5CB9",
			x"0000" when x"5CBA",
			x"0000" when x"5CBB",
			x"0000" when x"5CBC",
			x"0000" when x"5CBD",
			x"0000" when x"5CBE",
			x"0000" when x"5CBF",
			x"0000" when x"5CC0",
			x"0000" when x"5CC1",
			x"0000" when x"5CC2",
			x"0000" when x"5CC3",
			x"0000" when x"5CC4",
			x"0000" when x"5CC5",
			x"0000" when x"5CC6",
			x"0000" when x"5CC7",
			x"0000" when x"5CC8",
			x"0000" when x"5CC9",
			x"0000" when x"5CCA",
			x"0000" when x"5CCB",
			x"0000" when x"5CCC",
			x"0000" when x"5CCD",
			x"0000" when x"5CCE",
			x"0000" when x"5CCF",
			x"0000" when x"5CD0",
			x"0000" when x"5CD1",
			x"0000" when x"5CD2",
			x"0000" when x"5CD3",
			x"0000" when x"5CD4",
			x"0000" when x"5CD5",
			x"0000" when x"5CD6",
			x"0000" when x"5CD7",
			x"0000" when x"5CD8",
			x"0000" when x"5CD9",
			x"0000" when x"5CDA",
			x"0000" when x"5CDB",
			x"0000" when x"5CDC",
			x"0000" when x"5CDD",
			x"0000" when x"5CDE",
			x"0000" when x"5CDF",
			x"0000" when x"5CE0",
			x"0000" when x"5CE1",
			x"0000" when x"5CE2",
			x"0000" when x"5CE3",
			x"0000" when x"5CE4",
			x"0000" when x"5CE5",
			x"0000" when x"5CE6",
			x"0000" when x"5CE7",
			x"0000" when x"5CE8",
			x"0000" when x"5CE9",
			x"0000" when x"5CEA",
			x"0000" when x"5CEB",
			x"0000" when x"5CEC",
			x"0000" when x"5CED",
			x"0000" when x"5CEE",
			x"0000" when x"5CEF",
			x"0000" when x"5CF0",
			x"0000" when x"5CF1",
			x"0000" when x"5CF2",
			x"0000" when x"5CF3",
			x"0000" when x"5CF4",
			x"0000" when x"5CF5",
			x"0000" when x"5CF6",
			x"0000" when x"5CF7",
			x"0000" when x"5CF8",
			x"0000" when x"5CF9",
			x"0000" when x"5CFA",
			x"0000" when x"5CFB",
			x"0000" when x"5CFC",
			x"0000" when x"5CFD",
			x"0000" when x"5CFE",
			x"0000" when x"5CFF",
			x"0000" when x"5D00",
			x"0000" when x"5D01",
			x"0000" when x"5D02",
			x"0000" when x"5D03",
			x"0000" when x"5D04",
			x"0000" when x"5D05",
			x"0000" when x"5D06",
			x"0000" when x"5D07",
			x"0000" when x"5D08",
			x"0000" when x"5D09",
			x"0000" when x"5D0A",
			x"0000" when x"5D0B",
			x"0000" when x"5D0C",
			x"0000" when x"5D0D",
			x"0000" when x"5D0E",
			x"0000" when x"5D0F",
			x"0000" when x"5D10",
			x"0000" when x"5D11",
			x"0000" when x"5D12",
			x"0000" when x"5D13",
			x"0000" when x"5D14",
			x"0000" when x"5D15",
			x"0000" when x"5D16",
			x"0000" when x"5D17",
			x"0000" when x"5D18",
			x"0000" when x"5D19",
			x"0000" when x"5D1A",
			x"0000" when x"5D1B",
			x"0000" when x"5D1C",
			x"0000" when x"5D1D",
			x"0000" when x"5D1E",
			x"0000" when x"5D1F",
			x"0000" when x"5D20",
			x"0000" when x"5D21",
			x"0000" when x"5D22",
			x"0000" when x"5D23",
			x"0000" when x"5D24",
			x"0000" when x"5D25",
			x"0000" when x"5D26",
			x"0000" when x"5D27",
			x"0000" when x"5D28",
			x"0000" when x"5D29",
			x"0000" when x"5D2A",
			x"0000" when x"5D2B",
			x"0000" when x"5D2C",
			x"0000" when x"5D2D",
			x"0000" when x"5D2E",
			x"0000" when x"5D2F",
			x"0000" when x"5D30",
			x"0000" when x"5D31",
			x"0000" when x"5D32",
			x"0000" when x"5D33",
			x"0000" when x"5D34",
			x"0000" when x"5D35",
			x"0000" when x"5D36",
			x"0000" when x"5D37",
			x"0000" when x"5D38",
			x"0000" when x"5D39",
			x"0000" when x"5D3A",
			x"0000" when x"5D3B",
			x"0000" when x"5D3C",
			x"0000" when x"5D3D",
			x"0000" when x"5D3E",
			x"0000" when x"5D3F",
			x"0000" when x"5D40",
			x"0000" when x"5D41",
			x"0000" when x"5D42",
			x"0000" when x"5D43",
			x"0000" when x"5D44",
			x"0000" when x"5D45",
			x"0000" when x"5D46",
			x"0000" when x"5D47",
			x"0000" when x"5D48",
			x"0000" when x"5D49",
			x"0000" when x"5D4A",
			x"0000" when x"5D4B",
			x"0000" when x"5D4C",
			x"0000" when x"5D4D",
			x"0000" when x"5D4E",
			x"0000" when x"5D4F",
			x"0000" when x"5D50",
			x"0000" when x"5D51",
			x"0000" when x"5D52",
			x"0000" when x"5D53",
			x"0000" when x"5D54",
			x"0000" when x"5D55",
			x"0000" when x"5D56",
			x"0000" when x"5D57",
			x"0000" when x"5D58",
			x"0000" when x"5D59",
			x"0000" when x"5D5A",
			x"0000" when x"5D5B",
			x"0000" when x"5D5C",
			x"0000" when x"5D5D",
			x"0000" when x"5D5E",
			x"0000" when x"5D5F",
			x"0000" when x"5D60",
			x"0000" when x"5D61",
			x"0000" when x"5D62",
			x"0000" when x"5D63",
			x"0000" when x"5D64",
			x"0000" when x"5D65",
			x"0000" when x"5D66",
			x"0000" when x"5D67",
			x"0000" when x"5D68",
			x"0000" when x"5D69",
			x"0000" when x"5D6A",
			x"0000" when x"5D6B",
			x"0000" when x"5D6C",
			x"0000" when x"5D6D",
			x"0000" when x"5D6E",
			x"0000" when x"5D6F",
			x"0000" when x"5D70",
			x"0000" when x"5D71",
			x"0000" when x"5D72",
			x"0000" when x"5D73",
			x"0000" when x"5D74",
			x"0000" when x"5D75",
			x"0000" when x"5D76",
			x"0000" when x"5D77",
			x"0000" when x"5D78",
			x"0000" when x"5D79",
			x"0000" when x"5D7A",
			x"0000" when x"5D7B",
			x"0000" when x"5D7C",
			x"0000" when x"5D7D",
			x"0000" when x"5D7E",
			x"0000" when x"5D7F",
			x"0000" when x"5D80",
			x"0000" when x"5D81",
			x"0000" when x"5D82",
			x"0000" when x"5D83",
			x"0000" when x"5D84",
			x"0000" when x"5D85",
			x"0000" when x"5D86",
			x"0000" when x"5D87",
			x"0000" when x"5D88",
			x"0000" when x"5D89",
			x"0000" when x"5D8A",
			x"0000" when x"5D8B",
			x"0000" when x"5D8C",
			x"0000" when x"5D8D",
			x"0000" when x"5D8E",
			x"0000" when x"5D8F",
			x"0000" when x"5D90",
			x"0000" when x"5D91",
			x"0000" when x"5D92",
			x"0000" when x"5D93",
			x"0000" when x"5D94",
			x"0000" when x"5D95",
			x"0000" when x"5D96",
			x"0000" when x"5D97",
			x"0000" when x"5D98",
			x"0000" when x"5D99",
			x"0000" when x"5D9A",
			x"0000" when x"5D9B",
			x"0000" when x"5D9C",
			x"0000" when x"5D9D",
			x"0000" when x"5D9E",
			x"0000" when x"5D9F",
			x"0000" when x"5DA0",
			x"0000" when x"5DA1",
			x"0000" when x"5DA2",
			x"0000" when x"5DA3",
			x"0000" when x"5DA4",
			x"0000" when x"5DA5",
			x"0000" when x"5DA6",
			x"0000" when x"5DA7",
			x"0000" when x"5DA8",
			x"0000" when x"5DA9",
			x"0000" when x"5DAA",
			x"0000" when x"5DAB",
			x"0000" when x"5DAC",
			x"0000" when x"5DAD",
			x"0000" when x"5DAE",
			x"0000" when x"5DAF",
			x"0000" when x"5DB0",
			x"0000" when x"5DB1",
			x"0000" when x"5DB2",
			x"0000" when x"5DB3",
			x"0000" when x"5DB4",
			x"0000" when x"5DB5",
			x"0000" when x"5DB6",
			x"0000" when x"5DB7",
			x"0000" when x"5DB8",
			x"0000" when x"5DB9",
			x"0000" when x"5DBA",
			x"0000" when x"5DBB",
			x"0000" when x"5DBC",
			x"0000" when x"5DBD",
			x"0000" when x"5DBE",
			x"0000" when x"5DBF",
			x"0000" when x"5DC0",
			x"0000" when x"5DC1",
			x"0000" when x"5DC2",
			x"0000" when x"5DC3",
			x"0000" when x"5DC4",
			x"0000" when x"5DC5",
			x"0000" when x"5DC6",
			x"0000" when x"5DC7",
			x"0000" when x"5DC8",
			x"0000" when x"5DC9",
			x"0000" when x"5DCA",
			x"0000" when x"5DCB",
			x"0000" when x"5DCC",
			x"0000" when x"5DCD",
			x"0000" when x"5DCE",
			x"0000" when x"5DCF",
			x"0000" when x"5DD0",
			x"0000" when x"5DD1",
			x"0000" when x"5DD2",
			x"0000" when x"5DD3",
			x"0000" when x"5DD4",
			x"0000" when x"5DD5",
			x"0000" when x"5DD6",
			x"0000" when x"5DD7",
			x"0000" when x"5DD8",
			x"0000" when x"5DD9",
			x"0000" when x"5DDA",
			x"0000" when x"5DDB",
			x"0000" when x"5DDC",
			x"0000" when x"5DDD",
			x"0000" when x"5DDE",
			x"0000" when x"5DDF",
			x"0000" when x"5DE0",
			x"0000" when x"5DE1",
			x"0000" when x"5DE2",
			x"0000" when x"5DE3",
			x"0000" when x"5DE4",
			x"0000" when x"5DE5",
			x"0000" when x"5DE6",
			x"0000" when x"5DE7",
			x"0000" when x"5DE8",
			x"0000" when x"5DE9",
			x"0000" when x"5DEA",
			x"0000" when x"5DEB",
			x"0000" when x"5DEC",
			x"0000" when x"5DED",
			x"0000" when x"5DEE",
			x"0000" when x"5DEF",
			x"0000" when x"5DF0",
			x"0000" when x"5DF1",
			x"0000" when x"5DF2",
			x"0000" when x"5DF3",
			x"0000" when x"5DF4",
			x"0000" when x"5DF5",
			x"0000" when x"5DF6",
			x"0000" when x"5DF7",
			x"0000" when x"5DF8",
			x"0000" when x"5DF9",
			x"0000" when x"5DFA",
			x"0000" when x"5DFB",
			x"0000" when x"5DFC",
			x"0000" when x"5DFD",
			x"0000" when x"5DFE",
			x"0000" when x"5DFF",
			x"0000" when x"5E00",
			x"0000" when x"5E01",
			x"0000" when x"5E02",
			x"0000" when x"5E03",
			x"0000" when x"5E04",
			x"0000" when x"5E05",
			x"0000" when x"5E06",
			x"0000" when x"5E07",
			x"0000" when x"5E08",
			x"0000" when x"5E09",
			x"0000" when x"5E0A",
			x"0000" when x"5E0B",
			x"0000" when x"5E0C",
			x"0000" when x"5E0D",
			x"0000" when x"5E0E",
			x"0000" when x"5E0F",
			x"0000" when x"5E10",
			x"0000" when x"5E11",
			x"0000" when x"5E12",
			x"0000" when x"5E13",
			x"0000" when x"5E14",
			x"0000" when x"5E15",
			x"0000" when x"5E16",
			x"0000" when x"5E17",
			x"0000" when x"5E18",
			x"0000" when x"5E19",
			x"0000" when x"5E1A",
			x"0000" when x"5E1B",
			x"0000" when x"5E1C",
			x"0000" when x"5E1D",
			x"0000" when x"5E1E",
			x"0000" when x"5E1F",
			x"0000" when x"5E20",
			x"0000" when x"5E21",
			x"0000" when x"5E22",
			x"0000" when x"5E23",
			x"0000" when x"5E24",
			x"0000" when x"5E25",
			x"0000" when x"5E26",
			x"0000" when x"5E27",
			x"0000" when x"5E28",
			x"0000" when x"5E29",
			x"0000" when x"5E2A",
			x"0000" when x"5E2B",
			x"0000" when x"5E2C",
			x"0000" when x"5E2D",
			x"0000" when x"5E2E",
			x"0000" when x"5E2F",
			x"0000" when x"5E30",
			x"0000" when x"5E31",
			x"0000" when x"5E32",
			x"0000" when x"5E33",
			x"0000" when x"5E34",
			x"0000" when x"5E35",
			x"0000" when x"5E36",
			x"0000" when x"5E37",
			x"0000" when x"5E38",
			x"0000" when x"5E39",
			x"0000" when x"5E3A",
			x"0000" when x"5E3B",
			x"0000" when x"5E3C",
			x"0000" when x"5E3D",
			x"0000" when x"5E3E",
			x"0000" when x"5E3F",
			x"0000" when x"5E40",
			x"0000" when x"5E41",
			x"0000" when x"5E42",
			x"0000" when x"5E43",
			x"0000" when x"5E44",
			x"0000" when x"5E45",
			x"0000" when x"5E46",
			x"0000" when x"5E47",
			x"0000" when x"5E48",
			x"0000" when x"5E49",
			x"0000" when x"5E4A",
			x"0000" when x"5E4B",
			x"0000" when x"5E4C",
			x"0000" when x"5E4D",
			x"0000" when x"5E4E",
			x"0000" when x"5E4F",
			x"0000" when x"5E50",
			x"0000" when x"5E51",
			x"0000" when x"5E52",
			x"0000" when x"5E53",
			x"0000" when x"5E54",
			x"0000" when x"5E55",
			x"0000" when x"5E56",
			x"0000" when x"5E57",
			x"0000" when x"5E58",
			x"0000" when x"5E59",
			x"0000" when x"5E5A",
			x"0000" when x"5E5B",
			x"0000" when x"5E5C",
			x"0000" when x"5E5D",
			x"0000" when x"5E5E",
			x"0000" when x"5E5F",
			x"0000" when x"5E60",
			x"0000" when x"5E61",
			x"0000" when x"5E62",
			x"0000" when x"5E63",
			x"0000" when x"5E64",
			x"0000" when x"5E65",
			x"0000" when x"5E66",
			x"0000" when x"5E67",
			x"0000" when x"5E68",
			x"0000" when x"5E69",
			x"0000" when x"5E6A",
			x"0000" when x"5E6B",
			x"0000" when x"5E6C",
			x"0000" when x"5E6D",
			x"0000" when x"5E6E",
			x"0000" when x"5E6F",
			x"0000" when x"5E70",
			x"0000" when x"5E71",
			x"0000" when x"5E72",
			x"0000" when x"5E73",
			x"0000" when x"5E74",
			x"0000" when x"5E75",
			x"0000" when x"5E76",
			x"0000" when x"5E77",
			x"0000" when x"5E78",
			x"0000" when x"5E79",
			x"0000" when x"5E7A",
			x"0000" when x"5E7B",
			x"0000" when x"5E7C",
			x"0000" when x"5E7D",
			x"0000" when x"5E7E",
			x"0000" when x"5E7F",
			x"0000" when x"5E80",
			x"0000" when x"5E81",
			x"0000" when x"5E82",
			x"0000" when x"5E83",
			x"0000" when x"5E84",
			x"0000" when x"5E85",
			x"0000" when x"5E86",
			x"0000" when x"5E87",
			x"0000" when x"5E88",
			x"0000" when x"5E89",
			x"0000" when x"5E8A",
			x"0000" when x"5E8B",
			x"0000" when x"5E8C",
			x"0000" when x"5E8D",
			x"0000" when x"5E8E",
			x"0000" when x"5E8F",
			x"0000" when x"5E90",
			x"0000" when x"5E91",
			x"0000" when x"5E92",
			x"0000" when x"5E93",
			x"0000" when x"5E94",
			x"0000" when x"5E95",
			x"0000" when x"5E96",
			x"0000" when x"5E97",
			x"0000" when x"5E98",
			x"0000" when x"5E99",
			x"0000" when x"5E9A",
			x"0000" when x"5E9B",
			x"0000" when x"5E9C",
			x"0000" when x"5E9D",
			x"0000" when x"5E9E",
			x"0000" when x"5E9F",
			x"0000" when x"5EA0",
			x"0000" when x"5EA1",
			x"0000" when x"5EA2",
			x"0000" when x"5EA3",
			x"0000" when x"5EA4",
			x"0000" when x"5EA5",
			x"0000" when x"5EA6",
			x"0000" when x"5EA7",
			x"0000" when x"5EA8",
			x"0000" when x"5EA9",
			x"0000" when x"5EAA",
			x"0000" when x"5EAB",
			x"0000" when x"5EAC",
			x"0000" when x"5EAD",
			x"0000" when x"5EAE",
			x"0000" when x"5EAF",
			x"0000" when x"5EB0",
			x"0000" when x"5EB1",
			x"0000" when x"5EB2",
			x"0000" when x"5EB3",
			x"0000" when x"5EB4",
			x"0000" when x"5EB5",
			x"0000" when x"5EB6",
			x"0000" when x"5EB7",
			x"0000" when x"5EB8",
			x"0000" when x"5EB9",
			x"0000" when x"5EBA",
			x"0000" when x"5EBB",
			x"0000" when x"5EBC",
			x"0000" when x"5EBD",
			x"0000" when x"5EBE",
			x"0000" when x"5EBF",
			x"0000" when x"5EC0",
			x"0000" when x"5EC1",
			x"0000" when x"5EC2",
			x"0000" when x"5EC3",
			x"0000" when x"5EC4",
			x"0000" when x"5EC5",
			x"0000" when x"5EC6",
			x"0000" when x"5EC7",
			x"0000" when x"5EC8",
			x"0000" when x"5EC9",
			x"0000" when x"5ECA",
			x"0000" when x"5ECB",
			x"0000" when x"5ECC",
			x"0000" when x"5ECD",
			x"0000" when x"5ECE",
			x"0000" when x"5ECF",
			x"0000" when x"5ED0",
			x"0000" when x"5ED1",
			x"0000" when x"5ED2",
			x"0000" when x"5ED3",
			x"0000" when x"5ED4",
			x"0000" when x"5ED5",
			x"0000" when x"5ED6",
			x"0000" when x"5ED7",
			x"0000" when x"5ED8",
			x"0000" when x"5ED9",
			x"0000" when x"5EDA",
			x"0000" when x"5EDB",
			x"0000" when x"5EDC",
			x"0000" when x"5EDD",
			x"0000" when x"5EDE",
			x"0000" when x"5EDF",
			x"0000" when x"5EE0",
			x"0000" when x"5EE1",
			x"0000" when x"5EE2",
			x"0000" when x"5EE3",
			x"0000" when x"5EE4",
			x"0000" when x"5EE5",
			x"0000" when x"5EE6",
			x"0000" when x"5EE7",
			x"0000" when x"5EE8",
			x"0000" when x"5EE9",
			x"0000" when x"5EEA",
			x"0000" when x"5EEB",
			x"0000" when x"5EEC",
			x"0000" when x"5EED",
			x"0000" when x"5EEE",
			x"0000" when x"5EEF",
			x"0000" when x"5EF0",
			x"0000" when x"5EF1",
			x"0000" when x"5EF2",
			x"0000" when x"5EF3",
			x"0000" when x"5EF4",
			x"0000" when x"5EF5",
			x"0000" when x"5EF6",
			x"0000" when x"5EF7",
			x"0000" when x"5EF8",
			x"0000" when x"5EF9",
			x"0000" when x"5EFA",
			x"0000" when x"5EFB",
			x"0000" when x"5EFC",
			x"0000" when x"5EFD",
			x"0000" when x"5EFE",
			x"0000" when x"5EFF",
			x"0000" when x"5F00",
			x"0000" when x"5F01",
			x"0000" when x"5F02",
			x"0000" when x"5F03",
			x"0000" when x"5F04",
			x"0000" when x"5F05",
			x"0000" when x"5F06",
			x"0000" when x"5F07",
			x"0000" when x"5F08",
			x"0000" when x"5F09",
			x"0000" when x"5F0A",
			x"0000" when x"5F0B",
			x"0000" when x"5F0C",
			x"0000" when x"5F0D",
			x"0000" when x"5F0E",
			x"0000" when x"5F0F",
			x"0000" when x"5F10",
			x"0000" when x"5F11",
			x"0000" when x"5F12",
			x"0000" when x"5F13",
			x"0000" when x"5F14",
			x"0000" when x"5F15",
			x"0000" when x"5F16",
			x"0000" when x"5F17",
			x"0000" when x"5F18",
			x"0000" when x"5F19",
			x"0000" when x"5F1A",
			x"0000" when x"5F1B",
			x"0000" when x"5F1C",
			x"0000" when x"5F1D",
			x"0000" when x"5F1E",
			x"0000" when x"5F1F",
			x"0000" when x"5F20",
			x"0000" when x"5F21",
			x"0000" when x"5F22",
			x"0000" when x"5F23",
			x"0000" when x"5F24",
			x"0000" when x"5F25",
			x"0000" when x"5F26",
			x"0000" when x"5F27",
			x"0000" when x"5F28",
			x"0000" when x"5F29",
			x"0000" when x"5F2A",
			x"0000" when x"5F2B",
			x"0000" when x"5F2C",
			x"0000" when x"5F2D",
			x"0000" when x"5F2E",
			x"0000" when x"5F2F",
			x"0000" when x"5F30",
			x"0000" when x"5F31",
			x"0000" when x"5F32",
			x"0000" when x"5F33",
			x"0000" when x"5F34",
			x"0000" when x"5F35",
			x"0000" when x"5F36",
			x"0000" when x"5F37",
			x"0000" when x"5F38",
			x"0000" when x"5F39",
			x"0000" when x"5F3A",
			x"0000" when x"5F3B",
			x"0000" when x"5F3C",
			x"0000" when x"5F3D",
			x"0000" when x"5F3E",
			x"0000" when x"5F3F",
			x"0000" when x"5F40",
			x"0000" when x"5F41",
			x"0000" when x"5F42",
			x"0000" when x"5F43",
			x"0000" when x"5F44",
			x"0000" when x"5F45",
			x"0000" when x"5F46",
			x"0000" when x"5F47",
			x"0000" when x"5F48",
			x"0000" when x"5F49",
			x"0000" when x"5F4A",
			x"0000" when x"5F4B",
			x"0000" when x"5F4C",
			x"0000" when x"5F4D",
			x"0000" when x"5F4E",
			x"0000" when x"5F4F",
			x"0000" when x"5F50",
			x"0000" when x"5F51",
			x"0000" when x"5F52",
			x"0000" when x"5F53",
			x"0000" when x"5F54",
			x"0000" when x"5F55",
			x"0000" when x"5F56",
			x"0000" when x"5F57",
			x"0000" when x"5F58",
			x"0000" when x"5F59",
			x"0000" when x"5F5A",
			x"0000" when x"5F5B",
			x"0000" when x"5F5C",
			x"0000" when x"5F5D",
			x"0000" when x"5F5E",
			x"0000" when x"5F5F",
			x"0000" when x"5F60",
			x"0000" when x"5F61",
			x"0000" when x"5F62",
			x"0000" when x"5F63",
			x"0000" when x"5F64",
			x"0000" when x"5F65",
			x"0000" when x"5F66",
			x"0000" when x"5F67",
			x"0000" when x"5F68",
			x"0000" when x"5F69",
			x"0000" when x"5F6A",
			x"0000" when x"5F6B",
			x"0000" when x"5F6C",
			x"0000" when x"5F6D",
			x"0000" when x"5F6E",
			x"0000" when x"5F6F",
			x"0000" when x"5F70",
			x"0000" when x"5F71",
			x"0000" when x"5F72",
			x"0000" when x"5F73",
			x"0000" when x"5F74",
			x"0000" when x"5F75",
			x"0000" when x"5F76",
			x"0000" when x"5F77",
			x"0000" when x"5F78",
			x"0000" when x"5F79",
			x"0000" when x"5F7A",
			x"0000" when x"5F7B",
			x"0000" when x"5F7C",
			x"0000" when x"5F7D",
			x"0000" when x"5F7E",
			x"0000" when x"5F7F",
			x"0000" when x"5F80",
			x"0000" when x"5F81",
			x"0000" when x"5F82",
			x"0000" when x"5F83",
			x"0000" when x"5F84",
			x"0000" when x"5F85",
			x"0000" when x"5F86",
			x"0000" when x"5F87",
			x"0000" when x"5F88",
			x"0000" when x"5F89",
			x"0000" when x"5F8A",
			x"0000" when x"5F8B",
			x"0000" when x"5F8C",
			x"0000" when x"5F8D",
			x"0000" when x"5F8E",
			x"0000" when x"5F8F",
			x"0000" when x"5F90",
			x"0000" when x"5F91",
			x"0000" when x"5F92",
			x"0000" when x"5F93",
			x"0000" when x"5F94",
			x"0000" when x"5F95",
			x"0000" when x"5F96",
			x"0000" when x"5F97",
			x"0000" when x"5F98",
			x"0000" when x"5F99",
			x"0000" when x"5F9A",
			x"0000" when x"5F9B",
			x"0000" when x"5F9C",
			x"0000" when x"5F9D",
			x"0000" when x"5F9E",
			x"0000" when x"5F9F",
			x"0000" when x"5FA0",
			x"0000" when x"5FA1",
			x"0000" when x"5FA2",
			x"0000" when x"5FA3",
			x"0000" when x"5FA4",
			x"0000" when x"5FA5",
			x"0000" when x"5FA6",
			x"0000" when x"5FA7",
			x"0000" when x"5FA8",
			x"0000" when x"5FA9",
			x"0000" when x"5FAA",
			x"0000" when x"5FAB",
			x"0000" when x"5FAC",
			x"0000" when x"5FAD",
			x"0000" when x"5FAE",
			x"0000" when x"5FAF",
			x"0000" when x"5FB0",
			x"0000" when x"5FB1",
			x"0000" when x"5FB2",
			x"0000" when x"5FB3",
			x"0000" when x"5FB4",
			x"0000" when x"5FB5",
			x"0000" when x"5FB6",
			x"0000" when x"5FB7",
			x"0000" when x"5FB8",
			x"0000" when x"5FB9",
			x"0000" when x"5FBA",
			x"0000" when x"5FBB",
			x"0000" when x"5FBC",
			x"0000" when x"5FBD",
			x"0000" when x"5FBE",
			x"0000" when x"5FBF",
			x"0000" when x"5FC0",
			x"0000" when x"5FC1",
			x"0000" when x"5FC2",
			x"0000" when x"5FC3",
			x"0000" when x"5FC4",
			x"0000" when x"5FC5",
			x"0000" when x"5FC6",
			x"0000" when x"5FC7",
			x"0000" when x"5FC8",
			x"0000" when x"5FC9",
			x"0000" when x"5FCA",
			x"0000" when x"5FCB",
			x"0000" when x"5FCC",
			x"0000" when x"5FCD",
			x"0000" when x"5FCE",
			x"0000" when x"5FCF",
			x"0000" when x"5FD0",
			x"0000" when x"5FD1",
			x"0000" when x"5FD2",
			x"0000" when x"5FD3",
			x"0000" when x"5FD4",
			x"0000" when x"5FD5",
			x"0000" when x"5FD6",
			x"0000" when x"5FD7",
			x"0000" when x"5FD8",
			x"0000" when x"5FD9",
			x"0000" when x"5FDA",
			x"0000" when x"5FDB",
			x"0000" when x"5FDC",
			x"0000" when x"5FDD",
			x"0000" when x"5FDE",
			x"0000" when x"5FDF",
			x"0000" when x"5FE0",
			x"0000" when x"5FE1",
			x"0000" when x"5FE2",
			x"0000" when x"5FE3",
			x"0000" when x"5FE4",
			x"0000" when x"5FE5",
			x"0000" when x"5FE6",
			x"0000" when x"5FE7",
			x"0000" when x"5FE8",
			x"0000" when x"5FE9",
			x"0000" when x"5FEA",
			x"0000" when x"5FEB",
			x"0000" when x"5FEC",
			x"0000" when x"5FED",
			x"0000" when x"5FEE",
			x"0000" when x"5FEF",
			x"0000" when x"5FF0",
			x"0000" when x"5FF1",
			x"0000" when x"5FF2",
			x"0000" when x"5FF3",
			x"0000" when x"5FF4",
			x"0000" when x"5FF5",
			x"0000" when x"5FF6",
			x"0000" when x"5FF7",
			x"0000" when x"5FF8",
			x"0000" when x"5FF9",
			x"0000" when x"5FFA",
			x"0000" when x"5FFB",
			x"0000" when x"5FFC",
			x"0000" when x"5FFD",
			x"0000" when x"5FFE",
			x"0000" when x"5FFF",
			x"0000" when x"6000",
			x"0000" when x"6001",
			x"0000" when x"6002",
			x"0000" when x"6003",
			x"0000" when x"6004",
			x"0000" when x"6005",
			x"0000" when x"6006",
			x"0000" when x"6007",
			x"0000" when x"6008",
			x"0000" when x"6009",
			x"0000" when x"600A",
			x"0000" when x"600B",
			x"0000" when x"600C",
			x"0000" when x"600D",
			x"0000" when x"600E",
			x"0000" when x"600F",
			x"0000" when x"6010",
			x"0000" when x"6011",
			x"0000" when x"6012",
			x"0000" when x"6013",
			x"0000" when x"6014",
			x"0000" when x"6015",
			x"0000" when x"6016",
			x"0000" when x"6017",
			x"0000" when x"6018",
			x"0000" when x"6019",
			x"0000" when x"601A",
			x"0000" when x"601B",
			x"0000" when x"601C",
			x"0000" when x"601D",
			x"0000" when x"601E",
			x"0000" when x"601F",
			x"0000" when x"6020",
			x"0000" when x"6021",
			x"0000" when x"6022",
			x"0000" when x"6023",
			x"0000" when x"6024",
			x"0000" when x"6025",
			x"0000" when x"6026",
			x"0000" when x"6027",
			x"0000" when x"6028",
			x"0000" when x"6029",
			x"0000" when x"602A",
			x"0000" when x"602B",
			x"0000" when x"602C",
			x"0000" when x"602D",
			x"0000" when x"602E",
			x"0000" when x"602F",
			x"0000" when x"6030",
			x"0000" when x"6031",
			x"0000" when x"6032",
			x"0000" when x"6033",
			x"0000" when x"6034",
			x"0000" when x"6035",
			x"0000" when x"6036",
			x"0000" when x"6037",
			x"0000" when x"6038",
			x"0000" when x"6039",
			x"0000" when x"603A",
			x"0000" when x"603B",
			x"0000" when x"603C",
			x"0000" when x"603D",
			x"0000" when x"603E",
			x"0000" when x"603F",
			x"0000" when x"6040",
			x"0000" when x"6041",
			x"0000" when x"6042",
			x"0000" when x"6043",
			x"0000" when x"6044",
			x"0000" when x"6045",
			x"0000" when x"6046",
			x"0000" when x"6047",
			x"0000" when x"6048",
			x"0000" when x"6049",
			x"0000" when x"604A",
			x"0000" when x"604B",
			x"0000" when x"604C",
			x"0000" when x"604D",
			x"0000" when x"604E",
			x"0000" when x"604F",
			x"0000" when x"6050",
			x"0000" when x"6051",
			x"0000" when x"6052",
			x"0000" when x"6053",
			x"0000" when x"6054",
			x"0000" when x"6055",
			x"0000" when x"6056",
			x"0000" when x"6057",
			x"0000" when x"6058",
			x"0000" when x"6059",
			x"0000" when x"605A",
			x"0000" when x"605B",
			x"0000" when x"605C",
			x"0000" when x"605D",
			x"0000" when x"605E",
			x"0000" when x"605F",
			x"0000" when x"6060",
			x"0000" when x"6061",
			x"0000" when x"6062",
			x"0000" when x"6063",
			x"0000" when x"6064",
			x"0000" when x"6065",
			x"0000" when x"6066",
			x"0000" when x"6067",
			x"0000" when x"6068",
			x"0000" when x"6069",
			x"0000" when x"606A",
			x"0000" when x"606B",
			x"0000" when x"606C",
			x"0000" when x"606D",
			x"0000" when x"606E",
			x"0000" when x"606F",
			x"0000" when x"6070",
			x"0000" when x"6071",
			x"0000" when x"6072",
			x"0000" when x"6073",
			x"0000" when x"6074",
			x"0000" when x"6075",
			x"0000" when x"6076",
			x"0000" when x"6077",
			x"0000" when x"6078",
			x"0000" when x"6079",
			x"0000" when x"607A",
			x"0000" when x"607B",
			x"0000" when x"607C",
			x"0000" when x"607D",
			x"0000" when x"607E",
			x"0000" when x"607F",
			x"0000" when x"6080",
			x"0000" when x"6081",
			x"0000" when x"6082",
			x"0000" when x"6083",
			x"0000" when x"6084",
			x"0000" when x"6085",
			x"0000" when x"6086",
			x"0000" when x"6087",
			x"0000" when x"6088",
			x"0000" when x"6089",
			x"0000" when x"608A",
			x"0000" when x"608B",
			x"0000" when x"608C",
			x"0000" when x"608D",
			x"0000" when x"608E",
			x"0000" when x"608F",
			x"0000" when x"6090",
			x"0000" when x"6091",
			x"0000" when x"6092",
			x"0000" when x"6093",
			x"0000" when x"6094",
			x"0000" when x"6095",
			x"0000" when x"6096",
			x"0000" when x"6097",
			x"0000" when x"6098",
			x"0000" when x"6099",
			x"0000" when x"609A",
			x"0000" when x"609B",
			x"0000" when x"609C",
			x"0000" when x"609D",
			x"0000" when x"609E",
			x"0000" when x"609F",
			x"0000" when x"60A0",
			x"0000" when x"60A1",
			x"0000" when x"60A2",
			x"0000" when x"60A3",
			x"0000" when x"60A4",
			x"0000" when x"60A5",
			x"0000" when x"60A6",
			x"0000" when x"60A7",
			x"0000" when x"60A8",
			x"0000" when x"60A9",
			x"0000" when x"60AA",
			x"0000" when x"60AB",
			x"0000" when x"60AC",
			x"0000" when x"60AD",
			x"0000" when x"60AE",
			x"0000" when x"60AF",
			x"0000" when x"60B0",
			x"0000" when x"60B1",
			x"0000" when x"60B2",
			x"0000" when x"60B3",
			x"0000" when x"60B4",
			x"0000" when x"60B5",
			x"0000" when x"60B6",
			x"0000" when x"60B7",
			x"0000" when x"60B8",
			x"0000" when x"60B9",
			x"0000" when x"60BA",
			x"0000" when x"60BB",
			x"0000" when x"60BC",
			x"0000" when x"60BD",
			x"0000" when x"60BE",
			x"0000" when x"60BF",
			x"0000" when x"60C0",
			x"0000" when x"60C1",
			x"0000" when x"60C2",
			x"0000" when x"60C3",
			x"0000" when x"60C4",
			x"0000" when x"60C5",
			x"0000" when x"60C6",
			x"0000" when x"60C7",
			x"0000" when x"60C8",
			x"0000" when x"60C9",
			x"0000" when x"60CA",
			x"0000" when x"60CB",
			x"0000" when x"60CC",
			x"0000" when x"60CD",
			x"0000" when x"60CE",
			x"0000" when x"60CF",
			x"0000" when x"60D0",
			x"0000" when x"60D1",
			x"0000" when x"60D2",
			x"0000" when x"60D3",
			x"0000" when x"60D4",
			x"0000" when x"60D5",
			x"0000" when x"60D6",
			x"0000" when x"60D7",
			x"0000" when x"60D8",
			x"0000" when x"60D9",
			x"0000" when x"60DA",
			x"0000" when x"60DB",
			x"0000" when x"60DC",
			x"0000" when x"60DD",
			x"0000" when x"60DE",
			x"0000" when x"60DF",
			x"0000" when x"60E0",
			x"0000" when x"60E1",
			x"0000" when x"60E2",
			x"0000" when x"60E3",
			x"0000" when x"60E4",
			x"0000" when x"60E5",
			x"0000" when x"60E6",
			x"0000" when x"60E7",
			x"0000" when x"60E8",
			x"0000" when x"60E9",
			x"0000" when x"60EA",
			x"0000" when x"60EB",
			x"0000" when x"60EC",
			x"0000" when x"60ED",
			x"0000" when x"60EE",
			x"0000" when x"60EF",
			x"0000" when x"60F0",
			x"0000" when x"60F1",
			x"0000" when x"60F2",
			x"0000" when x"60F3",
			x"0000" when x"60F4",
			x"0000" when x"60F5",
			x"0000" when x"60F6",
			x"0000" when x"60F7",
			x"0000" when x"60F8",
			x"0000" when x"60F9",
			x"0000" when x"60FA",
			x"0000" when x"60FB",
			x"0000" when x"60FC",
			x"0000" when x"60FD",
			x"0000" when x"60FE",
			x"0000" when x"60FF",
			x"0000" when x"6100",
			x"0000" when x"6101",
			x"0000" when x"6102",
			x"0000" when x"6103",
			x"0000" when x"6104",
			x"0000" when x"6105",
			x"0000" when x"6106",
			x"0000" when x"6107",
			x"0000" when x"6108",
			x"0000" when x"6109",
			x"0000" when x"610A",
			x"0000" when x"610B",
			x"0000" when x"610C",
			x"0000" when x"610D",
			x"0000" when x"610E",
			x"0000" when x"610F",
			x"0000" when x"6110",
			x"0000" when x"6111",
			x"0000" when x"6112",
			x"0000" when x"6113",
			x"0000" when x"6114",
			x"0000" when x"6115",
			x"0000" when x"6116",
			x"0000" when x"6117",
			x"0000" when x"6118",
			x"0000" when x"6119",
			x"0000" when x"611A",
			x"0000" when x"611B",
			x"0000" when x"611C",
			x"0000" when x"611D",
			x"0000" when x"611E",
			x"0000" when x"611F",
			x"0000" when x"6120",
			x"0000" when x"6121",
			x"0000" when x"6122",
			x"0000" when x"6123",
			x"0000" when x"6124",
			x"0000" when x"6125",
			x"0000" when x"6126",
			x"0000" when x"6127",
			x"0000" when x"6128",
			x"0000" when x"6129",
			x"0000" when x"612A",
			x"0000" when x"612B",
			x"0000" when x"612C",
			x"0000" when x"612D",
			x"0000" when x"612E",
			x"0000" when x"612F",
			x"0000" when x"6130",
			x"0000" when x"6131",
			x"0000" when x"6132",
			x"0000" when x"6133",
			x"0000" when x"6134",
			x"0000" when x"6135",
			x"0000" when x"6136",
			x"0000" when x"6137",
			x"0000" when x"6138",
			x"0000" when x"6139",
			x"0000" when x"613A",
			x"0000" when x"613B",
			x"0000" when x"613C",
			x"0000" when x"613D",
			x"0000" when x"613E",
			x"0000" when x"613F",
			x"0000" when x"6140",
			x"0000" when x"6141",
			x"0000" when x"6142",
			x"0000" when x"6143",
			x"0000" when x"6144",
			x"0000" when x"6145",
			x"0000" when x"6146",
			x"0000" when x"6147",
			x"0000" when x"6148",
			x"0000" when x"6149",
			x"0000" when x"614A",
			x"0000" when x"614B",
			x"0000" when x"614C",
			x"0000" when x"614D",
			x"0000" when x"614E",
			x"0000" when x"614F",
			x"0000" when x"6150",
			x"0000" when x"6151",
			x"0000" when x"6152",
			x"0000" when x"6153",
			x"0000" when x"6154",
			x"0000" when x"6155",
			x"0000" when x"6156",
			x"0000" when x"6157",
			x"0000" when x"6158",
			x"0000" when x"6159",
			x"0000" when x"615A",
			x"0000" when x"615B",
			x"0000" when x"615C",
			x"0000" when x"615D",
			x"0000" when x"615E",
			x"0000" when x"615F",
			x"0000" when x"6160",
			x"0000" when x"6161",
			x"0000" when x"6162",
			x"0000" when x"6163",
			x"0000" when x"6164",
			x"0000" when x"6165",
			x"0000" when x"6166",
			x"0000" when x"6167",
			x"0000" when x"6168",
			x"0000" when x"6169",
			x"0000" when x"616A",
			x"0000" when x"616B",
			x"0000" when x"616C",
			x"0000" when x"616D",
			x"0000" when x"616E",
			x"0000" when x"616F",
			x"0000" when x"6170",
			x"0000" when x"6171",
			x"0000" when x"6172",
			x"0000" when x"6173",
			x"0000" when x"6174",
			x"0000" when x"6175",
			x"0000" when x"6176",
			x"0000" when x"6177",
			x"0000" when x"6178",
			x"0000" when x"6179",
			x"0000" when x"617A",
			x"0000" when x"617B",
			x"0000" when x"617C",
			x"0000" when x"617D",
			x"0000" when x"617E",
			x"0000" when x"617F",
			x"0000" when x"6180",
			x"0000" when x"6181",
			x"0000" when x"6182",
			x"0000" when x"6183",
			x"0000" when x"6184",
			x"0000" when x"6185",
			x"0000" when x"6186",
			x"0000" when x"6187",
			x"0000" when x"6188",
			x"0000" when x"6189",
			x"0000" when x"618A",
			x"0000" when x"618B",
			x"0000" when x"618C",
			x"0000" when x"618D",
			x"0000" when x"618E",
			x"0000" when x"618F",
			x"0000" when x"6190",
			x"0000" when x"6191",
			x"0000" when x"6192",
			x"0000" when x"6193",
			x"0000" when x"6194",
			x"0000" when x"6195",
			x"0000" when x"6196",
			x"0000" when x"6197",
			x"0000" when x"6198",
			x"0000" when x"6199",
			x"0000" when x"619A",
			x"0000" when x"619B",
			x"0000" when x"619C",
			x"0000" when x"619D",
			x"0000" when x"619E",
			x"0000" when x"619F",
			x"0000" when x"61A0",
			x"0000" when x"61A1",
			x"0000" when x"61A2",
			x"0000" when x"61A3",
			x"0000" when x"61A4",
			x"0000" when x"61A5",
			x"0000" when x"61A6",
			x"0000" when x"61A7",
			x"0000" when x"61A8",
			x"0000" when x"61A9",
			x"0000" when x"61AA",
			x"0000" when x"61AB",
			x"0000" when x"61AC",
			x"0000" when x"61AD",
			x"0000" when x"61AE",
			x"0000" when x"61AF",
			x"0000" when x"61B0",
			x"0000" when x"61B1",
			x"0000" when x"61B2",
			x"0000" when x"61B3",
			x"0000" when x"61B4",
			x"0000" when x"61B5",
			x"0000" when x"61B6",
			x"0000" when x"61B7",
			x"0000" when x"61B8",
			x"0000" when x"61B9",
			x"0000" when x"61BA",
			x"0000" when x"61BB",
			x"0000" when x"61BC",
			x"0000" when x"61BD",
			x"0000" when x"61BE",
			x"0000" when x"61BF",
			x"0000" when x"61C0",
			x"0000" when x"61C1",
			x"0000" when x"61C2",
			x"0000" when x"61C3",
			x"0000" when x"61C4",
			x"0000" when x"61C5",
			x"0000" when x"61C6",
			x"0000" when x"61C7",
			x"0000" when x"61C8",
			x"0000" when x"61C9",
			x"0000" when x"61CA",
			x"0000" when x"61CB",
			x"0000" when x"61CC",
			x"0000" when x"61CD",
			x"0000" when x"61CE",
			x"0000" when x"61CF",
			x"0000" when x"61D0",
			x"0000" when x"61D1",
			x"0000" when x"61D2",
			x"0000" when x"61D3",
			x"0000" when x"61D4",
			x"0000" when x"61D5",
			x"0000" when x"61D6",
			x"0000" when x"61D7",
			x"0000" when x"61D8",
			x"0000" when x"61D9",
			x"0000" when x"61DA",
			x"0000" when x"61DB",
			x"0000" when x"61DC",
			x"0000" when x"61DD",
			x"0000" when x"61DE",
			x"0000" when x"61DF",
			x"0000" when x"61E0",
			x"0000" when x"61E1",
			x"0000" when x"61E2",
			x"0000" when x"61E3",
			x"0000" when x"61E4",
			x"0000" when x"61E5",
			x"0000" when x"61E6",
			x"0000" when x"61E7",
			x"0000" when x"61E8",
			x"0000" when x"61E9",
			x"0000" when x"61EA",
			x"0000" when x"61EB",
			x"0000" when x"61EC",
			x"0000" when x"61ED",
			x"0000" when x"61EE",
			x"0000" when x"61EF",
			x"0000" when x"61F0",
			x"0000" when x"61F1",
			x"0000" when x"61F2",
			x"0000" when x"61F3",
			x"0000" when x"61F4",
			x"0000" when x"61F5",
			x"0000" when x"61F6",
			x"0000" when x"61F7",
			x"0000" when x"61F8",
			x"0000" when x"61F9",
			x"0000" when x"61FA",
			x"0000" when x"61FB",
			x"0000" when x"61FC",
			x"0000" when x"61FD",
			x"0000" when x"61FE",
			x"0000" when x"61FF",
			x"0000" when x"6200",
			x"0000" when x"6201",
			x"0000" when x"6202",
			x"0000" when x"6203",
			x"0000" when x"6204",
			x"0000" when x"6205",
			x"0000" when x"6206",
			x"0000" when x"6207",
			x"0000" when x"6208",
			x"0000" when x"6209",
			x"0000" when x"620A",
			x"0000" when x"620B",
			x"0000" when x"620C",
			x"0000" when x"620D",
			x"0000" when x"620E",
			x"0000" when x"620F",
			x"0000" when x"6210",
			x"0000" when x"6211",
			x"0000" when x"6212",
			x"0000" when x"6213",
			x"0000" when x"6214",
			x"0000" when x"6215",
			x"0000" when x"6216",
			x"0000" when x"6217",
			x"0000" when x"6218",
			x"0000" when x"6219",
			x"0000" when x"621A",
			x"0000" when x"621B",
			x"0000" when x"621C",
			x"0000" when x"621D",
			x"0000" when x"621E",
			x"0000" when x"621F",
			x"0000" when x"6220",
			x"0000" when x"6221",
			x"0000" when x"6222",
			x"0000" when x"6223",
			x"0000" when x"6224",
			x"0000" when x"6225",
			x"0000" when x"6226",
			x"0000" when x"6227",
			x"0000" when x"6228",
			x"0000" when x"6229",
			x"0000" when x"622A",
			x"0000" when x"622B",
			x"0000" when x"622C",
			x"0000" when x"622D",
			x"0000" when x"622E",
			x"0000" when x"622F",
			x"0000" when x"6230",
			x"0000" when x"6231",
			x"0000" when x"6232",
			x"0000" when x"6233",
			x"0000" when x"6234",
			x"0000" when x"6235",
			x"0000" when x"6236",
			x"0000" when x"6237",
			x"0000" when x"6238",
			x"0000" when x"6239",
			x"0000" when x"623A",
			x"0000" when x"623B",
			x"0000" when x"623C",
			x"0000" when x"623D",
			x"0000" when x"623E",
			x"0000" when x"623F",
			x"0000" when x"6240",
			x"0000" when x"6241",
			x"0000" when x"6242",
			x"0000" when x"6243",
			x"0000" when x"6244",
			x"0000" when x"6245",
			x"0000" when x"6246",
			x"0000" when x"6247",
			x"0000" when x"6248",
			x"0000" when x"6249",
			x"0000" when x"624A",
			x"0000" when x"624B",
			x"0000" when x"624C",
			x"0000" when x"624D",
			x"0000" when x"624E",
			x"0000" when x"624F",
			x"0000" when x"6250",
			x"0000" when x"6251",
			x"0000" when x"6252",
			x"0000" when x"6253",
			x"0000" when x"6254",
			x"0000" when x"6255",
			x"0000" when x"6256",
			x"0000" when x"6257",
			x"0000" when x"6258",
			x"0000" when x"6259",
			x"0000" when x"625A",
			x"0000" when x"625B",
			x"0000" when x"625C",
			x"0000" when x"625D",
			x"0000" when x"625E",
			x"0000" when x"625F",
			x"0000" when x"6260",
			x"0000" when x"6261",
			x"0000" when x"6262",
			x"0000" when x"6263",
			x"0000" when x"6264",
			x"0000" when x"6265",
			x"0000" when x"6266",
			x"0000" when x"6267",
			x"0000" when x"6268",
			x"0000" when x"6269",
			x"0000" when x"626A",
			x"0000" when x"626B",
			x"0000" when x"626C",
			x"0000" when x"626D",
			x"0000" when x"626E",
			x"0000" when x"626F",
			x"0000" when x"6270",
			x"0000" when x"6271",
			x"0000" when x"6272",
			x"0000" when x"6273",
			x"0000" when x"6274",
			x"0000" when x"6275",
			x"0000" when x"6276",
			x"0000" when x"6277",
			x"0000" when x"6278",
			x"0000" when x"6279",
			x"0000" when x"627A",
			x"0000" when x"627B",
			x"0000" when x"627C",
			x"0000" when x"627D",
			x"0000" when x"627E",
			x"0000" when x"627F",
			x"0000" when x"6280",
			x"0000" when x"6281",
			x"0000" when x"6282",
			x"0000" when x"6283",
			x"0000" when x"6284",
			x"0000" when x"6285",
			x"0000" when x"6286",
			x"0000" when x"6287",
			x"0000" when x"6288",
			x"0000" when x"6289",
			x"0000" when x"628A",
			x"0000" when x"628B",
			x"0000" when x"628C",
			x"0000" when x"628D",
			x"0000" when x"628E",
			x"0000" when x"628F",
			x"0000" when x"6290",
			x"0000" when x"6291",
			x"0000" when x"6292",
			x"0000" when x"6293",
			x"0000" when x"6294",
			x"0000" when x"6295",
			x"0000" when x"6296",
			x"0000" when x"6297",
			x"0000" when x"6298",
			x"0000" when x"6299",
			x"0000" when x"629A",
			x"0000" when x"629B",
			x"0000" when x"629C",
			x"0000" when x"629D",
			x"0000" when x"629E",
			x"0000" when x"629F",
			x"0000" when x"62A0",
			x"0000" when x"62A1",
			x"0000" when x"62A2",
			x"0000" when x"62A3",
			x"0000" when x"62A4",
			x"0000" when x"62A5",
			x"0000" when x"62A6",
			x"0000" when x"62A7",
			x"0000" when x"62A8",
			x"0000" when x"62A9",
			x"0000" when x"62AA",
			x"0000" when x"62AB",
			x"0000" when x"62AC",
			x"0000" when x"62AD",
			x"0000" when x"62AE",
			x"0000" when x"62AF",
			x"0000" when x"62B0",
			x"0000" when x"62B1",
			x"0000" when x"62B2",
			x"0000" when x"62B3",
			x"0000" when x"62B4",
			x"0000" when x"62B5",
			x"0000" when x"62B6",
			x"0000" when x"62B7",
			x"0000" when x"62B8",
			x"0000" when x"62B9",
			x"0000" when x"62BA",
			x"0000" when x"62BB",
			x"0000" when x"62BC",
			x"0000" when x"62BD",
			x"0000" when x"62BE",
			x"0000" when x"62BF",
			x"0000" when x"62C0",
			x"0000" when x"62C1",
			x"0000" when x"62C2",
			x"0000" when x"62C3",
			x"0000" when x"62C4",
			x"0000" when x"62C5",
			x"0000" when x"62C6",
			x"0000" when x"62C7",
			x"0000" when x"62C8",
			x"0000" when x"62C9",
			x"0000" when x"62CA",
			x"0000" when x"62CB",
			x"0000" when x"62CC",
			x"0000" when x"62CD",
			x"0000" when x"62CE",
			x"0000" when x"62CF",
			x"0000" when x"62D0",
			x"0000" when x"62D1",
			x"0000" when x"62D2",
			x"0000" when x"62D3",
			x"0000" when x"62D4",
			x"0000" when x"62D5",
			x"0000" when x"62D6",
			x"0000" when x"62D7",
			x"0000" when x"62D8",
			x"0000" when x"62D9",
			x"0000" when x"62DA",
			x"0000" when x"62DB",
			x"0000" when x"62DC",
			x"0000" when x"62DD",
			x"0000" when x"62DE",
			x"0000" when x"62DF",
			x"0000" when x"62E0",
			x"0000" when x"62E1",
			x"0000" when x"62E2",
			x"0000" when x"62E3",
			x"0000" when x"62E4",
			x"0000" when x"62E5",
			x"0000" when x"62E6",
			x"0000" when x"62E7",
			x"0000" when x"62E8",
			x"0000" when x"62E9",
			x"0000" when x"62EA",
			x"0000" when x"62EB",
			x"0000" when x"62EC",
			x"0000" when x"62ED",
			x"0000" when x"62EE",
			x"0000" when x"62EF",
			x"0000" when x"62F0",
			x"0000" when x"62F1",
			x"0000" when x"62F2",
			x"0000" when x"62F3",
			x"0000" when x"62F4",
			x"0000" when x"62F5",
			x"0000" when x"62F6",
			x"0000" when x"62F7",
			x"0000" when x"62F8",
			x"0000" when x"62F9",
			x"0000" when x"62FA",
			x"0000" when x"62FB",
			x"0000" when x"62FC",
			x"0000" when x"62FD",
			x"0000" when x"62FE",
			x"0000" when x"62FF",
			x"0000" when x"6300",
			x"0000" when x"6301",
			x"0000" when x"6302",
			x"0000" when x"6303",
			x"0000" when x"6304",
			x"0000" when x"6305",
			x"0000" when x"6306",
			x"0000" when x"6307",
			x"0000" when x"6308",
			x"0000" when x"6309",
			x"0000" when x"630A",
			x"0000" when x"630B",
			x"0000" when x"630C",
			x"0000" when x"630D",
			x"0000" when x"630E",
			x"0000" when x"630F",
			x"0000" when x"6310",
			x"0000" when x"6311",
			x"0000" when x"6312",
			x"0000" when x"6313",
			x"0000" when x"6314",
			x"0000" when x"6315",
			x"0000" when x"6316",
			x"0000" when x"6317",
			x"0000" when x"6318",
			x"0000" when x"6319",
			x"0000" when x"631A",
			x"0000" when x"631B",
			x"0000" when x"631C",
			x"0000" when x"631D",
			x"0000" when x"631E",
			x"0000" when x"631F",
			x"0000" when x"6320",
			x"0000" when x"6321",
			x"0000" when x"6322",
			x"0000" when x"6323",
			x"0000" when x"6324",
			x"0000" when x"6325",
			x"0000" when x"6326",
			x"0000" when x"6327",
			x"0000" when x"6328",
			x"0000" when x"6329",
			x"0000" when x"632A",
			x"0000" when x"632B",
			x"0000" when x"632C",
			x"0000" when x"632D",
			x"0000" when x"632E",
			x"0000" when x"632F",
			x"0000" when x"6330",
			x"0000" when x"6331",
			x"0000" when x"6332",
			x"0000" when x"6333",
			x"0000" when x"6334",
			x"0000" when x"6335",
			x"0000" when x"6336",
			x"0000" when x"6337",
			x"0000" when x"6338",
			x"0000" when x"6339",
			x"0000" when x"633A",
			x"0000" when x"633B",
			x"0000" when x"633C",
			x"0000" when x"633D",
			x"0000" when x"633E",
			x"0000" when x"633F",
			x"0000" when x"6340",
			x"0000" when x"6341",
			x"0000" when x"6342",
			x"0000" when x"6343",
			x"0000" when x"6344",
			x"0000" when x"6345",
			x"0000" when x"6346",
			x"0000" when x"6347",
			x"0000" when x"6348",
			x"0000" when x"6349",
			x"0000" when x"634A",
			x"0000" when x"634B",
			x"0000" when x"634C",
			x"0000" when x"634D",
			x"0000" when x"634E",
			x"0000" when x"634F",
			x"0000" when x"6350",
			x"0000" when x"6351",
			x"0000" when x"6352",
			x"0000" when x"6353",
			x"0000" when x"6354",
			x"0000" when x"6355",
			x"0000" when x"6356",
			x"0000" when x"6357",
			x"0000" when x"6358",
			x"0000" when x"6359",
			x"0000" when x"635A",
			x"0000" when x"635B",
			x"0000" when x"635C",
			x"0000" when x"635D",
			x"0000" when x"635E",
			x"0000" when x"635F",
			x"0000" when x"6360",
			x"0000" when x"6361",
			x"0000" when x"6362",
			x"0000" when x"6363",
			x"0000" when x"6364",
			x"0000" when x"6365",
			x"0000" when x"6366",
			x"0000" when x"6367",
			x"0000" when x"6368",
			x"0000" when x"6369",
			x"0000" when x"636A",
			x"0000" when x"636B",
			x"0000" when x"636C",
			x"0000" when x"636D",
			x"0000" when x"636E",
			x"0000" when x"636F",
			x"0000" when x"6370",
			x"0000" when x"6371",
			x"0000" when x"6372",
			x"0000" when x"6373",
			x"0000" when x"6374",
			x"0000" when x"6375",
			x"0000" when x"6376",
			x"0000" when x"6377",
			x"0000" when x"6378",
			x"0000" when x"6379",
			x"0000" when x"637A",
			x"0000" when x"637B",
			x"0000" when x"637C",
			x"0000" when x"637D",
			x"0000" when x"637E",
			x"0000" when x"637F",
			x"0000" when x"6380",
			x"0000" when x"6381",
			x"0000" when x"6382",
			x"0000" when x"6383",
			x"0000" when x"6384",
			x"0000" when x"6385",
			x"0000" when x"6386",
			x"0000" when x"6387",
			x"0000" when x"6388",
			x"0000" when x"6389",
			x"0000" when x"638A",
			x"0000" when x"638B",
			x"0000" when x"638C",
			x"0000" when x"638D",
			x"0000" when x"638E",
			x"0000" when x"638F",
			x"0000" when x"6390",
			x"0000" when x"6391",
			x"0000" when x"6392",
			x"0000" when x"6393",
			x"0000" when x"6394",
			x"0000" when x"6395",
			x"0000" when x"6396",
			x"0000" when x"6397",
			x"0000" when x"6398",
			x"0000" when x"6399",
			x"0000" when x"639A",
			x"0000" when x"639B",
			x"0000" when x"639C",
			x"0000" when x"639D",
			x"0000" when x"639E",
			x"0000" when x"639F",
			x"0000" when x"63A0",
			x"0000" when x"63A1",
			x"0000" when x"63A2",
			x"0000" when x"63A3",
			x"0000" when x"63A4",
			x"0000" when x"63A5",
			x"0000" when x"63A6",
			x"0000" when x"63A7",
			x"0000" when x"63A8",
			x"0000" when x"63A9",
			x"0000" when x"63AA",
			x"0000" when x"63AB",
			x"0000" when x"63AC",
			x"0000" when x"63AD",
			x"0000" when x"63AE",
			x"0000" when x"63AF",
			x"0000" when x"63B0",
			x"0000" when x"63B1",
			x"0000" when x"63B2",
			x"0000" when x"63B3",
			x"0000" when x"63B4",
			x"0000" when x"63B5",
			x"0000" when x"63B6",
			x"0000" when x"63B7",
			x"0000" when x"63B8",
			x"0000" when x"63B9",
			x"0000" when x"63BA",
			x"0000" when x"63BB",
			x"0000" when x"63BC",
			x"0000" when x"63BD",
			x"0000" when x"63BE",
			x"0000" when x"63BF",
			x"0000" when x"63C0",
			x"0000" when x"63C1",
			x"0000" when x"63C2",
			x"0000" when x"63C3",
			x"0000" when x"63C4",
			x"0000" when x"63C5",
			x"0000" when x"63C6",
			x"0000" when x"63C7",
			x"0000" when x"63C8",
			x"0000" when x"63C9",
			x"0000" when x"63CA",
			x"0000" when x"63CB",
			x"0000" when x"63CC",
			x"0000" when x"63CD",
			x"0000" when x"63CE",
			x"0000" when x"63CF",
			x"0000" when x"63D0",
			x"0000" when x"63D1",
			x"0000" when x"63D2",
			x"0000" when x"63D3",
			x"0000" when x"63D4",
			x"0000" when x"63D5",
			x"0000" when x"63D6",
			x"0000" when x"63D7",
			x"0000" when x"63D8",
			x"0000" when x"63D9",
			x"0000" when x"63DA",
			x"0000" when x"63DB",
			x"0000" when x"63DC",
			x"0000" when x"63DD",
			x"0000" when x"63DE",
			x"0000" when x"63DF",
			x"0000" when x"63E0",
			x"0000" when x"63E1",
			x"0000" when x"63E2",
			x"0000" when x"63E3",
			x"0000" when x"63E4",
			x"0000" when x"63E5",
			x"0000" when x"63E6",
			x"0000" when x"63E7",
			x"0000" when x"63E8",
			x"0000" when x"63E9",
			x"0000" when x"63EA",
			x"0000" when x"63EB",
			x"0000" when x"63EC",
			x"0000" when x"63ED",
			x"0000" when x"63EE",
			x"0000" when x"63EF",
			x"0000" when x"63F0",
			x"0000" when x"63F1",
			x"0000" when x"63F2",
			x"0000" when x"63F3",
			x"0000" when x"63F4",
			x"0000" when x"63F5",
			x"0000" when x"63F6",
			x"0000" when x"63F7",
			x"0000" when x"63F8",
			x"0000" when x"63F9",
			x"0000" when x"63FA",
			x"0000" when x"63FB",
			x"0000" when x"63FC",
			x"0000" when x"63FD",
			x"0000" when x"63FE",
			x"0000" when x"63FF",
			x"0000" when x"6400",
			x"0000" when x"6401",
			x"0000" when x"6402",
			x"0000" when x"6403",
			x"0000" when x"6404",
			x"0000" when x"6405",
			x"0000" when x"6406",
			x"0000" when x"6407",
			x"0000" when x"6408",
			x"0000" when x"6409",
			x"0000" when x"640A",
			x"0000" when x"640B",
			x"0000" when x"640C",
			x"0000" when x"640D",
			x"0000" when x"640E",
			x"0000" when x"640F",
			x"0000" when x"6410",
			x"0000" when x"6411",
			x"0000" when x"6412",
			x"0000" when x"6413",
			x"0000" when x"6414",
			x"0000" when x"6415",
			x"0000" when x"6416",
			x"0000" when x"6417",
			x"0000" when x"6418",
			x"0000" when x"6419",
			x"0000" when x"641A",
			x"0000" when x"641B",
			x"0000" when x"641C",
			x"0000" when x"641D",
			x"0000" when x"641E",
			x"0000" when x"641F",
			x"0000" when x"6420",
			x"0000" when x"6421",
			x"0000" when x"6422",
			x"0000" when x"6423",
			x"0000" when x"6424",
			x"0000" when x"6425",
			x"0000" when x"6426",
			x"0000" when x"6427",
			x"0000" when x"6428",
			x"0000" when x"6429",
			x"0000" when x"642A",
			x"0000" when x"642B",
			x"0000" when x"642C",
			x"0000" when x"642D",
			x"0000" when x"642E",
			x"0000" when x"642F",
			x"0000" when x"6430",
			x"0000" when x"6431",
			x"0000" when x"6432",
			x"0000" when x"6433",
			x"0000" when x"6434",
			x"0000" when x"6435",
			x"0000" when x"6436",
			x"0000" when x"6437",
			x"0000" when x"6438",
			x"0000" when x"6439",
			x"0000" when x"643A",
			x"0000" when x"643B",
			x"0000" when x"643C",
			x"0000" when x"643D",
			x"0000" when x"643E",
			x"0000" when x"643F",
			x"0000" when x"6440",
			x"0000" when x"6441",
			x"0000" when x"6442",
			x"0000" when x"6443",
			x"0000" when x"6444",
			x"0000" when x"6445",
			x"0000" when x"6446",
			x"0000" when x"6447",
			x"0000" when x"6448",
			x"0000" when x"6449",
			x"0000" when x"644A",
			x"0000" when x"644B",
			x"0000" when x"644C",
			x"0000" when x"644D",
			x"0000" when x"644E",
			x"0000" when x"644F",
			x"0000" when x"6450",
			x"0000" when x"6451",
			x"0000" when x"6452",
			x"0000" when x"6453",
			x"0000" when x"6454",
			x"0000" when x"6455",
			x"0000" when x"6456",
			x"0000" when x"6457",
			x"0000" when x"6458",
			x"0000" when x"6459",
			x"0000" when x"645A",
			x"0000" when x"645B",
			x"0000" when x"645C",
			x"0000" when x"645D",
			x"0000" when x"645E",
			x"0000" when x"645F",
			x"0000" when x"6460",
			x"0000" when x"6461",
			x"0000" when x"6462",
			x"0000" when x"6463",
			x"0000" when x"6464",
			x"0000" when x"6465",
			x"0000" when x"6466",
			x"0000" when x"6467",
			x"0000" when x"6468",
			x"0000" when x"6469",
			x"0000" when x"646A",
			x"0000" when x"646B",
			x"0000" when x"646C",
			x"0000" when x"646D",
			x"0000" when x"646E",
			x"0000" when x"646F",
			x"0000" when x"6470",
			x"0000" when x"6471",
			x"0000" when x"6472",
			x"0000" when x"6473",
			x"0000" when x"6474",
			x"0000" when x"6475",
			x"0000" when x"6476",
			x"0000" when x"6477",
			x"0000" when x"6478",
			x"0000" when x"6479",
			x"0000" when x"647A",
			x"0000" when x"647B",
			x"0000" when x"647C",
			x"0000" when x"647D",
			x"0000" when x"647E",
			x"0000" when x"647F",
			x"0000" when x"6480",
			x"0000" when x"6481",
			x"0000" when x"6482",
			x"0000" when x"6483",
			x"0000" when x"6484",
			x"0000" when x"6485",
			x"0000" when x"6486",
			x"0000" when x"6487",
			x"0000" when x"6488",
			x"0000" when x"6489",
			x"0000" when x"648A",
			x"0000" when x"648B",
			x"0000" when x"648C",
			x"0000" when x"648D",
			x"0000" when x"648E",
			x"0000" when x"648F",
			x"0000" when x"6490",
			x"0000" when x"6491",
			x"0000" when x"6492",
			x"0000" when x"6493",
			x"0000" when x"6494",
			x"0000" when x"6495",
			x"0000" when x"6496",
			x"0000" when x"6497",
			x"0000" when x"6498",
			x"0000" when x"6499",
			x"0000" when x"649A",
			x"0000" when x"649B",
			x"0000" when x"649C",
			x"0000" when x"649D",
			x"0000" when x"649E",
			x"0000" when x"649F",
			x"0000" when x"64A0",
			x"0000" when x"64A1",
			x"0000" when x"64A2",
			x"0000" when x"64A3",
			x"0000" when x"64A4",
			x"0000" when x"64A5",
			x"0000" when x"64A6",
			x"0000" when x"64A7",
			x"0000" when x"64A8",
			x"0000" when x"64A9",
			x"0000" when x"64AA",
			x"0000" when x"64AB",
			x"0000" when x"64AC",
			x"0000" when x"64AD",
			x"0000" when x"64AE",
			x"0000" when x"64AF",
			x"0000" when x"64B0",
			x"0000" when x"64B1",
			x"0000" when x"64B2",
			x"0000" when x"64B3",
			x"0000" when x"64B4",
			x"0000" when x"64B5",
			x"0000" when x"64B6",
			x"0000" when x"64B7",
			x"0000" when x"64B8",
			x"0000" when x"64B9",
			x"0000" when x"64BA",
			x"0000" when x"64BB",
			x"0000" when x"64BC",
			x"0000" when x"64BD",
			x"0000" when x"64BE",
			x"0000" when x"64BF",
			x"0000" when x"64C0",
			x"0000" when x"64C1",
			x"0000" when x"64C2",
			x"0000" when x"64C3",
			x"0000" when x"64C4",
			x"0000" when x"64C5",
			x"0000" when x"64C6",
			x"0000" when x"64C7",
			x"0000" when x"64C8",
			x"0000" when x"64C9",
			x"0000" when x"64CA",
			x"0000" when x"64CB",
			x"0000" when x"64CC",
			x"0000" when x"64CD",
			x"0000" when x"64CE",
			x"0000" when x"64CF",
			x"0000" when x"64D0",
			x"0000" when x"64D1",
			x"0000" when x"64D2",
			x"0000" when x"64D3",
			x"0000" when x"64D4",
			x"0000" when x"64D5",
			x"0000" when x"64D6",
			x"0000" when x"64D7",
			x"0000" when x"64D8",
			x"0000" when x"64D9",
			x"0000" when x"64DA",
			x"0000" when x"64DB",
			x"0000" when x"64DC",
			x"0000" when x"64DD",
			x"0000" when x"64DE",
			x"0000" when x"64DF",
			x"0000" when x"64E0",
			x"0000" when x"64E1",
			x"0000" when x"64E2",
			x"0000" when x"64E3",
			x"0000" when x"64E4",
			x"0000" when x"64E5",
			x"0000" when x"64E6",
			x"0000" when x"64E7",
			x"0000" when x"64E8",
			x"0000" when x"64E9",
			x"0000" when x"64EA",
			x"0000" when x"64EB",
			x"0000" when x"64EC",
			x"0000" when x"64ED",
			x"0000" when x"64EE",
			x"0000" when x"64EF",
			x"0000" when x"64F0",
			x"0000" when x"64F1",
			x"0000" when x"64F2",
			x"0000" when x"64F3",
			x"0000" when x"64F4",
			x"0000" when x"64F5",
			x"0000" when x"64F6",
			x"0000" when x"64F7",
			x"0000" when x"64F8",
			x"0000" when x"64F9",
			x"0000" when x"64FA",
			x"0000" when x"64FB",
			x"0000" when x"64FC",
			x"0000" when x"64FD",
			x"0000" when x"64FE",
			x"0000" when x"64FF",
			x"0000" when x"6500",
			x"0000" when x"6501",
			x"0000" when x"6502",
			x"0000" when x"6503",
			x"0000" when x"6504",
			x"0000" when x"6505",
			x"0000" when x"6506",
			x"0000" when x"6507",
			x"0000" when x"6508",
			x"0000" when x"6509",
			x"0000" when x"650A",
			x"0000" when x"650B",
			x"0000" when x"650C",
			x"0000" when x"650D",
			x"0000" when x"650E",
			x"0000" when x"650F",
			x"0000" when x"6510",
			x"0000" when x"6511",
			x"0000" when x"6512",
			x"0000" when x"6513",
			x"0000" when x"6514",
			x"0000" when x"6515",
			x"0000" when x"6516",
			x"0000" when x"6517",
			x"0000" when x"6518",
			x"0000" when x"6519",
			x"0000" when x"651A",
			x"0000" when x"651B",
			x"0000" when x"651C",
			x"0000" when x"651D",
			x"0000" when x"651E",
			x"0000" when x"651F",
			x"0000" when x"6520",
			x"0000" when x"6521",
			x"0000" when x"6522",
			x"0000" when x"6523",
			x"0000" when x"6524",
			x"0000" when x"6525",
			x"0000" when x"6526",
			x"0000" when x"6527",
			x"0000" when x"6528",
			x"0000" when x"6529",
			x"0000" when x"652A",
			x"0000" when x"652B",
			x"0000" when x"652C",
			x"0000" when x"652D",
			x"0000" when x"652E",
			x"0000" when x"652F",
			x"0000" when x"6530",
			x"0000" when x"6531",
			x"0000" when x"6532",
			x"0000" when x"6533",
			x"0000" when x"6534",
			x"0000" when x"6535",
			x"0000" when x"6536",
			x"0000" when x"6537",
			x"0000" when x"6538",
			x"0000" when x"6539",
			x"0000" when x"653A",
			x"0000" when x"653B",
			x"0000" when x"653C",
			x"0000" when x"653D",
			x"0000" when x"653E",
			x"0000" when x"653F",
			x"0000" when x"6540",
			x"0000" when x"6541",
			x"0000" when x"6542",
			x"0000" when x"6543",
			x"0000" when x"6544",
			x"0000" when x"6545",
			x"0000" when x"6546",
			x"0000" when x"6547",
			x"0000" when x"6548",
			x"0000" when x"6549",
			x"0000" when x"654A",
			x"0000" when x"654B",
			x"0000" when x"654C",
			x"0000" when x"654D",
			x"0000" when x"654E",
			x"0000" when x"654F",
			x"0000" when x"6550",
			x"0000" when x"6551",
			x"0000" when x"6552",
			x"0000" when x"6553",
			x"0000" when x"6554",
			x"0000" when x"6555",
			x"0000" when x"6556",
			x"0000" when x"6557",
			x"0000" when x"6558",
			x"0000" when x"6559",
			x"0000" when x"655A",
			x"0000" when x"655B",
			x"0000" when x"655C",
			x"0000" when x"655D",
			x"0000" when x"655E",
			x"0000" when x"655F",
			x"0000" when x"6560",
			x"0000" when x"6561",
			x"0000" when x"6562",
			x"0000" when x"6563",
			x"0000" when x"6564",
			x"0000" when x"6565",
			x"0000" when x"6566",
			x"0000" when x"6567",
			x"0000" when x"6568",
			x"0000" when x"6569",
			x"0000" when x"656A",
			x"0000" when x"656B",
			x"0000" when x"656C",
			x"0000" when x"656D",
			x"0000" when x"656E",
			x"0000" when x"656F",
			x"0000" when x"6570",
			x"0000" when x"6571",
			x"0000" when x"6572",
			x"0000" when x"6573",
			x"0000" when x"6574",
			x"0000" when x"6575",
			x"0000" when x"6576",
			x"0000" when x"6577",
			x"0000" when x"6578",
			x"0000" when x"6579",
			x"0000" when x"657A",
			x"0000" when x"657B",
			x"0000" when x"657C",
			x"0000" when x"657D",
			x"0000" when x"657E",
			x"0000" when x"657F",
			x"0000" when x"6580",
			x"0000" when x"6581",
			x"0000" when x"6582",
			x"0000" when x"6583",
			x"0000" when x"6584",
			x"0000" when x"6585",
			x"0000" when x"6586",
			x"0000" when x"6587",
			x"0000" when x"6588",
			x"0000" when x"6589",
			x"0000" when x"658A",
			x"0000" when x"658B",
			x"0000" when x"658C",
			x"0000" when x"658D",
			x"0000" when x"658E",
			x"0000" when x"658F",
			x"0000" when x"6590",
			x"0000" when x"6591",
			x"0000" when x"6592",
			x"0000" when x"6593",
			x"0000" when x"6594",
			x"0000" when x"6595",
			x"0000" when x"6596",
			x"0000" when x"6597",
			x"0000" when x"6598",
			x"0000" when x"6599",
			x"0000" when x"659A",
			x"0000" when x"659B",
			x"0000" when x"659C",
			x"0000" when x"659D",
			x"0000" when x"659E",
			x"0000" when x"659F",
			x"0000" when x"65A0",
			x"0000" when x"65A1",
			x"0000" when x"65A2",
			x"0000" when x"65A3",
			x"0000" when x"65A4",
			x"0000" when x"65A5",
			x"0000" when x"65A6",
			x"0000" when x"65A7",
			x"0000" when x"65A8",
			x"0000" when x"65A9",
			x"0000" when x"65AA",
			x"0000" when x"65AB",
			x"0000" when x"65AC",
			x"0000" when x"65AD",
			x"0000" when x"65AE",
			x"0000" when x"65AF",
			x"0000" when x"65B0",
			x"0000" when x"65B1",
			x"0000" when x"65B2",
			x"0000" when x"65B3",
			x"0000" when x"65B4",
			x"0000" when x"65B5",
			x"0000" when x"65B6",
			x"0000" when x"65B7",
			x"0000" when x"65B8",
			x"0000" when x"65B9",
			x"0000" when x"65BA",
			x"0000" when x"65BB",
			x"0000" when x"65BC",
			x"0000" when x"65BD",
			x"0000" when x"65BE",
			x"0000" when x"65BF",
			x"0000" when x"65C0",
			x"0000" when x"65C1",
			x"0000" when x"65C2",
			x"0000" when x"65C3",
			x"0000" when x"65C4",
			x"0000" when x"65C5",
			x"0000" when x"65C6",
			x"0000" when x"65C7",
			x"0000" when x"65C8",
			x"0000" when x"65C9",
			x"0000" when x"65CA",
			x"0000" when x"65CB",
			x"0000" when x"65CC",
			x"0000" when x"65CD",
			x"0000" when x"65CE",
			x"0000" when x"65CF",
			x"0000" when x"65D0",
			x"0000" when x"65D1",
			x"0000" when x"65D2",
			x"0000" when x"65D3",
			x"0000" when x"65D4",
			x"0000" when x"65D5",
			x"0000" when x"65D6",
			x"0000" when x"65D7",
			x"0000" when x"65D8",
			x"0000" when x"65D9",
			x"0000" when x"65DA",
			x"0000" when x"65DB",
			x"0000" when x"65DC",
			x"0000" when x"65DD",
			x"0000" when x"65DE",
			x"0000" when x"65DF",
			x"0000" when x"65E0",
			x"0000" when x"65E1",
			x"0000" when x"65E2",
			x"0000" when x"65E3",
			x"0000" when x"65E4",
			x"0000" when x"65E5",
			x"0000" when x"65E6",
			x"0000" when x"65E7",
			x"0000" when x"65E8",
			x"0000" when x"65E9",
			x"0000" when x"65EA",
			x"0000" when x"65EB",
			x"0000" when x"65EC",
			x"0000" when x"65ED",
			x"0000" when x"65EE",
			x"0000" when x"65EF",
			x"0000" when x"65F0",
			x"0000" when x"65F1",
			x"0000" when x"65F2",
			x"0000" when x"65F3",
			x"0000" when x"65F4",
			x"0000" when x"65F5",
			x"0000" when x"65F6",
			x"0000" when x"65F7",
			x"0000" when x"65F8",
			x"0000" when x"65F9",
			x"0000" when x"65FA",
			x"0000" when x"65FB",
			x"0000" when x"65FC",
			x"0000" when x"65FD",
			x"0000" when x"65FE",
			x"0000" when x"65FF",
			x"0000" when x"6600",
			x"0000" when x"6601",
			x"0000" when x"6602",
			x"0000" when x"6603",
			x"0000" when x"6604",
			x"0000" when x"6605",
			x"0000" when x"6606",
			x"0000" when x"6607",
			x"0000" when x"6608",
			x"0000" when x"6609",
			x"0000" when x"660A",
			x"0000" when x"660B",
			x"0000" when x"660C",
			x"0000" when x"660D",
			x"0000" when x"660E",
			x"0000" when x"660F",
			x"0000" when x"6610",
			x"0000" when x"6611",
			x"0000" when x"6612",
			x"0000" when x"6613",
			x"0000" when x"6614",
			x"0000" when x"6615",
			x"0000" when x"6616",
			x"0000" when x"6617",
			x"0000" when x"6618",
			x"0000" when x"6619",
			x"0000" when x"661A",
			x"0000" when x"661B",
			x"0000" when x"661C",
			x"0000" when x"661D",
			x"0000" when x"661E",
			x"0000" when x"661F",
			x"0000" when x"6620",
			x"0000" when x"6621",
			x"0000" when x"6622",
			x"0000" when x"6623",
			x"0000" when x"6624",
			x"0000" when x"6625",
			x"0000" when x"6626",
			x"0000" when x"6627",
			x"0000" when x"6628",
			x"0000" when x"6629",
			x"0000" when x"662A",
			x"0000" when x"662B",
			x"0000" when x"662C",
			x"0000" when x"662D",
			x"0000" when x"662E",
			x"0000" when x"662F",
			x"0000" when x"6630",
			x"0000" when x"6631",
			x"0000" when x"6632",
			x"0000" when x"6633",
			x"0000" when x"6634",
			x"0000" when x"6635",
			x"0000" when x"6636",
			x"0000" when x"6637",
			x"0000" when x"6638",
			x"0000" when x"6639",
			x"0000" when x"663A",
			x"0000" when x"663B",
			x"0000" when x"663C",
			x"0000" when x"663D",
			x"0000" when x"663E",
			x"0000" when x"663F",
			x"0000" when x"6640",
			x"0000" when x"6641",
			x"0000" when x"6642",
			x"0000" when x"6643",
			x"0000" when x"6644",
			x"0000" when x"6645",
			x"0000" when x"6646",
			x"0000" when x"6647",
			x"0000" when x"6648",
			x"0000" when x"6649",
			x"0000" when x"664A",
			x"0000" when x"664B",
			x"0000" when x"664C",
			x"0000" when x"664D",
			x"0000" when x"664E",
			x"0000" when x"664F",
			x"0000" when x"6650",
			x"0000" when x"6651",
			x"0000" when x"6652",
			x"0000" when x"6653",
			x"0000" when x"6654",
			x"0000" when x"6655",
			x"0000" when x"6656",
			x"0000" when x"6657",
			x"0000" when x"6658",
			x"0000" when x"6659",
			x"0000" when x"665A",
			x"0000" when x"665B",
			x"0000" when x"665C",
			x"0000" when x"665D",
			x"0000" when x"665E",
			x"0000" when x"665F",
			x"0000" when x"6660",
			x"0000" when x"6661",
			x"0000" when x"6662",
			x"0000" when x"6663",
			x"0000" when x"6664",
			x"0000" when x"6665",
			x"0000" when x"6666",
			x"0000" when x"6667",
			x"0000" when x"6668",
			x"0000" when x"6669",
			x"0000" when x"666A",
			x"0000" when x"666B",
			x"0000" when x"666C",
			x"0000" when x"666D",
			x"0000" when x"666E",
			x"0000" when x"666F",
			x"0000" when x"6670",
			x"0000" when x"6671",
			x"0000" when x"6672",
			x"0000" when x"6673",
			x"0000" when x"6674",
			x"0000" when x"6675",
			x"0000" when x"6676",
			x"0000" when x"6677",
			x"0000" when x"6678",
			x"0000" when x"6679",
			x"0000" when x"667A",
			x"0000" when x"667B",
			x"0000" when x"667C",
			x"0000" when x"667D",
			x"0000" when x"667E",
			x"0000" when x"667F",
			x"0000" when x"6680",
			x"0000" when x"6681",
			x"0000" when x"6682",
			x"0000" when x"6683",
			x"0000" when x"6684",
			x"0000" when x"6685",
			x"0000" when x"6686",
			x"0000" when x"6687",
			x"0000" when x"6688",
			x"0000" when x"6689",
			x"0000" when x"668A",
			x"0000" when x"668B",
			x"0000" when x"668C",
			x"0000" when x"668D",
			x"0000" when x"668E",
			x"0000" when x"668F",
			x"0000" when x"6690",
			x"0000" when x"6691",
			x"0000" when x"6692",
			x"0000" when x"6693",
			x"0000" when x"6694",
			x"0000" when x"6695",
			x"0000" when x"6696",
			x"0000" when x"6697",
			x"0000" when x"6698",
			x"0000" when x"6699",
			x"0000" when x"669A",
			x"0000" when x"669B",
			x"0000" when x"669C",
			x"0000" when x"669D",
			x"0000" when x"669E",
			x"0000" when x"669F",
			x"0000" when x"66A0",
			x"0000" when x"66A1",
			x"0000" when x"66A2",
			x"0000" when x"66A3",
			x"0000" when x"66A4",
			x"0000" when x"66A5",
			x"0000" when x"66A6",
			x"0000" when x"66A7",
			x"0000" when x"66A8",
			x"0000" when x"66A9",
			x"0000" when x"66AA",
			x"0000" when x"66AB",
			x"0000" when x"66AC",
			x"0000" when x"66AD",
			x"0000" when x"66AE",
			x"0000" when x"66AF",
			x"0000" when x"66B0",
			x"0000" when x"66B1",
			x"0000" when x"66B2",
			x"0000" when x"66B3",
			x"0000" when x"66B4",
			x"0000" when x"66B5",
			x"0000" when x"66B6",
			x"0000" when x"66B7",
			x"0000" when x"66B8",
			x"0000" when x"66B9",
			x"0000" when x"66BA",
			x"0000" when x"66BB",
			x"0000" when x"66BC",
			x"0000" when x"66BD",
			x"0000" when x"66BE",
			x"0000" when x"66BF",
			x"0000" when x"66C0",
			x"0000" when x"66C1",
			x"0000" when x"66C2",
			x"0000" when x"66C3",
			x"0000" when x"66C4",
			x"0000" when x"66C5",
			x"0000" when x"66C6",
			x"0000" when x"66C7",
			x"0000" when x"66C8",
			x"0000" when x"66C9",
			x"0000" when x"66CA",
			x"0000" when x"66CB",
			x"0000" when x"66CC",
			x"0000" when x"66CD",
			x"0000" when x"66CE",
			x"0000" when x"66CF",
			x"0000" when x"66D0",
			x"0000" when x"66D1",
			x"0000" when x"66D2",
			x"0000" when x"66D3",
			x"0000" when x"66D4",
			x"0000" when x"66D5",
			x"0000" when x"66D6",
			x"0000" when x"66D7",
			x"0000" when x"66D8",
			x"0000" when x"66D9",
			x"0000" when x"66DA",
			x"0000" when x"66DB",
			x"0000" when x"66DC",
			x"0000" when x"66DD",
			x"0000" when x"66DE",
			x"0000" when x"66DF",
			x"0000" when x"66E0",
			x"0000" when x"66E1",
			x"0000" when x"66E2",
			x"0000" when x"66E3",
			x"0000" when x"66E4",
			x"0000" when x"66E5",
			x"0000" when x"66E6",
			x"0000" when x"66E7",
			x"0000" when x"66E8",
			x"0000" when x"66E9",
			x"0000" when x"66EA",
			x"0000" when x"66EB",
			x"0000" when x"66EC",
			x"0000" when x"66ED",
			x"0000" when x"66EE",
			x"0000" when x"66EF",
			x"0000" when x"66F0",
			x"0000" when x"66F1",
			x"0000" when x"66F2",
			x"0000" when x"66F3",
			x"0000" when x"66F4",
			x"0000" when x"66F5",
			x"0000" when x"66F6",
			x"0000" when x"66F7",
			x"0000" when x"66F8",
			x"0000" when x"66F9",
			x"0000" when x"66FA",
			x"0000" when x"66FB",
			x"0000" when x"66FC",
			x"0000" when x"66FD",
			x"0000" when x"66FE",
			x"0000" when x"66FF",
			x"0000" when x"6700",
			x"0000" when x"6701",
			x"0000" when x"6702",
			x"0000" when x"6703",
			x"0000" when x"6704",
			x"0000" when x"6705",
			x"0000" when x"6706",
			x"0000" when x"6707",
			x"0000" when x"6708",
			x"0000" when x"6709",
			x"0000" when x"670A",
			x"0000" when x"670B",
			x"0000" when x"670C",
			x"0000" when x"670D",
			x"0000" when x"670E",
			x"0000" when x"670F",
			x"0000" when x"6710",
			x"0000" when x"6711",
			x"0000" when x"6712",
			x"0000" when x"6713",
			x"0000" when x"6714",
			x"0000" when x"6715",
			x"0000" when x"6716",
			x"0000" when x"6717",
			x"0000" when x"6718",
			x"0000" when x"6719",
			x"0000" when x"671A",
			x"0000" when x"671B",
			x"0000" when x"671C",
			x"0000" when x"671D",
			x"0000" when x"671E",
			x"0000" when x"671F",
			x"0000" when x"6720",
			x"0000" when x"6721",
			x"0000" when x"6722",
			x"0000" when x"6723",
			x"0000" when x"6724",
			x"0000" when x"6725",
			x"0000" when x"6726",
			x"0000" when x"6727",
			x"0000" when x"6728",
			x"0000" when x"6729",
			x"0000" when x"672A",
			x"0000" when x"672B",
			x"0000" when x"672C",
			x"0000" when x"672D",
			x"0000" when x"672E",
			x"0000" when x"672F",
			x"0000" when x"6730",
			x"0000" when x"6731",
			x"0000" when x"6732",
			x"0000" when x"6733",
			x"0000" when x"6734",
			x"0000" when x"6735",
			x"0000" when x"6736",
			x"0000" when x"6737",
			x"0000" when x"6738",
			x"0000" when x"6739",
			x"0000" when x"673A",
			x"0000" when x"673B",
			x"0000" when x"673C",
			x"0000" when x"673D",
			x"0000" when x"673E",
			x"0000" when x"673F",
			x"0000" when x"6740",
			x"0000" when x"6741",
			x"0000" when x"6742",
			x"0000" when x"6743",
			x"0000" when x"6744",
			x"0000" when x"6745",
			x"0000" when x"6746",
			x"0000" when x"6747",
			x"0000" when x"6748",
			x"0000" when x"6749",
			x"0000" when x"674A",
			x"0000" when x"674B",
			x"0000" when x"674C",
			x"0000" when x"674D",
			x"0000" when x"674E",
			x"0000" when x"674F",
			x"0000" when x"6750",
			x"0000" when x"6751",
			x"0000" when x"6752",
			x"0000" when x"6753",
			x"0000" when x"6754",
			x"0000" when x"6755",
			x"0000" when x"6756",
			x"0000" when x"6757",
			x"0000" when x"6758",
			x"0000" when x"6759",
			x"0000" when x"675A",
			x"0000" when x"675B",
			x"0000" when x"675C",
			x"0000" when x"675D",
			x"0000" when x"675E",
			x"0000" when x"675F",
			x"0000" when x"6760",
			x"0000" when x"6761",
			x"0000" when x"6762",
			x"0000" when x"6763",
			x"0000" when x"6764",
			x"0000" when x"6765",
			x"0000" when x"6766",
			x"0000" when x"6767",
			x"0000" when x"6768",
			x"0000" when x"6769",
			x"0000" when x"676A",
			x"0000" when x"676B",
			x"0000" when x"676C",
			x"0000" when x"676D",
			x"0000" when x"676E",
			x"0000" when x"676F",
			x"0000" when x"6770",
			x"0000" when x"6771",
			x"0000" when x"6772",
			x"0000" when x"6773",
			x"0000" when x"6774",
			x"0000" when x"6775",
			x"0000" when x"6776",
			x"0000" when x"6777",
			x"0000" when x"6778",
			x"0000" when x"6779",
			x"0000" when x"677A",
			x"0000" when x"677B",
			x"0000" when x"677C",
			x"0000" when x"677D",
			x"0000" when x"677E",
			x"0000" when x"677F",
			x"0000" when x"6780",
			x"0000" when x"6781",
			x"0000" when x"6782",
			x"0000" when x"6783",
			x"0000" when x"6784",
			x"0000" when x"6785",
			x"0000" when x"6786",
			x"0000" when x"6787",
			x"0000" when x"6788",
			x"0000" when x"6789",
			x"0000" when x"678A",
			x"0000" when x"678B",
			x"0000" when x"678C",
			x"0000" when x"678D",
			x"0000" when x"678E",
			x"0000" when x"678F",
			x"0000" when x"6790",
			x"0000" when x"6791",
			x"0000" when x"6792",
			x"0000" when x"6793",
			x"0000" when x"6794",
			x"0000" when x"6795",
			x"0000" when x"6796",
			x"0000" when x"6797",
			x"0000" when x"6798",
			x"0000" when x"6799",
			x"0000" when x"679A",
			x"0000" when x"679B",
			x"0000" when x"679C",
			x"0000" when x"679D",
			x"0000" when x"679E",
			x"0000" when x"679F",
			x"0000" when x"67A0",
			x"0000" when x"67A1",
			x"0000" when x"67A2",
			x"0000" when x"67A3",
			x"0000" when x"67A4",
			x"0000" when x"67A5",
			x"0000" when x"67A6",
			x"0000" when x"67A7",
			x"0000" when x"67A8",
			x"0000" when x"67A9",
			x"0000" when x"67AA",
			x"0000" when x"67AB",
			x"0000" when x"67AC",
			x"0000" when x"67AD",
			x"0000" when x"67AE",
			x"0000" when x"67AF",
			x"0000" when x"67B0",
			x"0000" when x"67B1",
			x"0000" when x"67B2",
			x"0000" when x"67B3",
			x"0000" when x"67B4",
			x"0000" when x"67B5",
			x"0000" when x"67B6",
			x"0000" when x"67B7",
			x"0000" when x"67B8",
			x"0000" when x"67B9",
			x"0000" when x"67BA",
			x"0000" when x"67BB",
			x"0000" when x"67BC",
			x"0000" when x"67BD",
			x"0000" when x"67BE",
			x"0000" when x"67BF",
			x"0000" when x"67C0",
			x"0000" when x"67C1",
			x"0000" when x"67C2",
			x"0000" when x"67C3",
			x"0000" when x"67C4",
			x"0000" when x"67C5",
			x"0000" when x"67C6",
			x"0000" when x"67C7",
			x"0000" when x"67C8",
			x"0000" when x"67C9",
			x"0000" when x"67CA",
			x"0000" when x"67CB",
			x"0000" when x"67CC",
			x"0000" when x"67CD",
			x"0000" when x"67CE",
			x"0000" when x"67CF",
			x"0000" when x"67D0",
			x"0000" when x"67D1",
			x"0000" when x"67D2",
			x"0000" when x"67D3",
			x"0000" when x"67D4",
			x"0000" when x"67D5",
			x"0000" when x"67D6",
			x"0000" when x"67D7",
			x"0000" when x"67D8",
			x"0000" when x"67D9",
			x"0000" when x"67DA",
			x"0000" when x"67DB",
			x"0000" when x"67DC",
			x"0000" when x"67DD",
			x"0000" when x"67DE",
			x"0000" when x"67DF",
			x"0000" when x"67E0",
			x"0000" when x"67E1",
			x"0000" when x"67E2",
			x"0000" when x"67E3",
			x"0000" when x"67E4",
			x"0000" when x"67E5",
			x"0000" when x"67E6",
			x"0000" when x"67E7",
			x"0000" when x"67E8",
			x"0000" when x"67E9",
			x"0000" when x"67EA",
			x"0000" when x"67EB",
			x"0000" when x"67EC",
			x"0000" when x"67ED",
			x"0000" when x"67EE",
			x"0000" when x"67EF",
			x"0000" when x"67F0",
			x"0000" when x"67F1",
			x"0000" when x"67F2",
			x"0000" when x"67F3",
			x"0000" when x"67F4",
			x"0000" when x"67F5",
			x"0000" when x"67F6",
			x"0000" when x"67F7",
			x"0000" when x"67F8",
			x"0000" when x"67F9",
			x"0000" when x"67FA",
			x"0000" when x"67FB",
			x"0000" when x"67FC",
			x"0000" when x"67FD",
			x"0000" when x"67FE",
			x"0000" when x"67FF",
			x"0000" when x"6800",
			x"0000" when x"6801",
			x"0000" when x"6802",
			x"0000" when x"6803",
			x"0000" when x"6804",
			x"0000" when x"6805",
			x"0000" when x"6806",
			x"0000" when x"6807",
			x"0000" when x"6808",
			x"0000" when x"6809",
			x"0000" when x"680A",
			x"0000" when x"680B",
			x"0000" when x"680C",
			x"0000" when x"680D",
			x"0000" when x"680E",
			x"0000" when x"680F",
			x"0000" when x"6810",
			x"0000" when x"6811",
			x"0000" when x"6812",
			x"0000" when x"6813",
			x"0000" when x"6814",
			x"0000" when x"6815",
			x"0000" when x"6816",
			x"0000" when x"6817",
			x"0000" when x"6818",
			x"0000" when x"6819",
			x"0000" when x"681A",
			x"0000" when x"681B",
			x"0000" when x"681C",
			x"0000" when x"681D",
			x"0000" when x"681E",
			x"0000" when x"681F",
			x"0000" when x"6820",
			x"0000" when x"6821",
			x"0000" when x"6822",
			x"0000" when x"6823",
			x"0000" when x"6824",
			x"0000" when x"6825",
			x"0000" when x"6826",
			x"0000" when x"6827",
			x"0000" when x"6828",
			x"0000" when x"6829",
			x"0000" when x"682A",
			x"0000" when x"682B",
			x"0000" when x"682C",
			x"0000" when x"682D",
			x"0000" when x"682E",
			x"0000" when x"682F",
			x"0000" when x"6830",
			x"0000" when x"6831",
			x"0000" when x"6832",
			x"0000" when x"6833",
			x"0000" when x"6834",
			x"0000" when x"6835",
			x"0000" when x"6836",
			x"0000" when x"6837",
			x"0000" when x"6838",
			x"0000" when x"6839",
			x"0000" when x"683A",
			x"0000" when x"683B",
			x"0000" when x"683C",
			x"0000" when x"683D",
			x"0000" when x"683E",
			x"0000" when x"683F",
			x"0000" when x"6840",
			x"0000" when x"6841",
			x"0000" when x"6842",
			x"0000" when x"6843",
			x"0000" when x"6844",
			x"0000" when x"6845",
			x"0000" when x"6846",
			x"0000" when x"6847",
			x"0000" when x"6848",
			x"0000" when x"6849",
			x"0000" when x"684A",
			x"0000" when x"684B",
			x"0000" when x"684C",
			x"0000" when x"684D",
			x"0000" when x"684E",
			x"0000" when x"684F",
			x"0000" when x"6850",
			x"0000" when x"6851",
			x"0000" when x"6852",
			x"0000" when x"6853",
			x"0000" when x"6854",
			x"0000" when x"6855",
			x"0000" when x"6856",
			x"0000" when x"6857",
			x"0000" when x"6858",
			x"0000" when x"6859",
			x"0000" when x"685A",
			x"0000" when x"685B",
			x"0000" when x"685C",
			x"0000" when x"685D",
			x"0000" when x"685E",
			x"0000" when x"685F",
			x"0000" when x"6860",
			x"0000" when x"6861",
			x"0000" when x"6862",
			x"0000" when x"6863",
			x"0000" when x"6864",
			x"0000" when x"6865",
			x"0000" when x"6866",
			x"0000" when x"6867",
			x"0000" when x"6868",
			x"0000" when x"6869",
			x"0000" when x"686A",
			x"0000" when x"686B",
			x"0000" when x"686C",
			x"0000" when x"686D",
			x"0000" when x"686E",
			x"0000" when x"686F",
			x"0000" when x"6870",
			x"0000" when x"6871",
			x"0000" when x"6872",
			x"0000" when x"6873",
			x"0000" when x"6874",
			x"0000" when x"6875",
			x"0000" when x"6876",
			x"0000" when x"6877",
			x"0000" when x"6878",
			x"0000" when x"6879",
			x"0000" when x"687A",
			x"0000" when x"687B",
			x"0000" when x"687C",
			x"0000" when x"687D",
			x"0000" when x"687E",
			x"0000" when x"687F",
			x"0000" when x"6880",
			x"0000" when x"6881",
			x"0000" when x"6882",
			x"0000" when x"6883",
			x"0000" when x"6884",
			x"0000" when x"6885",
			x"0000" when x"6886",
			x"0000" when x"6887",
			x"0000" when x"6888",
			x"0000" when x"6889",
			x"0000" when x"688A",
			x"0000" when x"688B",
			x"0000" when x"688C",
			x"0000" when x"688D",
			x"0000" when x"688E",
			x"0000" when x"688F",
			x"0000" when x"6890",
			x"0000" when x"6891",
			x"0000" when x"6892",
			x"0000" when x"6893",
			x"0000" when x"6894",
			x"0000" when x"6895",
			x"0000" when x"6896",
			x"0000" when x"6897",
			x"0000" when x"6898",
			x"0000" when x"6899",
			x"0000" when x"689A",
			x"0000" when x"689B",
			x"0000" when x"689C",
			x"0000" when x"689D",
			x"0000" when x"689E",
			x"0000" when x"689F",
			x"0000" when x"68A0",
			x"0000" when x"68A1",
			x"0000" when x"68A2",
			x"0000" when x"68A3",
			x"0000" when x"68A4",
			x"0000" when x"68A5",
			x"0000" when x"68A6",
			x"0000" when x"68A7",
			x"0000" when x"68A8",
			x"0000" when x"68A9",
			x"0000" when x"68AA",
			x"0000" when x"68AB",
			x"0000" when x"68AC",
			x"0000" when x"68AD",
			x"0000" when x"68AE",
			x"0000" when x"68AF",
			x"0000" when x"68B0",
			x"0000" when x"68B1",
			x"0000" when x"68B2",
			x"0000" when x"68B3",
			x"0000" when x"68B4",
			x"0000" when x"68B5",
			x"0000" when x"68B6",
			x"0000" when x"68B7",
			x"0000" when x"68B8",
			x"0000" when x"68B9",
			x"0000" when x"68BA",
			x"0000" when x"68BB",
			x"0000" when x"68BC",
			x"0000" when x"68BD",
			x"0000" when x"68BE",
			x"0000" when x"68BF",
			x"0000" when x"68C0",
			x"0000" when x"68C1",
			x"0000" when x"68C2",
			x"0000" when x"68C3",
			x"0000" when x"68C4",
			x"0000" when x"68C5",
			x"0000" when x"68C6",
			x"0000" when x"68C7",
			x"0000" when x"68C8",
			x"0000" when x"68C9",
			x"0000" when x"68CA",
			x"0000" when x"68CB",
			x"0000" when x"68CC",
			x"0000" when x"68CD",
			x"0000" when x"68CE",
			x"0000" when x"68CF",
			x"0000" when x"68D0",
			x"0000" when x"68D1",
			x"0000" when x"68D2",
			x"0000" when x"68D3",
			x"0000" when x"68D4",
			x"0000" when x"68D5",
			x"0000" when x"68D6",
			x"0000" when x"68D7",
			x"0000" when x"68D8",
			x"0000" when x"68D9",
			x"0000" when x"68DA",
			x"0000" when x"68DB",
			x"0000" when x"68DC",
			x"0000" when x"68DD",
			x"0000" when x"68DE",
			x"0000" when x"68DF",
			x"0000" when x"68E0",
			x"0000" when x"68E1",
			x"0000" when x"68E2",
			x"0000" when x"68E3",
			x"0000" when x"68E4",
			x"0000" when x"68E5",
			x"0000" when x"68E6",
			x"0000" when x"68E7",
			x"0000" when x"68E8",
			x"0000" when x"68E9",
			x"0000" when x"68EA",
			x"0000" when x"68EB",
			x"0000" when x"68EC",
			x"0000" when x"68ED",
			x"0000" when x"68EE",
			x"0000" when x"68EF",
			x"0000" when x"68F0",
			x"0000" when x"68F1",
			x"0000" when x"68F2",
			x"0000" when x"68F3",
			x"0000" when x"68F4",
			x"0000" when x"68F5",
			x"0000" when x"68F6",
			x"0000" when x"68F7",
			x"0000" when x"68F8",
			x"0000" when x"68F9",
			x"0000" when x"68FA",
			x"0000" when x"68FB",
			x"0000" when x"68FC",
			x"0000" when x"68FD",
			x"0000" when x"68FE",
			x"0000" when x"68FF",
			x"0000" when x"6900",
			x"0000" when x"6901",
			x"0000" when x"6902",
			x"0000" when x"6903",
			x"0000" when x"6904",
			x"0000" when x"6905",
			x"0000" when x"6906",
			x"0000" when x"6907",
			x"0000" when x"6908",
			x"0000" when x"6909",
			x"0000" when x"690A",
			x"0000" when x"690B",
			x"0000" when x"690C",
			x"0000" when x"690D",
			x"0000" when x"690E",
			x"0000" when x"690F",
			x"0000" when x"6910",
			x"0000" when x"6911",
			x"0000" when x"6912",
			x"0000" when x"6913",
			x"0000" when x"6914",
			x"0000" when x"6915",
			x"0000" when x"6916",
			x"0000" when x"6917",
			x"0000" when x"6918",
			x"0000" when x"6919",
			x"0000" when x"691A",
			x"0000" when x"691B",
			x"0000" when x"691C",
			x"0000" when x"691D",
			x"0000" when x"691E",
			x"0000" when x"691F",
			x"0000" when x"6920",
			x"0000" when x"6921",
			x"0000" when x"6922",
			x"0000" when x"6923",
			x"0000" when x"6924",
			x"0000" when x"6925",
			x"0000" when x"6926",
			x"0000" when x"6927",
			x"0000" when x"6928",
			x"0000" when x"6929",
			x"0000" when x"692A",
			x"0000" when x"692B",
			x"0000" when x"692C",
			x"0000" when x"692D",
			x"0000" when x"692E",
			x"0000" when x"692F",
			x"0000" when x"6930",
			x"0000" when x"6931",
			x"0000" when x"6932",
			x"0000" when x"6933",
			x"0000" when x"6934",
			x"0000" when x"6935",
			x"0000" when x"6936",
			x"0000" when x"6937",
			x"0000" when x"6938",
			x"0000" when x"6939",
			x"0000" when x"693A",
			x"0000" when x"693B",
			x"0000" when x"693C",
			x"0000" when x"693D",
			x"0000" when x"693E",
			x"0000" when x"693F",
			x"0000" when x"6940",
			x"0000" when x"6941",
			x"0000" when x"6942",
			x"0000" when x"6943",
			x"0000" when x"6944",
			x"0000" when x"6945",
			x"0000" when x"6946",
			x"0000" when x"6947",
			x"0000" when x"6948",
			x"0000" when x"6949",
			x"0000" when x"694A",
			x"0000" when x"694B",
			x"0000" when x"694C",
			x"0000" when x"694D",
			x"0000" when x"694E",
			x"0000" when x"694F",
			x"0000" when x"6950",
			x"0000" when x"6951",
			x"0000" when x"6952",
			x"0000" when x"6953",
			x"0000" when x"6954",
			x"0000" when x"6955",
			x"0000" when x"6956",
			x"0000" when x"6957",
			x"0000" when x"6958",
			x"0000" when x"6959",
			x"0000" when x"695A",
			x"0000" when x"695B",
			x"0000" when x"695C",
			x"0000" when x"695D",
			x"0000" when x"695E",
			x"0000" when x"695F",
			x"0000" when x"6960",
			x"0000" when x"6961",
			x"0000" when x"6962",
			x"0000" when x"6963",
			x"0000" when x"6964",
			x"0000" when x"6965",
			x"0000" when x"6966",
			x"0000" when x"6967",
			x"0000" when x"6968",
			x"0000" when x"6969",
			x"0000" when x"696A",
			x"0000" when x"696B",
			x"0000" when x"696C",
			x"0000" when x"696D",
			x"0000" when x"696E",
			x"0000" when x"696F",
			x"0000" when x"6970",
			x"0000" when x"6971",
			x"0000" when x"6972",
			x"0000" when x"6973",
			x"0000" when x"6974",
			x"0000" when x"6975",
			x"0000" when x"6976",
			x"0000" when x"6977",
			x"0000" when x"6978",
			x"0000" when x"6979",
			x"0000" when x"697A",
			x"0000" when x"697B",
			x"0000" when x"697C",
			x"0000" when x"697D",
			x"0000" when x"697E",
			x"0000" when x"697F",
			x"0000" when x"6980",
			x"0000" when x"6981",
			x"0000" when x"6982",
			x"0000" when x"6983",
			x"0000" when x"6984",
			x"0000" when x"6985",
			x"0000" when x"6986",
			x"0000" when x"6987",
			x"0000" when x"6988",
			x"0000" when x"6989",
			x"0000" when x"698A",
			x"0000" when x"698B",
			x"0000" when x"698C",
			x"0000" when x"698D",
			x"0000" when x"698E",
			x"0000" when x"698F",
			x"0000" when x"6990",
			x"0000" when x"6991",
			x"0000" when x"6992",
			x"0000" when x"6993",
			x"0000" when x"6994",
			x"0000" when x"6995",
			x"0000" when x"6996",
			x"0000" when x"6997",
			x"0000" when x"6998",
			x"0000" when x"6999",
			x"0000" when x"699A",
			x"0000" when x"699B",
			x"0000" when x"699C",
			x"0000" when x"699D",
			x"0000" when x"699E",
			x"0000" when x"699F",
			x"0000" when x"69A0",
			x"0000" when x"69A1",
			x"0000" when x"69A2",
			x"0000" when x"69A3",
			x"0000" when x"69A4",
			x"0000" when x"69A5",
			x"0000" when x"69A6",
			x"0000" when x"69A7",
			x"0000" when x"69A8",
			x"0000" when x"69A9",
			x"0000" when x"69AA",
			x"0000" when x"69AB",
			x"0000" when x"69AC",
			x"0000" when x"69AD",
			x"0000" when x"69AE",
			x"0000" when x"69AF",
			x"0000" when x"69B0",
			x"0000" when x"69B1",
			x"0000" when x"69B2",
			x"0000" when x"69B3",
			x"0000" when x"69B4",
			x"0000" when x"69B5",
			x"0000" when x"69B6",
			x"0000" when x"69B7",
			x"0000" when x"69B8",
			x"0000" when x"69B9",
			x"0000" when x"69BA",
			x"0000" when x"69BB",
			x"0000" when x"69BC",
			x"0000" when x"69BD",
			x"0000" when x"69BE",
			x"0000" when x"69BF",
			x"0000" when x"69C0",
			x"0000" when x"69C1",
			x"0000" when x"69C2",
			x"0000" when x"69C3",
			x"0000" when x"69C4",
			x"0000" when x"69C5",
			x"0000" when x"69C6",
			x"0000" when x"69C7",
			x"0000" when x"69C8",
			x"0000" when x"69C9",
			x"0000" when x"69CA",
			x"0000" when x"69CB",
			x"0000" when x"69CC",
			x"0000" when x"69CD",
			x"0000" when x"69CE",
			x"0000" when x"69CF",
			x"0000" when x"69D0",
			x"0000" when x"69D1",
			x"0000" when x"69D2",
			x"0000" when x"69D3",
			x"0000" when x"69D4",
			x"0000" when x"69D5",
			x"0000" when x"69D6",
			x"0000" when x"69D7",
			x"0000" when x"69D8",
			x"0000" when x"69D9",
			x"0000" when x"69DA",
			x"0000" when x"69DB",
			x"0000" when x"69DC",
			x"0000" when x"69DD",
			x"0000" when x"69DE",
			x"0000" when x"69DF",
			x"0000" when x"69E0",
			x"0000" when x"69E1",
			x"0000" when x"69E2",
			x"0000" when x"69E3",
			x"0000" when x"69E4",
			x"0000" when x"69E5",
			x"0000" when x"69E6",
			x"0000" when x"69E7",
			x"0000" when x"69E8",
			x"0000" when x"69E9",
			x"0000" when x"69EA",
			x"0000" when x"69EB",
			x"0000" when x"69EC",
			x"0000" when x"69ED",
			x"0000" when x"69EE",
			x"0000" when x"69EF",
			x"0000" when x"69F0",
			x"0000" when x"69F1",
			x"0000" when x"69F2",
			x"0000" when x"69F3",
			x"0000" when x"69F4",
			x"0000" when x"69F5",
			x"0000" when x"69F6",
			x"0000" when x"69F7",
			x"0000" when x"69F8",
			x"0000" when x"69F9",
			x"0000" when x"69FA",
			x"0000" when x"69FB",
			x"0000" when x"69FC",
			x"0000" when x"69FD",
			x"0000" when x"69FE",
			x"0000" when x"69FF",
			x"0000" when x"6A00",
			x"0000" when x"6A01",
			x"0000" when x"6A02",
			x"0000" when x"6A03",
			x"0000" when x"6A04",
			x"0000" when x"6A05",
			x"0000" when x"6A06",
			x"0000" when x"6A07",
			x"0000" when x"6A08",
			x"0000" when x"6A09",
			x"0000" when x"6A0A",
			x"0000" when x"6A0B",
			x"0000" when x"6A0C",
			x"0000" when x"6A0D",
			x"0000" when x"6A0E",
			x"0000" when x"6A0F",
			x"0000" when x"6A10",
			x"0000" when x"6A11",
			x"0000" when x"6A12",
			x"0000" when x"6A13",
			x"0000" when x"6A14",
			x"0000" when x"6A15",
			x"0000" when x"6A16",
			x"0000" when x"6A17",
			x"0000" when x"6A18",
			x"0000" when x"6A19",
			x"0000" when x"6A1A",
			x"0000" when x"6A1B",
			x"0000" when x"6A1C",
			x"0000" when x"6A1D",
			x"0000" when x"6A1E",
			x"0000" when x"6A1F",
			x"0000" when x"6A20",
			x"0000" when x"6A21",
			x"0000" when x"6A22",
			x"0000" when x"6A23",
			x"0000" when x"6A24",
			x"0000" when x"6A25",
			x"0000" when x"6A26",
			x"0000" when x"6A27",
			x"0000" when x"6A28",
			x"0000" when x"6A29",
			x"0000" when x"6A2A",
			x"0000" when x"6A2B",
			x"0000" when x"6A2C",
			x"0000" when x"6A2D",
			x"0000" when x"6A2E",
			x"0000" when x"6A2F",
			x"0000" when x"6A30",
			x"0000" when x"6A31",
			x"0000" when x"6A32",
			x"0000" when x"6A33",
			x"0000" when x"6A34",
			x"0000" when x"6A35",
			x"0000" when x"6A36",
			x"0000" when x"6A37",
			x"0000" when x"6A38",
			x"0000" when x"6A39",
			x"0000" when x"6A3A",
			x"0000" when x"6A3B",
			x"0000" when x"6A3C",
			x"0000" when x"6A3D",
			x"0000" when x"6A3E",
			x"0000" when x"6A3F",
			x"0000" when x"6A40",
			x"0000" when x"6A41",
			x"0000" when x"6A42",
			x"0000" when x"6A43",
			x"0000" when x"6A44",
			x"0000" when x"6A45",
			x"0000" when x"6A46",
			x"0000" when x"6A47",
			x"0000" when x"6A48",
			x"0000" when x"6A49",
			x"0000" when x"6A4A",
			x"0000" when x"6A4B",
			x"0000" when x"6A4C",
			x"0000" when x"6A4D",
			x"0000" when x"6A4E",
			x"0000" when x"6A4F",
			x"0000" when x"6A50",
			x"0000" when x"6A51",
			x"0000" when x"6A52",
			x"0000" when x"6A53",
			x"0000" when x"6A54",
			x"0000" when x"6A55",
			x"0000" when x"6A56",
			x"0000" when x"6A57",
			x"0000" when x"6A58",
			x"0000" when x"6A59",
			x"0000" when x"6A5A",
			x"0000" when x"6A5B",
			x"0000" when x"6A5C",
			x"0000" when x"6A5D",
			x"0000" when x"6A5E",
			x"0000" when x"6A5F",
			x"0000" when x"6A60",
			x"0000" when x"6A61",
			x"0000" when x"6A62",
			x"0000" when x"6A63",
			x"0000" when x"6A64",
			x"0000" when x"6A65",
			x"0000" when x"6A66",
			x"0000" when x"6A67",
			x"0000" when x"6A68",
			x"0000" when x"6A69",
			x"0000" when x"6A6A",
			x"0000" when x"6A6B",
			x"0000" when x"6A6C",
			x"0000" when x"6A6D",
			x"0000" when x"6A6E",
			x"0000" when x"6A6F",
			x"0000" when x"6A70",
			x"0000" when x"6A71",
			x"0000" when x"6A72",
			x"0000" when x"6A73",
			x"0000" when x"6A74",
			x"0000" when x"6A75",
			x"0000" when x"6A76",
			x"0000" when x"6A77",
			x"0000" when x"6A78",
			x"0000" when x"6A79",
			x"0000" when x"6A7A",
			x"0000" when x"6A7B",
			x"0000" when x"6A7C",
			x"0000" when x"6A7D",
			x"0000" when x"6A7E",
			x"0000" when x"6A7F",
			x"0000" when x"6A80",
			x"0000" when x"6A81",
			x"0000" when x"6A82",
			x"0000" when x"6A83",
			x"0000" when x"6A84",
			x"0000" when x"6A85",
			x"0000" when x"6A86",
			x"0000" when x"6A87",
			x"0000" when x"6A88",
			x"0000" when x"6A89",
			x"0000" when x"6A8A",
			x"0000" when x"6A8B",
			x"0000" when x"6A8C",
			x"0000" when x"6A8D",
			x"0000" when x"6A8E",
			x"0000" when x"6A8F",
			x"0000" when x"6A90",
			x"0000" when x"6A91",
			x"0000" when x"6A92",
			x"0000" when x"6A93",
			x"0000" when x"6A94",
			x"0000" when x"6A95",
			x"0000" when x"6A96",
			x"0000" when x"6A97",
			x"0000" when x"6A98",
			x"0000" when x"6A99",
			x"0000" when x"6A9A",
			x"0000" when x"6A9B",
			x"0000" when x"6A9C",
			x"0000" when x"6A9D",
			x"0000" when x"6A9E",
			x"0000" when x"6A9F",
			x"0000" when x"6AA0",
			x"0000" when x"6AA1",
			x"0000" when x"6AA2",
			x"0000" when x"6AA3",
			x"0000" when x"6AA4",
			x"0000" when x"6AA5",
			x"0000" when x"6AA6",
			x"0000" when x"6AA7",
			x"0000" when x"6AA8",
			x"0000" when x"6AA9",
			x"0000" when x"6AAA",
			x"0000" when x"6AAB",
			x"0000" when x"6AAC",
			x"0000" when x"6AAD",
			x"0000" when x"6AAE",
			x"0000" when x"6AAF",
			x"0000" when x"6AB0",
			x"0000" when x"6AB1",
			x"0000" when x"6AB2",
			x"0000" when x"6AB3",
			x"0000" when x"6AB4",
			x"0000" when x"6AB5",
			x"0000" when x"6AB6",
			x"0000" when x"6AB7",
			x"0000" when x"6AB8",
			x"0000" when x"6AB9",
			x"0000" when x"6ABA",
			x"0000" when x"6ABB",
			x"0000" when x"6ABC",
			x"0000" when x"6ABD",
			x"0000" when x"6ABE",
			x"0000" when x"6ABF",
			x"0000" when x"6AC0",
			x"0000" when x"6AC1",
			x"0000" when x"6AC2",
			x"0000" when x"6AC3",
			x"0000" when x"6AC4",
			x"0000" when x"6AC5",
			x"0000" when x"6AC6",
			x"0000" when x"6AC7",
			x"0000" when x"6AC8",
			x"0000" when x"6AC9",
			x"0000" when x"6ACA",
			x"0000" when x"6ACB",
			x"0000" when x"6ACC",
			x"0000" when x"6ACD",
			x"0000" when x"6ACE",
			x"0000" when x"6ACF",
			x"0000" when x"6AD0",
			x"0000" when x"6AD1",
			x"0000" when x"6AD2",
			x"0000" when x"6AD3",
			x"0000" when x"6AD4",
			x"0000" when x"6AD5",
			x"0000" when x"6AD6",
			x"0000" when x"6AD7",
			x"0000" when x"6AD8",
			x"0000" when x"6AD9",
			x"0000" when x"6ADA",
			x"0000" when x"6ADB",
			x"0000" when x"6ADC",
			x"0000" when x"6ADD",
			x"0000" when x"6ADE",
			x"0000" when x"6ADF",
			x"0000" when x"6AE0",
			x"0000" when x"6AE1",
			x"0000" when x"6AE2",
			x"0000" when x"6AE3",
			x"0000" when x"6AE4",
			x"0000" when x"6AE5",
			x"0000" when x"6AE6",
			x"0000" when x"6AE7",
			x"0000" when x"6AE8",
			x"0000" when x"6AE9",
			x"0000" when x"6AEA",
			x"0000" when x"6AEB",
			x"0000" when x"6AEC",
			x"0000" when x"6AED",
			x"0000" when x"6AEE",
			x"0000" when x"6AEF",
			x"0000" when x"6AF0",
			x"0000" when x"6AF1",
			x"0000" when x"6AF2",
			x"0000" when x"6AF3",
			x"0000" when x"6AF4",
			x"0000" when x"6AF5",
			x"0000" when x"6AF6",
			x"0000" when x"6AF7",
			x"0000" when x"6AF8",
			x"0000" when x"6AF9",
			x"0000" when x"6AFA",
			x"0000" when x"6AFB",
			x"0000" when x"6AFC",
			x"0000" when x"6AFD",
			x"0000" when x"6AFE",
			x"0000" when x"6AFF",
			x"0000" when x"6B00",
			x"0000" when x"6B01",
			x"0000" when x"6B02",
			x"0000" when x"6B03",
			x"0000" when x"6B04",
			x"0000" when x"6B05",
			x"0000" when x"6B06",
			x"0000" when x"6B07",
			x"0000" when x"6B08",
			x"0000" when x"6B09",
			x"0000" when x"6B0A",
			x"0000" when x"6B0B",
			x"0000" when x"6B0C",
			x"0000" when x"6B0D",
			x"0000" when x"6B0E",
			x"0000" when x"6B0F",
			x"0000" when x"6B10",
			x"0000" when x"6B11",
			x"0000" when x"6B12",
			x"0000" when x"6B13",
			x"0000" when x"6B14",
			x"0000" when x"6B15",
			x"0000" when x"6B16",
			x"0000" when x"6B17",
			x"0000" when x"6B18",
			x"0000" when x"6B19",
			x"0000" when x"6B1A",
			x"0000" when x"6B1B",
			x"0000" when x"6B1C",
			x"0000" when x"6B1D",
			x"0000" when x"6B1E",
			x"0000" when x"6B1F",
			x"0000" when x"6B20",
			x"0000" when x"6B21",
			x"0000" when x"6B22",
			x"0000" when x"6B23",
			x"0000" when x"6B24",
			x"0000" when x"6B25",
			x"0000" when x"6B26",
			x"0000" when x"6B27",
			x"0000" when x"6B28",
			x"0000" when x"6B29",
			x"0000" when x"6B2A",
			x"0000" when x"6B2B",
			x"0000" when x"6B2C",
			x"0000" when x"6B2D",
			x"0000" when x"6B2E",
			x"0000" when x"6B2F",
			x"0000" when x"6B30",
			x"0000" when x"6B31",
			x"0000" when x"6B32",
			x"0000" when x"6B33",
			x"0000" when x"6B34",
			x"0000" when x"6B35",
			x"0000" when x"6B36",
			x"0000" when x"6B37",
			x"0000" when x"6B38",
			x"0000" when x"6B39",
			x"0000" when x"6B3A",
			x"0000" when x"6B3B",
			x"0000" when x"6B3C",
			x"0000" when x"6B3D",
			x"0000" when x"6B3E",
			x"0000" when x"6B3F",
			x"0000" when x"6B40",
			x"0000" when x"6B41",
			x"0000" when x"6B42",
			x"0000" when x"6B43",
			x"0000" when x"6B44",
			x"0000" when x"6B45",
			x"0000" when x"6B46",
			x"0000" when x"6B47",
			x"0000" when x"6B48",
			x"0000" when x"6B49",
			x"0000" when x"6B4A",
			x"0000" when x"6B4B",
			x"0000" when x"6B4C",
			x"0000" when x"6B4D",
			x"0000" when x"6B4E",
			x"0000" when x"6B4F",
			x"0000" when x"6B50",
			x"0000" when x"6B51",
			x"0000" when x"6B52",
			x"0000" when x"6B53",
			x"0000" when x"6B54",
			x"0000" when x"6B55",
			x"0000" when x"6B56",
			x"0000" when x"6B57",
			x"0000" when x"6B58",
			x"0000" when x"6B59",
			x"0000" when x"6B5A",
			x"0000" when x"6B5B",
			x"0000" when x"6B5C",
			x"0000" when x"6B5D",
			x"0000" when x"6B5E",
			x"0000" when x"6B5F",
			x"0000" when x"6B60",
			x"0000" when x"6B61",
			x"0000" when x"6B62",
			x"0000" when x"6B63",
			x"0000" when x"6B64",
			x"0000" when x"6B65",
			x"0000" when x"6B66",
			x"0000" when x"6B67",
			x"0000" when x"6B68",
			x"0000" when x"6B69",
			x"0000" when x"6B6A",
			x"0000" when x"6B6B",
			x"0000" when x"6B6C",
			x"0000" when x"6B6D",
			x"0000" when x"6B6E",
			x"0000" when x"6B6F",
			x"0000" when x"6B70",
			x"0000" when x"6B71",
			x"0000" when x"6B72",
			x"0000" when x"6B73",
			x"0000" when x"6B74",
			x"0000" when x"6B75",
			x"0000" when x"6B76",
			x"0000" when x"6B77",
			x"0000" when x"6B78",
			x"0000" when x"6B79",
			x"0000" when x"6B7A",
			x"0000" when x"6B7B",
			x"0000" when x"6B7C",
			x"0000" when x"6B7D",
			x"0000" when x"6B7E",
			x"0000" when x"6B7F",
			x"0000" when x"6B80",
			x"0000" when x"6B81",
			x"0000" when x"6B82",
			x"0000" when x"6B83",
			x"0000" when x"6B84",
			x"0000" when x"6B85",
			x"0000" when x"6B86",
			x"0000" when x"6B87",
			x"0000" when x"6B88",
			x"0000" when x"6B89",
			x"0000" when x"6B8A",
			x"0000" when x"6B8B",
			x"0000" when x"6B8C",
			x"0000" when x"6B8D",
			x"0000" when x"6B8E",
			x"0000" when x"6B8F",
			x"0000" when x"6B90",
			x"0000" when x"6B91",
			x"0000" when x"6B92",
			x"0000" when x"6B93",
			x"0000" when x"6B94",
			x"0000" when x"6B95",
			x"0000" when x"6B96",
			x"0000" when x"6B97",
			x"0000" when x"6B98",
			x"0000" when x"6B99",
			x"0000" when x"6B9A",
			x"0000" when x"6B9B",
			x"0000" when x"6B9C",
			x"0000" when x"6B9D",
			x"0000" when x"6B9E",
			x"0000" when x"6B9F",
			x"0000" when x"6BA0",
			x"0000" when x"6BA1",
			x"0000" when x"6BA2",
			x"0000" when x"6BA3",
			x"0000" when x"6BA4",
			x"0000" when x"6BA5",
			x"0000" when x"6BA6",
			x"0000" when x"6BA7",
			x"0000" when x"6BA8",
			x"0000" when x"6BA9",
			x"0000" when x"6BAA",
			x"0000" when x"6BAB",
			x"0000" when x"6BAC",
			x"0000" when x"6BAD",
			x"0000" when x"6BAE",
			x"0000" when x"6BAF",
			x"0000" when x"6BB0",
			x"0000" when x"6BB1",
			x"0000" when x"6BB2",
			x"0000" when x"6BB3",
			x"0000" when x"6BB4",
			x"0000" when x"6BB5",
			x"0000" when x"6BB6",
			x"0000" when x"6BB7",
			x"0000" when x"6BB8",
			x"0000" when x"6BB9",
			x"0000" when x"6BBA",
			x"0000" when x"6BBB",
			x"0000" when x"6BBC",
			x"0000" when x"6BBD",
			x"0000" when x"6BBE",
			x"0000" when x"6BBF",
			x"0000" when x"6BC0",
			x"0000" when x"6BC1",
			x"0000" when x"6BC2",
			x"0000" when x"6BC3",
			x"0000" when x"6BC4",
			x"0000" when x"6BC5",
			x"0000" when x"6BC6",
			x"0000" when x"6BC7",
			x"0000" when x"6BC8",
			x"0000" when x"6BC9",
			x"0000" when x"6BCA",
			x"0000" when x"6BCB",
			x"0000" when x"6BCC",
			x"0000" when x"6BCD",
			x"0000" when x"6BCE",
			x"0000" when x"6BCF",
			x"0000" when x"6BD0",
			x"0000" when x"6BD1",
			x"0000" when x"6BD2",
			x"0000" when x"6BD3",
			x"0000" when x"6BD4",
			x"0000" when x"6BD5",
			x"0000" when x"6BD6",
			x"0000" when x"6BD7",
			x"0000" when x"6BD8",
			x"0000" when x"6BD9",
			x"0000" when x"6BDA",
			x"0000" when x"6BDB",
			x"0000" when x"6BDC",
			x"0000" when x"6BDD",
			x"0000" when x"6BDE",
			x"0000" when x"6BDF",
			x"0000" when x"6BE0",
			x"0000" when x"6BE1",
			x"0000" when x"6BE2",
			x"0000" when x"6BE3",
			x"0000" when x"6BE4",
			x"0000" when x"6BE5",
			x"0000" when x"6BE6",
			x"0000" when x"6BE7",
			x"0000" when x"6BE8",
			x"0000" when x"6BE9",
			x"0000" when x"6BEA",
			x"0000" when x"6BEB",
			x"0000" when x"6BEC",
			x"0000" when x"6BED",
			x"0000" when x"6BEE",
			x"0000" when x"6BEF",
			x"0000" when x"6BF0",
			x"0000" when x"6BF1",
			x"0000" when x"6BF2",
			x"0000" when x"6BF3",
			x"0000" when x"6BF4",
			x"0000" when x"6BF5",
			x"0000" when x"6BF6",
			x"0000" when x"6BF7",
			x"0000" when x"6BF8",
			x"0000" when x"6BF9",
			x"0000" when x"6BFA",
			x"0000" when x"6BFB",
			x"0000" when x"6BFC",
			x"0000" when x"6BFD",
			x"0000" when x"6BFE",
			x"0000" when x"6BFF",
			x"0000" when x"6C00",
			x"0000" when x"6C01",
			x"0000" when x"6C02",
			x"0000" when x"6C03",
			x"0000" when x"6C04",
			x"0000" when x"6C05",
			x"0000" when x"6C06",
			x"0000" when x"6C07",
			x"0000" when x"6C08",
			x"0000" when x"6C09",
			x"0000" when x"6C0A",
			x"0000" when x"6C0B",
			x"0000" when x"6C0C",
			x"0000" when x"6C0D",
			x"0000" when x"6C0E",
			x"0000" when x"6C0F",
			x"0000" when x"6C10",
			x"0000" when x"6C11",
			x"0000" when x"6C12",
			x"0000" when x"6C13",
			x"0000" when x"6C14",
			x"0000" when x"6C15",
			x"0000" when x"6C16",
			x"0000" when x"6C17",
			x"0000" when x"6C18",
			x"0000" when x"6C19",
			x"0000" when x"6C1A",
			x"0000" when x"6C1B",
			x"0000" when x"6C1C",
			x"0000" when x"6C1D",
			x"0000" when x"6C1E",
			x"0000" when x"6C1F",
			x"0000" when x"6C20",
			x"0000" when x"6C21",
			x"0000" when x"6C22",
			x"0000" when x"6C23",
			x"0000" when x"6C24",
			x"0000" when x"6C25",
			x"0000" when x"6C26",
			x"0000" when x"6C27",
			x"0000" when x"6C28",
			x"0000" when x"6C29",
			x"0000" when x"6C2A",
			x"0000" when x"6C2B",
			x"0000" when x"6C2C",
			x"0000" when x"6C2D",
			x"0000" when x"6C2E",
			x"0000" when x"6C2F",
			x"0000" when x"6C30",
			x"0000" when x"6C31",
			x"0000" when x"6C32",
			x"0000" when x"6C33",
			x"0000" when x"6C34",
			x"0000" when x"6C35",
			x"0000" when x"6C36",
			x"0000" when x"6C37",
			x"0000" when x"6C38",
			x"0000" when x"6C39",
			x"0000" when x"6C3A",
			x"0000" when x"6C3B",
			x"0000" when x"6C3C",
			x"0000" when x"6C3D",
			x"0000" when x"6C3E",
			x"0000" when x"6C3F",
			x"0000" when x"6C40",
			x"0000" when x"6C41",
			x"0000" when x"6C42",
			x"0000" when x"6C43",
			x"0000" when x"6C44",
			x"0000" when x"6C45",
			x"0000" when x"6C46",
			x"0000" when x"6C47",
			x"0000" when x"6C48",
			x"0000" when x"6C49",
			x"0000" when x"6C4A",
			x"0000" when x"6C4B",
			x"0000" when x"6C4C",
			x"0000" when x"6C4D",
			x"0000" when x"6C4E",
			x"0000" when x"6C4F",
			x"0000" when x"6C50",
			x"0000" when x"6C51",
			x"0000" when x"6C52",
			x"0000" when x"6C53",
			x"0000" when x"6C54",
			x"0000" when x"6C55",
			x"0000" when x"6C56",
			x"0000" when x"6C57",
			x"0000" when x"6C58",
			x"0000" when x"6C59",
			x"0000" when x"6C5A",
			x"0000" when x"6C5B",
			x"0000" when x"6C5C",
			x"0000" when x"6C5D",
			x"0000" when x"6C5E",
			x"0000" when x"6C5F",
			x"0000" when x"6C60",
			x"0000" when x"6C61",
			x"0000" when x"6C62",
			x"0000" when x"6C63",
			x"0000" when x"6C64",
			x"0000" when x"6C65",
			x"0000" when x"6C66",
			x"0000" when x"6C67",
			x"0000" when x"6C68",
			x"0000" when x"6C69",
			x"0000" when x"6C6A",
			x"0000" when x"6C6B",
			x"0000" when x"6C6C",
			x"0000" when x"6C6D",
			x"0000" when x"6C6E",
			x"0000" when x"6C6F",
			x"0000" when x"6C70",
			x"0000" when x"6C71",
			x"0000" when x"6C72",
			x"0000" when x"6C73",
			x"0000" when x"6C74",
			x"0000" when x"6C75",
			x"0000" when x"6C76",
			x"0000" when x"6C77",
			x"0000" when x"6C78",
			x"0000" when x"6C79",
			x"0000" when x"6C7A",
			x"0000" when x"6C7B",
			x"0000" when x"6C7C",
			x"0000" when x"6C7D",
			x"0000" when x"6C7E",
			x"0000" when x"6C7F",
			x"0000" when x"6C80",
			x"0000" when x"6C81",
			x"0000" when x"6C82",
			x"0000" when x"6C83",
			x"0000" when x"6C84",
			x"0000" when x"6C85",
			x"0000" when x"6C86",
			x"0000" when x"6C87",
			x"0000" when x"6C88",
			x"0000" when x"6C89",
			x"0000" when x"6C8A",
			x"0000" when x"6C8B",
			x"0000" when x"6C8C",
			x"0000" when x"6C8D",
			x"0000" when x"6C8E",
			x"0000" when x"6C8F",
			x"0000" when x"6C90",
			x"0000" when x"6C91",
			x"0000" when x"6C92",
			x"0000" when x"6C93",
			x"0000" when x"6C94",
			x"0000" when x"6C95",
			x"0000" when x"6C96",
			x"0000" when x"6C97",
			x"0000" when x"6C98",
			x"0000" when x"6C99",
			x"0000" when x"6C9A",
			x"0000" when x"6C9B",
			x"0000" when x"6C9C",
			x"0000" when x"6C9D",
			x"0000" when x"6C9E",
			x"0000" when x"6C9F",
			x"0000" when x"6CA0",
			x"0000" when x"6CA1",
			x"0000" when x"6CA2",
			x"0000" when x"6CA3",
			x"0000" when x"6CA4",
			x"0000" when x"6CA5",
			x"0000" when x"6CA6",
			x"0000" when x"6CA7",
			x"0000" when x"6CA8",
			x"0000" when x"6CA9",
			x"0000" when x"6CAA",
			x"0000" when x"6CAB",
			x"0000" when x"6CAC",
			x"0000" when x"6CAD",
			x"0000" when x"6CAE",
			x"0000" when x"6CAF",
			x"0000" when x"6CB0",
			x"0000" when x"6CB1",
			x"0000" when x"6CB2",
			x"0000" when x"6CB3",
			x"0000" when x"6CB4",
			x"0000" when x"6CB5",
			x"0000" when x"6CB6",
			x"0000" when x"6CB7",
			x"0000" when x"6CB8",
			x"0000" when x"6CB9",
			x"0000" when x"6CBA",
			x"0000" when x"6CBB",
			x"0000" when x"6CBC",
			x"0000" when x"6CBD",
			x"0000" when x"6CBE",
			x"0000" when x"6CBF",
			x"0000" when x"6CC0",
			x"0000" when x"6CC1",
			x"0000" when x"6CC2",
			x"0000" when x"6CC3",
			x"0000" when x"6CC4",
			x"0000" when x"6CC5",
			x"0000" when x"6CC6",
			x"0000" when x"6CC7",
			x"0000" when x"6CC8",
			x"0000" when x"6CC9",
			x"0000" when x"6CCA",
			x"0000" when x"6CCB",
			x"0000" when x"6CCC",
			x"0000" when x"6CCD",
			x"0000" when x"6CCE",
			x"0000" when x"6CCF",
			x"0000" when x"6CD0",
			x"0000" when x"6CD1",
			x"0000" when x"6CD2",
			x"0000" when x"6CD3",
			x"0000" when x"6CD4",
			x"0000" when x"6CD5",
			x"0000" when x"6CD6",
			x"0000" when x"6CD7",
			x"0000" when x"6CD8",
			x"0000" when x"6CD9",
			x"0000" when x"6CDA",
			x"0000" when x"6CDB",
			x"0000" when x"6CDC",
			x"0000" when x"6CDD",
			x"0000" when x"6CDE",
			x"0000" when x"6CDF",
			x"0000" when x"6CE0",
			x"0000" when x"6CE1",
			x"0000" when x"6CE2",
			x"0000" when x"6CE3",
			x"0000" when x"6CE4",
			x"0000" when x"6CE5",
			x"0000" when x"6CE6",
			x"0000" when x"6CE7",
			x"0000" when x"6CE8",
			x"0000" when x"6CE9",
			x"0000" when x"6CEA",
			x"0000" when x"6CEB",
			x"0000" when x"6CEC",
			x"0000" when x"6CED",
			x"0000" when x"6CEE",
			x"0000" when x"6CEF",
			x"0000" when x"6CF0",
			x"0000" when x"6CF1",
			x"0000" when x"6CF2",
			x"0000" when x"6CF3",
			x"0000" when x"6CF4",
			x"0000" when x"6CF5",
			x"0000" when x"6CF6",
			x"0000" when x"6CF7",
			x"0000" when x"6CF8",
			x"0000" when x"6CF9",
			x"0000" when x"6CFA",
			x"0000" when x"6CFB",
			x"0000" when x"6CFC",
			x"0000" when x"6CFD",
			x"0000" when x"6CFE",
			x"0000" when x"6CFF",
			x"0000" when x"6D00",
			x"0000" when x"6D01",
			x"0000" when x"6D02",
			x"0000" when x"6D03",
			x"0000" when x"6D04",
			x"0000" when x"6D05",
			x"0000" when x"6D06",
			x"0000" when x"6D07",
			x"0000" when x"6D08",
			x"0000" when x"6D09",
			x"0000" when x"6D0A",
			x"0000" when x"6D0B",
			x"0000" when x"6D0C",
			x"0000" when x"6D0D",
			x"0000" when x"6D0E",
			x"0000" when x"6D0F",
			x"0000" when x"6D10",
			x"0000" when x"6D11",
			x"0000" when x"6D12",
			x"0000" when x"6D13",
			x"0000" when x"6D14",
			x"0000" when x"6D15",
			x"0000" when x"6D16",
			x"0000" when x"6D17",
			x"0000" when x"6D18",
			x"0000" when x"6D19",
			x"0000" when x"6D1A",
			x"0000" when x"6D1B",
			x"0000" when x"6D1C",
			x"0000" when x"6D1D",
			x"0000" when x"6D1E",
			x"0000" when x"6D1F",
			x"0000" when x"6D20",
			x"0000" when x"6D21",
			x"0000" when x"6D22",
			x"0000" when x"6D23",
			x"0000" when x"6D24",
			x"0000" when x"6D25",
			x"0000" when x"6D26",
			x"0000" when x"6D27",
			x"0000" when x"6D28",
			x"0000" when x"6D29",
			x"0000" when x"6D2A",
			x"0000" when x"6D2B",
			x"0000" when x"6D2C",
			x"0000" when x"6D2D",
			x"0000" when x"6D2E",
			x"0000" when x"6D2F",
			x"0000" when x"6D30",
			x"0000" when x"6D31",
			x"0000" when x"6D32",
			x"0000" when x"6D33",
			x"0000" when x"6D34",
			x"0000" when x"6D35",
			x"0000" when x"6D36",
			x"0000" when x"6D37",
			x"0000" when x"6D38",
			x"0000" when x"6D39",
			x"0000" when x"6D3A",
			x"0000" when x"6D3B",
			x"0000" when x"6D3C",
			x"0000" when x"6D3D",
			x"0000" when x"6D3E",
			x"0000" when x"6D3F",
			x"0000" when x"6D40",
			x"0000" when x"6D41",
			x"0000" when x"6D42",
			x"0000" when x"6D43",
			x"0000" when x"6D44",
			x"0000" when x"6D45",
			x"0000" when x"6D46",
			x"0000" when x"6D47",
			x"0000" when x"6D48",
			x"0000" when x"6D49",
			x"0000" when x"6D4A",
			x"0000" when x"6D4B",
			x"0000" when x"6D4C",
			x"0000" when x"6D4D",
			x"0000" when x"6D4E",
			x"0000" when x"6D4F",
			x"0000" when x"6D50",
			x"0000" when x"6D51",
			x"0000" when x"6D52",
			x"0000" when x"6D53",
			x"0000" when x"6D54",
			x"0000" when x"6D55",
			x"0000" when x"6D56",
			x"0000" when x"6D57",
			x"0000" when x"6D58",
			x"0000" when x"6D59",
			x"0000" when x"6D5A",
			x"0000" when x"6D5B",
			x"0000" when x"6D5C",
			x"0000" when x"6D5D",
			x"0000" when x"6D5E",
			x"0000" when x"6D5F",
			x"0000" when x"6D60",
			x"0000" when x"6D61",
			x"0000" when x"6D62",
			x"0000" when x"6D63",
			x"0000" when x"6D64",
			x"0000" when x"6D65",
			x"0000" when x"6D66",
			x"0000" when x"6D67",
			x"0000" when x"6D68",
			x"0000" when x"6D69",
			x"0000" when x"6D6A",
			x"0000" when x"6D6B",
			x"0000" when x"6D6C",
			x"0000" when x"6D6D",
			x"0000" when x"6D6E",
			x"0000" when x"6D6F",
			x"0000" when x"6D70",
			x"0000" when x"6D71",
			x"0000" when x"6D72",
			x"0000" when x"6D73",
			x"0000" when x"6D74",
			x"0000" when x"6D75",
			x"0000" when x"6D76",
			x"0000" when x"6D77",
			x"0000" when x"6D78",
			x"0000" when x"6D79",
			x"0000" when x"6D7A",
			x"0000" when x"6D7B",
			x"0000" when x"6D7C",
			x"0000" when x"6D7D",
			x"0000" when x"6D7E",
			x"0000" when x"6D7F",
			x"0000" when x"6D80",
			x"0000" when x"6D81",
			x"0000" when x"6D82",
			x"0000" when x"6D83",
			x"0000" when x"6D84",
			x"0000" when x"6D85",
			x"0000" when x"6D86",
			x"0000" when x"6D87",
			x"0000" when x"6D88",
			x"0000" when x"6D89",
			x"0000" when x"6D8A",
			x"0000" when x"6D8B",
			x"0000" when x"6D8C",
			x"0000" when x"6D8D",
			x"0000" when x"6D8E",
			x"0000" when x"6D8F",
			x"0000" when x"6D90",
			x"0000" when x"6D91",
			x"0000" when x"6D92",
			x"0000" when x"6D93",
			x"0000" when x"6D94",
			x"0000" when x"6D95",
			x"0000" when x"6D96",
			x"0000" when x"6D97",
			x"0000" when x"6D98",
			x"0000" when x"6D99",
			x"0000" when x"6D9A",
			x"0000" when x"6D9B",
			x"0000" when x"6D9C",
			x"0000" when x"6D9D",
			x"0000" when x"6D9E",
			x"0000" when x"6D9F",
			x"0000" when x"6DA0",
			x"0000" when x"6DA1",
			x"0000" when x"6DA2",
			x"0000" when x"6DA3",
			x"0000" when x"6DA4",
			x"0000" when x"6DA5",
			x"0000" when x"6DA6",
			x"0000" when x"6DA7",
			x"0000" when x"6DA8",
			x"0000" when x"6DA9",
			x"0000" when x"6DAA",
			x"0000" when x"6DAB",
			x"0000" when x"6DAC",
			x"0000" when x"6DAD",
			x"0000" when x"6DAE",
			x"0000" when x"6DAF",
			x"0000" when x"6DB0",
			x"0000" when x"6DB1",
			x"0000" when x"6DB2",
			x"0000" when x"6DB3",
			x"0000" when x"6DB4",
			x"0000" when x"6DB5",
			x"0000" when x"6DB6",
			x"0000" when x"6DB7",
			x"0000" when x"6DB8",
			x"0000" when x"6DB9",
			x"0000" when x"6DBA",
			x"0000" when x"6DBB",
			x"0000" when x"6DBC",
			x"0000" when x"6DBD",
			x"0000" when x"6DBE",
			x"0000" when x"6DBF",
			x"0000" when x"6DC0",
			x"0000" when x"6DC1",
			x"0000" when x"6DC2",
			x"0000" when x"6DC3",
			x"0000" when x"6DC4",
			x"0000" when x"6DC5",
			x"0000" when x"6DC6",
			x"0000" when x"6DC7",
			x"0000" when x"6DC8",
			x"0000" when x"6DC9",
			x"0000" when x"6DCA",
			x"0000" when x"6DCB",
			x"0000" when x"6DCC",
			x"0000" when x"6DCD",
			x"0000" when x"6DCE",
			x"0000" when x"6DCF",
			x"0000" when x"6DD0",
			x"0000" when x"6DD1",
			x"0000" when x"6DD2",
			x"0000" when x"6DD3",
			x"0000" when x"6DD4",
			x"0000" when x"6DD5",
			x"0000" when x"6DD6",
			x"0000" when x"6DD7",
			x"0000" when x"6DD8",
			x"0000" when x"6DD9",
			x"0000" when x"6DDA",
			x"0000" when x"6DDB",
			x"0000" when x"6DDC",
			x"0000" when x"6DDD",
			x"0000" when x"6DDE",
			x"0000" when x"6DDF",
			x"0000" when x"6DE0",
			x"0000" when x"6DE1",
			x"0000" when x"6DE2",
			x"0000" when x"6DE3",
			x"0000" when x"6DE4",
			x"0000" when x"6DE5",
			x"0000" when x"6DE6",
			x"0000" when x"6DE7",
			x"0000" when x"6DE8",
			x"0000" when x"6DE9",
			x"0000" when x"6DEA",
			x"0000" when x"6DEB",
			x"0000" when x"6DEC",
			x"0000" when x"6DED",
			x"0000" when x"6DEE",
			x"0000" when x"6DEF",
			x"0000" when x"6DF0",
			x"0000" when x"6DF1",
			x"0000" when x"6DF2",
			x"0000" when x"6DF3",
			x"0000" when x"6DF4",
			x"0000" when x"6DF5",
			x"0000" when x"6DF6",
			x"0000" when x"6DF7",
			x"0000" when x"6DF8",
			x"0000" when x"6DF9",
			x"0000" when x"6DFA",
			x"0000" when x"6DFB",
			x"0000" when x"6DFC",
			x"0000" when x"6DFD",
			x"0000" when x"6DFE",
			x"0000" when x"6DFF",
			x"0000" when x"6E00",
			x"0000" when x"6E01",
			x"0000" when x"6E02",
			x"0000" when x"6E03",
			x"0000" when x"6E04",
			x"0000" when x"6E05",
			x"0000" when x"6E06",
			x"0000" when x"6E07",
			x"0000" when x"6E08",
			x"0000" when x"6E09",
			x"0000" when x"6E0A",
			x"0000" when x"6E0B",
			x"0000" when x"6E0C",
			x"0000" when x"6E0D",
			x"0000" when x"6E0E",
			x"0000" when x"6E0F",
			x"0000" when x"6E10",
			x"0000" when x"6E11",
			x"0000" when x"6E12",
			x"0000" when x"6E13",
			x"0000" when x"6E14",
			x"0000" when x"6E15",
			x"0000" when x"6E16",
			x"0000" when x"6E17",
			x"0000" when x"6E18",
			x"0000" when x"6E19",
			x"0000" when x"6E1A",
			x"0000" when x"6E1B",
			x"0000" when x"6E1C",
			x"0000" when x"6E1D",
			x"0000" when x"6E1E",
			x"0000" when x"6E1F",
			x"0000" when x"6E20",
			x"0000" when x"6E21",
			x"0000" when x"6E22",
			x"0000" when x"6E23",
			x"0000" when x"6E24",
			x"0000" when x"6E25",
			x"0000" when x"6E26",
			x"0000" when x"6E27",
			x"0000" when x"6E28",
			x"0000" when x"6E29",
			x"0000" when x"6E2A",
			x"0000" when x"6E2B",
			x"0000" when x"6E2C",
			x"0000" when x"6E2D",
			x"0000" when x"6E2E",
			x"0000" when x"6E2F",
			x"0000" when x"6E30",
			x"0000" when x"6E31",
			x"0000" when x"6E32",
			x"0000" when x"6E33",
			x"0000" when x"6E34",
			x"0000" when x"6E35",
			x"0000" when x"6E36",
			x"0000" when x"6E37",
			x"0000" when x"6E38",
			x"0000" when x"6E39",
			x"0000" when x"6E3A",
			x"0000" when x"6E3B",
			x"0000" when x"6E3C",
			x"0000" when x"6E3D",
			x"0000" when x"6E3E",
			x"0000" when x"6E3F",
			x"0000" when x"6E40",
			x"0000" when x"6E41",
			x"0000" when x"6E42",
			x"0000" when x"6E43",
			x"0000" when x"6E44",
			x"0000" when x"6E45",
			x"0000" when x"6E46",
			x"0000" when x"6E47",
			x"0000" when x"6E48",
			x"0000" when x"6E49",
			x"0000" when x"6E4A",
			x"0000" when x"6E4B",
			x"0000" when x"6E4C",
			x"0000" when x"6E4D",
			x"0000" when x"6E4E",
			x"0000" when x"6E4F",
			x"0000" when x"6E50",
			x"0000" when x"6E51",
			x"0000" when x"6E52",
			x"0000" when x"6E53",
			x"0000" when x"6E54",
			x"0000" when x"6E55",
			x"0000" when x"6E56",
			x"0000" when x"6E57",
			x"0000" when x"6E58",
			x"0000" when x"6E59",
			x"0000" when x"6E5A",
			x"0000" when x"6E5B",
			x"0000" when x"6E5C",
			x"0000" when x"6E5D",
			x"0000" when x"6E5E",
			x"0000" when x"6E5F",
			x"0000" when x"6E60",
			x"0000" when x"6E61",
			x"0000" when x"6E62",
			x"0000" when x"6E63",
			x"0000" when x"6E64",
			x"0000" when x"6E65",
			x"0000" when x"6E66",
			x"0000" when x"6E67",
			x"0000" when x"6E68",
			x"0000" when x"6E69",
			x"0000" when x"6E6A",
			x"0000" when x"6E6B",
			x"0000" when x"6E6C",
			x"0000" when x"6E6D",
			x"0000" when x"6E6E",
			x"0000" when x"6E6F",
			x"0000" when x"6E70",
			x"0000" when x"6E71",
			x"0000" when x"6E72",
			x"0000" when x"6E73",
			x"0000" when x"6E74",
			x"0000" when x"6E75",
			x"0000" when x"6E76",
			x"0000" when x"6E77",
			x"0000" when x"6E78",
			x"0000" when x"6E79",
			x"0000" when x"6E7A",
			x"0000" when x"6E7B",
			x"0000" when x"6E7C",
			x"0000" when x"6E7D",
			x"0000" when x"6E7E",
			x"0000" when x"6E7F",
			x"0000" when x"6E80",
			x"0000" when x"6E81",
			x"0000" when x"6E82",
			x"0000" when x"6E83",
			x"0000" when x"6E84",
			x"0000" when x"6E85",
			x"0000" when x"6E86",
			x"0000" when x"6E87",
			x"0000" when x"6E88",
			x"0000" when x"6E89",
			x"0000" when x"6E8A",
			x"0000" when x"6E8B",
			x"0000" when x"6E8C",
			x"0000" when x"6E8D",
			x"0000" when x"6E8E",
			x"0000" when x"6E8F",
			x"0000" when x"6E90",
			x"0000" when x"6E91",
			x"0000" when x"6E92",
			x"0000" when x"6E93",
			x"0000" when x"6E94",
			x"0000" when x"6E95",
			x"0000" when x"6E96",
			x"0000" when x"6E97",
			x"0000" when x"6E98",
			x"0000" when x"6E99",
			x"0000" when x"6E9A",
			x"0000" when x"6E9B",
			x"0000" when x"6E9C",
			x"0000" when x"6E9D",
			x"0000" when x"6E9E",
			x"0000" when x"6E9F",
			x"0000" when x"6EA0",
			x"0000" when x"6EA1",
			x"0000" when x"6EA2",
			x"0000" when x"6EA3",
			x"0000" when x"6EA4",
			x"0000" when x"6EA5",
			x"0000" when x"6EA6",
			x"0000" when x"6EA7",
			x"0000" when x"6EA8",
			x"0000" when x"6EA9",
			x"0000" when x"6EAA",
			x"0000" when x"6EAB",
			x"0000" when x"6EAC",
			x"0000" when x"6EAD",
			x"0000" when x"6EAE",
			x"0000" when x"6EAF",
			x"0000" when x"6EB0",
			x"0000" when x"6EB1",
			x"0000" when x"6EB2",
			x"0000" when x"6EB3",
			x"0000" when x"6EB4",
			x"0000" when x"6EB5",
			x"0000" when x"6EB6",
			x"0000" when x"6EB7",
			x"0000" when x"6EB8",
			x"0000" when x"6EB9",
			x"0000" when x"6EBA",
			x"0000" when x"6EBB",
			x"0000" when x"6EBC",
			x"0000" when x"6EBD",
			x"0000" when x"6EBE",
			x"0000" when x"6EBF",
			x"0000" when x"6EC0",
			x"0000" when x"6EC1",
			x"0000" when x"6EC2",
			x"0000" when x"6EC3",
			x"0000" when x"6EC4",
			x"0000" when x"6EC5",
			x"0000" when x"6EC6",
			x"0000" when x"6EC7",
			x"0000" when x"6EC8",
			x"0000" when x"6EC9",
			x"0000" when x"6ECA",
			x"0000" when x"6ECB",
			x"0000" when x"6ECC",
			x"0000" when x"6ECD",
			x"0000" when x"6ECE",
			x"0000" when x"6ECF",
			x"0000" when x"6ED0",
			x"0000" when x"6ED1",
			x"0000" when x"6ED2",
			x"0000" when x"6ED3",
			x"0000" when x"6ED4",
			x"0000" when x"6ED5",
			x"0000" when x"6ED6",
			x"0000" when x"6ED7",
			x"0000" when x"6ED8",
			x"0000" when x"6ED9",
			x"0000" when x"6EDA",
			x"0000" when x"6EDB",
			x"0000" when x"6EDC",
			x"0000" when x"6EDD",
			x"0000" when x"6EDE",
			x"0000" when x"6EDF",
			x"0000" when x"6EE0",
			x"0000" when x"6EE1",
			x"0000" when x"6EE2",
			x"0000" when x"6EE3",
			x"0000" when x"6EE4",
			x"0000" when x"6EE5",
			x"0000" when x"6EE6",
			x"0000" when x"6EE7",
			x"0000" when x"6EE8",
			x"0000" when x"6EE9",
			x"0000" when x"6EEA",
			x"0000" when x"6EEB",
			x"0000" when x"6EEC",
			x"0000" when x"6EED",
			x"0000" when x"6EEE",
			x"0000" when x"6EEF",
			x"0000" when x"6EF0",
			x"0000" when x"6EF1",
			x"0000" when x"6EF2",
			x"0000" when x"6EF3",
			x"0000" when x"6EF4",
			x"0000" when x"6EF5",
			x"0000" when x"6EF6",
			x"0000" when x"6EF7",
			x"0000" when x"6EF8",
			x"0000" when x"6EF9",
			x"0000" when x"6EFA",
			x"0000" when x"6EFB",
			x"0000" when x"6EFC",
			x"0000" when x"6EFD",
			x"0000" when x"6EFE",
			x"0000" when x"6EFF",
			x"0000" when x"6F00",
			x"0000" when x"6F01",
			x"0000" when x"6F02",
			x"0000" when x"6F03",
			x"0000" when x"6F04",
			x"0000" when x"6F05",
			x"0000" when x"6F06",
			x"0000" when x"6F07",
			x"0000" when x"6F08",
			x"0000" when x"6F09",
			x"0000" when x"6F0A",
			x"0000" when x"6F0B",
			x"0000" when x"6F0C",
			x"0000" when x"6F0D",
			x"0000" when x"6F0E",
			x"0000" when x"6F0F",
			x"0000" when x"6F10",
			x"0000" when x"6F11",
			x"0000" when x"6F12",
			x"0000" when x"6F13",
			x"0000" when x"6F14",
			x"0000" when x"6F15",
			x"0000" when x"6F16",
			x"0000" when x"6F17",
			x"0000" when x"6F18",
			x"0000" when x"6F19",
			x"0000" when x"6F1A",
			x"0000" when x"6F1B",
			x"0000" when x"6F1C",
			x"0000" when x"6F1D",
			x"0000" when x"6F1E",
			x"0000" when x"6F1F",
			x"0000" when x"6F20",
			x"0000" when x"6F21",
			x"0000" when x"6F22",
			x"0000" when x"6F23",
			x"0000" when x"6F24",
			x"0000" when x"6F25",
			x"0000" when x"6F26",
			x"0000" when x"6F27",
			x"0000" when x"6F28",
			x"0000" when x"6F29",
			x"0000" when x"6F2A",
			x"0000" when x"6F2B",
			x"0000" when x"6F2C",
			x"0000" when x"6F2D",
			x"0000" when x"6F2E",
			x"0000" when x"6F2F",
			x"0000" when x"6F30",
			x"0000" when x"6F31",
			x"0000" when x"6F32",
			x"0000" when x"6F33",
			x"0000" when x"6F34",
			x"0000" when x"6F35",
			x"0000" when x"6F36",
			x"0000" when x"6F37",
			x"0000" when x"6F38",
			x"0000" when x"6F39",
			x"0000" when x"6F3A",
			x"0000" when x"6F3B",
			x"0000" when x"6F3C",
			x"0000" when x"6F3D",
			x"0000" when x"6F3E",
			x"0000" when x"6F3F",
			x"0000" when x"6F40",
			x"0000" when x"6F41",
			x"0000" when x"6F42",
			x"0000" when x"6F43",
			x"0000" when x"6F44",
			x"0000" when x"6F45",
			x"0000" when x"6F46",
			x"0000" when x"6F47",
			x"0000" when x"6F48",
			x"0000" when x"6F49",
			x"0000" when x"6F4A",
			x"0000" when x"6F4B",
			x"0000" when x"6F4C",
			x"0000" when x"6F4D",
			x"0000" when x"6F4E",
			x"0000" when x"6F4F",
			x"0000" when x"6F50",
			x"0000" when x"6F51",
			x"0000" when x"6F52",
			x"0000" when x"6F53",
			x"0000" when x"6F54",
			x"0000" when x"6F55",
			x"0000" when x"6F56",
			x"0000" when x"6F57",
			x"0000" when x"6F58",
			x"0000" when x"6F59",
			x"0000" when x"6F5A",
			x"0000" when x"6F5B",
			x"0000" when x"6F5C",
			x"0000" when x"6F5D",
			x"0000" when x"6F5E",
			x"0000" when x"6F5F",
			x"0000" when x"6F60",
			x"0000" when x"6F61",
			x"0000" when x"6F62",
			x"0000" when x"6F63",
			x"0000" when x"6F64",
			x"0000" when x"6F65",
			x"0000" when x"6F66",
			x"0000" when x"6F67",
			x"0000" when x"6F68",
			x"0000" when x"6F69",
			x"0000" when x"6F6A",
			x"0000" when x"6F6B",
			x"0000" when x"6F6C",
			x"0000" when x"6F6D",
			x"0000" when x"6F6E",
			x"0000" when x"6F6F",
			x"0000" when x"6F70",
			x"0000" when x"6F71",
			x"0000" when x"6F72",
			x"0000" when x"6F73",
			x"0000" when x"6F74",
			x"0000" when x"6F75",
			x"0000" when x"6F76",
			x"0000" when x"6F77",
			x"0000" when x"6F78",
			x"0000" when x"6F79",
			x"0000" when x"6F7A",
			x"0000" when x"6F7B",
			x"0000" when x"6F7C",
			x"0000" when x"6F7D",
			x"0000" when x"6F7E",
			x"0000" when x"6F7F",
			x"0000" when x"6F80",
			x"0000" when x"6F81",
			x"0000" when x"6F82",
			x"0000" when x"6F83",
			x"0000" when x"6F84",
			x"0000" when x"6F85",
			x"0000" when x"6F86",
			x"0000" when x"6F87",
			x"0000" when x"6F88",
			x"0000" when x"6F89",
			x"0000" when x"6F8A",
			x"0000" when x"6F8B",
			x"0000" when x"6F8C",
			x"0000" when x"6F8D",
			x"0000" when x"6F8E",
			x"0000" when x"6F8F",
			x"0000" when x"6F90",
			x"0000" when x"6F91",
			x"0000" when x"6F92",
			x"0000" when x"6F93",
			x"0000" when x"6F94",
			x"0000" when x"6F95",
			x"0000" when x"6F96",
			x"0000" when x"6F97",
			x"0000" when x"6F98",
			x"0000" when x"6F99",
			x"0000" when x"6F9A",
			x"0000" when x"6F9B",
			x"0000" when x"6F9C",
			x"0000" when x"6F9D",
			x"0000" when x"6F9E",
			x"0000" when x"6F9F",
			x"0000" when x"6FA0",
			x"0000" when x"6FA1",
			x"0000" when x"6FA2",
			x"0000" when x"6FA3",
			x"0000" when x"6FA4",
			x"0000" when x"6FA5",
			x"0000" when x"6FA6",
			x"0000" when x"6FA7",
			x"0000" when x"6FA8",
			x"0000" when x"6FA9",
			x"0000" when x"6FAA",
			x"0000" when x"6FAB",
			x"0000" when x"6FAC",
			x"0000" when x"6FAD",
			x"0000" when x"6FAE",
			x"0000" when x"6FAF",
			x"0000" when x"6FB0",
			x"0000" when x"6FB1",
			x"0000" when x"6FB2",
			x"0000" when x"6FB3",
			x"0000" when x"6FB4",
			x"0000" when x"6FB5",
			x"0000" when x"6FB6",
			x"0000" when x"6FB7",
			x"0000" when x"6FB8",
			x"0000" when x"6FB9",
			x"0000" when x"6FBA",
			x"0000" when x"6FBB",
			x"0000" when x"6FBC",
			x"0000" when x"6FBD",
			x"0000" when x"6FBE",
			x"0000" when x"6FBF",
			x"0000" when x"6FC0",
			x"0000" when x"6FC1",
			x"0000" when x"6FC2",
			x"0000" when x"6FC3",
			x"0000" when x"6FC4",
			x"0000" when x"6FC5",
			x"0000" when x"6FC6",
			x"0000" when x"6FC7",
			x"0000" when x"6FC8",
			x"0000" when x"6FC9",
			x"0000" when x"6FCA",
			x"0000" when x"6FCB",
			x"0000" when x"6FCC",
			x"0000" when x"6FCD",
			x"0000" when x"6FCE",
			x"0000" when x"6FCF",
			x"0000" when x"6FD0",
			x"0000" when x"6FD1",
			x"0000" when x"6FD2",
			x"0000" when x"6FD3",
			x"0000" when x"6FD4",
			x"0000" when x"6FD5",
			x"0000" when x"6FD6",
			x"0000" when x"6FD7",
			x"0000" when x"6FD8",
			x"0000" when x"6FD9",
			x"0000" when x"6FDA",
			x"0000" when x"6FDB",
			x"0000" when x"6FDC",
			x"0000" when x"6FDD",
			x"0000" when x"6FDE",
			x"0000" when x"6FDF",
			x"0000" when x"6FE0",
			x"0000" when x"6FE1",
			x"0000" when x"6FE2",
			x"0000" when x"6FE3",
			x"0000" when x"6FE4",
			x"0000" when x"6FE5",
			x"0000" when x"6FE6",
			x"0000" when x"6FE7",
			x"0000" when x"6FE8",
			x"0000" when x"6FE9",
			x"0000" when x"6FEA",
			x"0000" when x"6FEB",
			x"0000" when x"6FEC",
			x"0000" when x"6FED",
			x"0000" when x"6FEE",
			x"0000" when x"6FEF",
			x"0000" when x"6FF0",
			x"0000" when x"6FF1",
			x"0000" when x"6FF2",
			x"0000" when x"6FF3",
			x"0000" when x"6FF4",
			x"0000" when x"6FF5",
			x"0000" when x"6FF6",
			x"0000" when x"6FF7",
			x"0000" when x"6FF8",
			x"0000" when x"6FF9",
			x"0000" when x"6FFA",
			x"0000" when x"6FFB",
			x"0000" when x"6FFC",
			x"0000" when x"6FFD",
			x"0000" when x"6FFE",
			x"0000" when x"6FFF",
			x"0000" when x"7000",
			x"0000" when x"7001",
			x"0000" when x"7002",
			x"0000" when x"7003",
			x"0000" when x"7004",
			x"0000" when x"7005",
			x"0000" when x"7006",
			x"0000" when x"7007",
			x"0000" when x"7008",
			x"0000" when x"7009",
			x"0000" when x"700A",
			x"0000" when x"700B",
			x"0000" when x"700C",
			x"0000" when x"700D",
			x"0000" when x"700E",
			x"0000" when x"700F",
			x"0000" when x"7010",
			x"0000" when x"7011",
			x"0000" when x"7012",
			x"0000" when x"7013",
			x"0000" when x"7014",
			x"0000" when x"7015",
			x"0000" when x"7016",
			x"0000" when x"7017",
			x"0000" when x"7018",
			x"0000" when x"7019",
			x"0000" when x"701A",
			x"0000" when x"701B",
			x"0000" when x"701C",
			x"0000" when x"701D",
			x"0000" when x"701E",
			x"0000" when x"701F",
			x"0000" when x"7020",
			x"0000" when x"7021",
			x"0000" when x"7022",
			x"0000" when x"7023",
			x"0000" when x"7024",
			x"0000" when x"7025",
			x"0000" when x"7026",
			x"0000" when x"7027",
			x"0000" when x"7028",
			x"0000" when x"7029",
			x"0000" when x"702A",
			x"0000" when x"702B",
			x"0000" when x"702C",
			x"0000" when x"702D",
			x"0000" when x"702E",
			x"0000" when x"702F",
			x"0000" when x"7030",
			x"0000" when x"7031",
			x"0000" when x"7032",
			x"0000" when x"7033",
			x"0000" when x"7034",
			x"0000" when x"7035",
			x"0000" when x"7036",
			x"0000" when x"7037",
			x"0000" when x"7038",
			x"0000" when x"7039",
			x"0000" when x"703A",
			x"0000" when x"703B",
			x"0000" when x"703C",
			x"0000" when x"703D",
			x"0000" when x"703E",
			x"0000" when x"703F",
			x"0000" when x"7040",
			x"0000" when x"7041",
			x"0000" when x"7042",
			x"0000" when x"7043",
			x"0000" when x"7044",
			x"0000" when x"7045",
			x"0000" when x"7046",
			x"0000" when x"7047",
			x"0000" when x"7048",
			x"0000" when x"7049",
			x"0000" when x"704A",
			x"0000" when x"704B",
			x"0000" when x"704C",
			x"0000" when x"704D",
			x"0000" when x"704E",
			x"0000" when x"704F",
			x"0000" when x"7050",
			x"0000" when x"7051",
			x"0000" when x"7052",
			x"0000" when x"7053",
			x"0000" when x"7054",
			x"0000" when x"7055",
			x"0000" when x"7056",
			x"0000" when x"7057",
			x"0000" when x"7058",
			x"0000" when x"7059",
			x"0000" when x"705A",
			x"0000" when x"705B",
			x"0000" when x"705C",
			x"0000" when x"705D",
			x"0000" when x"705E",
			x"0000" when x"705F",
			x"0000" when x"7060",
			x"0000" when x"7061",
			x"0000" when x"7062",
			x"0000" when x"7063",
			x"0000" when x"7064",
			x"0000" when x"7065",
			x"0000" when x"7066",
			x"0000" when x"7067",
			x"0000" when x"7068",
			x"0000" when x"7069",
			x"0000" when x"706A",
			x"0000" when x"706B",
			x"0000" when x"706C",
			x"0000" when x"706D",
			x"0000" when x"706E",
			x"0000" when x"706F",
			x"0000" when x"7070",
			x"0000" when x"7071",
			x"0000" when x"7072",
			x"0000" when x"7073",
			x"0000" when x"7074",
			x"0000" when x"7075",
			x"0000" when x"7076",
			x"0000" when x"7077",
			x"0000" when x"7078",
			x"0000" when x"7079",
			x"0000" when x"707A",
			x"0000" when x"707B",
			x"0000" when x"707C",
			x"0000" when x"707D",
			x"0000" when x"707E",
			x"0000" when x"707F",
			x"0000" when x"7080",
			x"0000" when x"7081",
			x"0000" when x"7082",
			x"0000" when x"7083",
			x"0000" when x"7084",
			x"0000" when x"7085",
			x"0000" when x"7086",
			x"0000" when x"7087",
			x"0000" when x"7088",
			x"0000" when x"7089",
			x"0000" when x"708A",
			x"0000" when x"708B",
			x"0000" when x"708C",
			x"0000" when x"708D",
			x"0000" when x"708E",
			x"0000" when x"708F",
			x"0000" when x"7090",
			x"0000" when x"7091",
			x"0000" when x"7092",
			x"0000" when x"7093",
			x"0000" when x"7094",
			x"0000" when x"7095",
			x"0000" when x"7096",
			x"0000" when x"7097",
			x"0000" when x"7098",
			x"0000" when x"7099",
			x"0000" when x"709A",
			x"0000" when x"709B",
			x"0000" when x"709C",
			x"0000" when x"709D",
			x"0000" when x"709E",
			x"0000" when x"709F",
			x"0000" when x"70A0",
			x"0000" when x"70A1",
			x"0000" when x"70A2",
			x"0000" when x"70A3",
			x"0000" when x"70A4",
			x"0000" when x"70A5",
			x"0000" when x"70A6",
			x"0000" when x"70A7",
			x"0000" when x"70A8",
			x"0000" when x"70A9",
			x"0000" when x"70AA",
			x"0000" when x"70AB",
			x"0000" when x"70AC",
			x"0000" when x"70AD",
			x"0000" when x"70AE",
			x"0000" when x"70AF",
			x"0000" when x"70B0",
			x"0000" when x"70B1",
			x"0000" when x"70B2",
			x"0000" when x"70B3",
			x"0000" when x"70B4",
			x"0000" when x"70B5",
			x"0000" when x"70B6",
			x"0000" when x"70B7",
			x"0000" when x"70B8",
			x"0000" when x"70B9",
			x"0000" when x"70BA",
			x"0000" when x"70BB",
			x"0000" when x"70BC",
			x"0000" when x"70BD",
			x"0000" when x"70BE",
			x"0000" when x"70BF",
			x"0000" when x"70C0",
			x"0000" when x"70C1",
			x"0000" when x"70C2",
			x"0000" when x"70C3",
			x"0000" when x"70C4",
			x"0000" when x"70C5",
			x"0000" when x"70C6",
			x"0000" when x"70C7",
			x"0000" when x"70C8",
			x"0000" when x"70C9",
			x"0000" when x"70CA",
			x"0000" when x"70CB",
			x"0000" when x"70CC",
			x"0000" when x"70CD",
			x"0000" when x"70CE",
			x"0000" when x"70CF",
			x"0000" when x"70D0",
			x"0000" when x"70D1",
			x"0000" when x"70D2",
			x"0000" when x"70D3",
			x"0000" when x"70D4",
			x"0000" when x"70D5",
			x"0000" when x"70D6",
			x"0000" when x"70D7",
			x"0000" when x"70D8",
			x"0000" when x"70D9",
			x"0000" when x"70DA",
			x"0000" when x"70DB",
			x"0000" when x"70DC",
			x"0000" when x"70DD",
			x"0000" when x"70DE",
			x"0000" when x"70DF",
			x"0000" when x"70E0",
			x"0000" when x"70E1",
			x"0000" when x"70E2",
			x"0000" when x"70E3",
			x"0000" when x"70E4",
			x"0000" when x"70E5",
			x"0000" when x"70E6",
			x"0000" when x"70E7",
			x"0000" when x"70E8",
			x"0000" when x"70E9",
			x"0000" when x"70EA",
			x"0000" when x"70EB",
			x"0000" when x"70EC",
			x"0000" when x"70ED",
			x"0000" when x"70EE",
			x"0000" when x"70EF",
			x"0000" when x"70F0",
			x"0000" when x"70F1",
			x"0000" when x"70F2",
			x"0000" when x"70F3",
			x"0000" when x"70F4",
			x"0000" when x"70F5",
			x"0000" when x"70F6",
			x"0000" when x"70F7",
			x"0000" when x"70F8",
			x"0000" when x"70F9",
			x"0000" when x"70FA",
			x"0000" when x"70FB",
			x"0000" when x"70FC",
			x"0000" when x"70FD",
			x"0000" when x"70FE",
			x"0000" when x"70FF",
			x"0000" when x"7100",
			x"0000" when x"7101",
			x"0000" when x"7102",
			x"0000" when x"7103",
			x"0000" when x"7104",
			x"0000" when x"7105",
			x"0000" when x"7106",
			x"0000" when x"7107",
			x"0000" when x"7108",
			x"0000" when x"7109",
			x"0000" when x"710A",
			x"0000" when x"710B",
			x"0000" when x"710C",
			x"0000" when x"710D",
			x"0000" when x"710E",
			x"0000" when x"710F",
			x"0000" when x"7110",
			x"0000" when x"7111",
			x"0000" when x"7112",
			x"0000" when x"7113",
			x"0000" when x"7114",
			x"0000" when x"7115",
			x"0000" when x"7116",
			x"0000" when x"7117",
			x"0000" when x"7118",
			x"0000" when x"7119",
			x"0000" when x"711A",
			x"0000" when x"711B",
			x"0000" when x"711C",
			x"0000" when x"711D",
			x"0000" when x"711E",
			x"0000" when x"711F",
			x"0000" when x"7120",
			x"0000" when x"7121",
			x"0000" when x"7122",
			x"0000" when x"7123",
			x"0000" when x"7124",
			x"0000" when x"7125",
			x"0000" when x"7126",
			x"0000" when x"7127",
			x"0000" when x"7128",
			x"0000" when x"7129",
			x"0000" when x"712A",
			x"0000" when x"712B",
			x"0000" when x"712C",
			x"0000" when x"712D",
			x"0000" when x"712E",
			x"0000" when x"712F",
			x"0000" when x"7130",
			x"0000" when x"7131",
			x"0000" when x"7132",
			x"0000" when x"7133",
			x"0000" when x"7134",
			x"0000" when x"7135",
			x"0000" when x"7136",
			x"0000" when x"7137",
			x"0000" when x"7138",
			x"0000" when x"7139",
			x"0000" when x"713A",
			x"0000" when x"713B",
			x"0000" when x"713C",
			x"0000" when x"713D",
			x"0000" when x"713E",
			x"0000" when x"713F",
			x"0000" when x"7140",
			x"0000" when x"7141",
			x"0000" when x"7142",
			x"0000" when x"7143",
			x"0000" when x"7144",
			x"0000" when x"7145",
			x"0000" when x"7146",
			x"0000" when x"7147",
			x"0000" when x"7148",
			x"0000" when x"7149",
			x"0000" when x"714A",
			x"0000" when x"714B",
			x"0000" when x"714C",
			x"0000" when x"714D",
			x"0000" when x"714E",
			x"0000" when x"714F",
			x"0000" when x"7150",
			x"0000" when x"7151",
			x"0000" when x"7152",
			x"0000" when x"7153",
			x"0000" when x"7154",
			x"0000" when x"7155",
			x"0000" when x"7156",
			x"0000" when x"7157",
			x"0000" when x"7158",
			x"0000" when x"7159",
			x"0000" when x"715A",
			x"0000" when x"715B",
			x"0000" when x"715C",
			x"0000" when x"715D",
			x"0000" when x"715E",
			x"0000" when x"715F",
			x"0000" when x"7160",
			x"0000" when x"7161",
			x"0000" when x"7162",
			x"0000" when x"7163",
			x"0000" when x"7164",
			x"0000" when x"7165",
			x"0000" when x"7166",
			x"0000" when x"7167",
			x"0000" when x"7168",
			x"0000" when x"7169",
			x"0000" when x"716A",
			x"0000" when x"716B",
			x"0000" when x"716C",
			x"0000" when x"716D",
			x"0000" when x"716E",
			x"0000" when x"716F",
			x"0000" when x"7170",
			x"0000" when x"7171",
			x"0000" when x"7172",
			x"0000" when x"7173",
			x"0000" when x"7174",
			x"0000" when x"7175",
			x"0000" when x"7176",
			x"0000" when x"7177",
			x"0000" when x"7178",
			x"0000" when x"7179",
			x"0000" when x"717A",
			x"0000" when x"717B",
			x"0000" when x"717C",
			x"0000" when x"717D",
			x"0000" when x"717E",
			x"0000" when x"717F",
			x"0000" when x"7180",
			x"0000" when x"7181",
			x"0000" when x"7182",
			x"0000" when x"7183",
			x"0000" when x"7184",
			x"0000" when x"7185",
			x"0000" when x"7186",
			x"0000" when x"7187",
			x"0000" when x"7188",
			x"0000" when x"7189",
			x"0000" when x"718A",
			x"0000" when x"718B",
			x"0000" when x"718C",
			x"0000" when x"718D",
			x"0000" when x"718E",
			x"0000" when x"718F",
			x"0000" when x"7190",
			x"0000" when x"7191",
			x"0000" when x"7192",
			x"0000" when x"7193",
			x"0000" when x"7194",
			x"0000" when x"7195",
			x"0000" when x"7196",
			x"0000" when x"7197",
			x"0000" when x"7198",
			x"0000" when x"7199",
			x"0000" when x"719A",
			x"0000" when x"719B",
			x"0000" when x"719C",
			x"0000" when x"719D",
			x"0000" when x"719E",
			x"0000" when x"719F",
			x"0000" when x"71A0",
			x"0000" when x"71A1",
			x"0000" when x"71A2",
			x"0000" when x"71A3",
			x"0000" when x"71A4",
			x"0000" when x"71A5",
			x"0000" when x"71A6",
			x"0000" when x"71A7",
			x"0000" when x"71A8",
			x"0000" when x"71A9",
			x"0000" when x"71AA",
			x"0000" when x"71AB",
			x"0000" when x"71AC",
			x"0000" when x"71AD",
			x"0000" when x"71AE",
			x"0000" when x"71AF",
			x"0000" when x"71B0",
			x"0000" when x"71B1",
			x"0000" when x"71B2",
			x"0000" when x"71B3",
			x"0000" when x"71B4",
			x"0000" when x"71B5",
			x"0000" when x"71B6",
			x"0000" when x"71B7",
			x"0000" when x"71B8",
			x"0000" when x"71B9",
			x"0000" when x"71BA",
			x"0000" when x"71BB",
			x"0000" when x"71BC",
			x"0000" when x"71BD",
			x"0000" when x"71BE",
			x"0000" when x"71BF",
			x"0000" when x"71C0",
			x"0000" when x"71C1",
			x"0000" when x"71C2",
			x"0000" when x"71C3",
			x"0000" when x"71C4",
			x"0000" when x"71C5",
			x"0000" when x"71C6",
			x"0000" when x"71C7",
			x"0000" when x"71C8",
			x"0000" when x"71C9",
			x"0000" when x"71CA",
			x"0000" when x"71CB",
			x"0000" when x"71CC",
			x"0000" when x"71CD",
			x"0000" when x"71CE",
			x"0000" when x"71CF",
			x"0000" when x"71D0",
			x"0000" when x"71D1",
			x"0000" when x"71D2",
			x"0000" when x"71D3",
			x"0000" when x"71D4",
			x"0000" when x"71D5",
			x"0000" when x"71D6",
			x"0000" when x"71D7",
			x"0000" when x"71D8",
			x"0000" when x"71D9",
			x"0000" when x"71DA",
			x"0000" when x"71DB",
			x"0000" when x"71DC",
			x"0000" when x"71DD",
			x"0000" when x"71DE",
			x"0000" when x"71DF",
			x"0000" when x"71E0",
			x"0000" when x"71E1",
			x"0000" when x"71E2",
			x"0000" when x"71E3",
			x"0000" when x"71E4",
			x"0000" when x"71E5",
			x"0000" when x"71E6",
			x"0000" when x"71E7",
			x"0000" when x"71E8",
			x"0000" when x"71E9",
			x"0000" when x"71EA",
			x"0000" when x"71EB",
			x"0000" when x"71EC",
			x"0000" when x"71ED",
			x"0000" when x"71EE",
			x"0000" when x"71EF",
			x"0000" when x"71F0",
			x"0000" when x"71F1",
			x"0000" when x"71F2",
			x"0000" when x"71F3",
			x"0000" when x"71F4",
			x"0000" when x"71F5",
			x"0000" when x"71F6",
			x"0000" when x"71F7",
			x"0000" when x"71F8",
			x"0000" when x"71F9",
			x"0000" when x"71FA",
			x"0000" when x"71FB",
			x"0000" when x"71FC",
			x"0000" when x"71FD",
			x"0000" when x"71FE",
			x"0000" when x"71FF",
			x"0000" when x"7200",
			x"0000" when x"7201",
			x"0000" when x"7202",
			x"0000" when x"7203",
			x"0000" when x"7204",
			x"0000" when x"7205",
			x"0000" when x"7206",
			x"0000" when x"7207",
			x"0000" when x"7208",
			x"0000" when x"7209",
			x"0000" when x"720A",
			x"0000" when x"720B",
			x"0000" when x"720C",
			x"0000" when x"720D",
			x"0000" when x"720E",
			x"0000" when x"720F",
			x"0000" when x"7210",
			x"0000" when x"7211",
			x"0000" when x"7212",
			x"0000" when x"7213",
			x"0000" when x"7214",
			x"0000" when x"7215",
			x"0000" when x"7216",
			x"0000" when x"7217",
			x"0000" when x"7218",
			x"0000" when x"7219",
			x"0000" when x"721A",
			x"0000" when x"721B",
			x"0000" when x"721C",
			x"0000" when x"721D",
			x"0000" when x"721E",
			x"0000" when x"721F",
			x"0000" when x"7220",
			x"0000" when x"7221",
			x"0000" when x"7222",
			x"0000" when x"7223",
			x"0000" when x"7224",
			x"0000" when x"7225",
			x"0000" when x"7226",
			x"0000" when x"7227",
			x"0000" when x"7228",
			x"0000" when x"7229",
			x"0000" when x"722A",
			x"0000" when x"722B",
			x"0000" when x"722C",
			x"0000" when x"722D",
			x"0000" when x"722E",
			x"0000" when x"722F",
			x"0000" when x"7230",
			x"0000" when x"7231",
			x"0000" when x"7232",
			x"0000" when x"7233",
			x"0000" when x"7234",
			x"0000" when x"7235",
			x"0000" when x"7236",
			x"0000" when x"7237",
			x"0000" when x"7238",
			x"0000" when x"7239",
			x"0000" when x"723A",
			x"0000" when x"723B",
			x"0000" when x"723C",
			x"0000" when x"723D",
			x"0000" when x"723E",
			x"0000" when x"723F",
			x"0000" when x"7240",
			x"0000" when x"7241",
			x"0000" when x"7242",
			x"0000" when x"7243",
			x"0000" when x"7244",
			x"0000" when x"7245",
			x"0000" when x"7246",
			x"0000" when x"7247",
			x"0000" when x"7248",
			x"0000" when x"7249",
			x"0000" when x"724A",
			x"0000" when x"724B",
			x"0000" when x"724C",
			x"0000" when x"724D",
			x"0000" when x"724E",
			x"0000" when x"724F",
			x"0000" when x"7250",
			x"0000" when x"7251",
			x"0000" when x"7252",
			x"0000" when x"7253",
			x"0000" when x"7254",
			x"0000" when x"7255",
			x"0000" when x"7256",
			x"0000" when x"7257",
			x"0000" when x"7258",
			x"0000" when x"7259",
			x"0000" when x"725A",
			x"0000" when x"725B",
			x"0000" when x"725C",
			x"0000" when x"725D",
			x"0000" when x"725E",
			x"0000" when x"725F",
			x"0000" when x"7260",
			x"0000" when x"7261",
			x"0000" when x"7262",
			x"0000" when x"7263",
			x"0000" when x"7264",
			x"0000" when x"7265",
			x"0000" when x"7266",
			x"0000" when x"7267",
			x"0000" when x"7268",
			x"0000" when x"7269",
			x"0000" when x"726A",
			x"0000" when x"726B",
			x"0000" when x"726C",
			x"0000" when x"726D",
			x"0000" when x"726E",
			x"0000" when x"726F",
			x"0000" when x"7270",
			x"0000" when x"7271",
			x"0000" when x"7272",
			x"0000" when x"7273",
			x"0000" when x"7274",
			x"0000" when x"7275",
			x"0000" when x"7276",
			x"0000" when x"7277",
			x"0000" when x"7278",
			x"0000" when x"7279",
			x"0000" when x"727A",
			x"0000" when x"727B",
			x"0000" when x"727C",
			x"0000" when x"727D",
			x"0000" when x"727E",
			x"0000" when x"727F",
			x"0000" when x"7280",
			x"0000" when x"7281",
			x"0000" when x"7282",
			x"0000" when x"7283",
			x"0000" when x"7284",
			x"0000" when x"7285",
			x"0000" when x"7286",
			x"0000" when x"7287",
			x"0000" when x"7288",
			x"0000" when x"7289",
			x"0000" when x"728A",
			x"0000" when x"728B",
			x"0000" when x"728C",
			x"0000" when x"728D",
			x"0000" when x"728E",
			x"0000" when x"728F",
			x"0000" when x"7290",
			x"0000" when x"7291",
			x"0000" when x"7292",
			x"0000" when x"7293",
			x"0000" when x"7294",
			x"0000" when x"7295",
			x"0000" when x"7296",
			x"0000" when x"7297",
			x"0000" when x"7298",
			x"0000" when x"7299",
			x"0000" when x"729A",
			x"0000" when x"729B",
			x"0000" when x"729C",
			x"0000" when x"729D",
			x"0000" when x"729E",
			x"0000" when x"729F",
			x"0000" when x"72A0",
			x"0000" when x"72A1",
			x"0000" when x"72A2",
			x"0000" when x"72A3",
			x"0000" when x"72A4",
			x"0000" when x"72A5",
			x"0000" when x"72A6",
			x"0000" when x"72A7",
			x"0000" when x"72A8",
			x"0000" when x"72A9",
			x"0000" when x"72AA",
			x"0000" when x"72AB",
			x"0000" when x"72AC",
			x"0000" when x"72AD",
			x"0000" when x"72AE",
			x"0000" when x"72AF",
			x"0000" when x"72B0",
			x"0000" when x"72B1",
			x"0000" when x"72B2",
			x"0000" when x"72B3",
			x"0000" when x"72B4",
			x"0000" when x"72B5",
			x"0000" when x"72B6",
			x"0000" when x"72B7",
			x"0000" when x"72B8",
			x"0000" when x"72B9",
			x"0000" when x"72BA",
			x"0000" when x"72BB",
			x"0000" when x"72BC",
			x"0000" when x"72BD",
			x"0000" when x"72BE",
			x"0000" when x"72BF",
			x"0000" when x"72C0",
			x"0000" when x"72C1",
			x"0000" when x"72C2",
			x"0000" when x"72C3",
			x"0000" when x"72C4",
			x"0000" when x"72C5",
			x"0000" when x"72C6",
			x"0000" when x"72C7",
			x"0000" when x"72C8",
			x"0000" when x"72C9",
			x"0000" when x"72CA",
			x"0000" when x"72CB",
			x"0000" when x"72CC",
			x"0000" when x"72CD",
			x"0000" when x"72CE",
			x"0000" when x"72CF",
			x"0000" when x"72D0",
			x"0000" when x"72D1",
			x"0000" when x"72D2",
			x"0000" when x"72D3",
			x"0000" when x"72D4",
			x"0000" when x"72D5",
			x"0000" when x"72D6",
			x"0000" when x"72D7",
			x"0000" when x"72D8",
			x"0000" when x"72D9",
			x"0000" when x"72DA",
			x"0000" when x"72DB",
			x"0000" when x"72DC",
			x"0000" when x"72DD",
			x"0000" when x"72DE",
			x"0000" when x"72DF",
			x"0000" when x"72E0",
			x"0000" when x"72E1",
			x"0000" when x"72E2",
			x"0000" when x"72E3",
			x"0000" when x"72E4",
			x"0000" when x"72E5",
			x"0000" when x"72E6",
			x"0000" when x"72E7",
			x"0000" when x"72E8",
			x"0000" when x"72E9",
			x"0000" when x"72EA",
			x"0000" when x"72EB",
			x"0000" when x"72EC",
			x"0000" when x"72ED",
			x"0000" when x"72EE",
			x"0000" when x"72EF",
			x"0000" when x"72F0",
			x"0000" when x"72F1",
			x"0000" when x"72F2",
			x"0000" when x"72F3",
			x"0000" when x"72F4",
			x"0000" when x"72F5",
			x"0000" when x"72F6",
			x"0000" when x"72F7",
			x"0000" when x"72F8",
			x"0000" when x"72F9",
			x"0000" when x"72FA",
			x"0000" when x"72FB",
			x"0000" when x"72FC",
			x"0000" when x"72FD",
			x"0000" when x"72FE",
			x"0000" when x"72FF",
			x"0000" when x"7300",
			x"0000" when x"7301",
			x"0000" when x"7302",
			x"0000" when x"7303",
			x"0000" when x"7304",
			x"0000" when x"7305",
			x"0000" when x"7306",
			x"0000" when x"7307",
			x"0000" when x"7308",
			x"0000" when x"7309",
			x"0000" when x"730A",
			x"0000" when x"730B",
			x"0000" when x"730C",
			x"0000" when x"730D",
			x"0000" when x"730E",
			x"0000" when x"730F",
			x"0000" when x"7310",
			x"0000" when x"7311",
			x"0000" when x"7312",
			x"0000" when x"7313",
			x"0000" when x"7314",
			x"0000" when x"7315",
			x"0000" when x"7316",
			x"0000" when x"7317",
			x"0000" when x"7318",
			x"0000" when x"7319",
			x"0000" when x"731A",
			x"0000" when x"731B",
			x"0000" when x"731C",
			x"0000" when x"731D",
			x"0000" when x"731E",
			x"0000" when x"731F",
			x"0000" when x"7320",
			x"0000" when x"7321",
			x"0000" when x"7322",
			x"0000" when x"7323",
			x"0000" when x"7324",
			x"0000" when x"7325",
			x"0000" when x"7326",
			x"0000" when x"7327",
			x"0000" when x"7328",
			x"0000" when x"7329",
			x"0000" when x"732A",
			x"0000" when x"732B",
			x"0000" when x"732C",
			x"0000" when x"732D",
			x"0000" when x"732E",
			x"0000" when x"732F",
			x"0000" when x"7330",
			x"0000" when x"7331",
			x"0000" when x"7332",
			x"0000" when x"7333",
			x"0000" when x"7334",
			x"0000" when x"7335",
			x"0000" when x"7336",
			x"0000" when x"7337",
			x"0000" when x"7338",
			x"0000" when x"7339",
			x"0000" when x"733A",
			x"0000" when x"733B",
			x"0000" when x"733C",
			x"0000" when x"733D",
			x"0000" when x"733E",
			x"0000" when x"733F",
			x"0000" when x"7340",
			x"0000" when x"7341",
			x"0000" when x"7342",
			x"0000" when x"7343",
			x"0000" when x"7344",
			x"0000" when x"7345",
			x"0000" when x"7346",
			x"0000" when x"7347",
			x"0000" when x"7348",
			x"0000" when x"7349",
			x"0000" when x"734A",
			x"0000" when x"734B",
			x"0000" when x"734C",
			x"0000" when x"734D",
			x"0000" when x"734E",
			x"0000" when x"734F",
			x"0000" when x"7350",
			x"0000" when x"7351",
			x"0000" when x"7352",
			x"0000" when x"7353",
			x"0000" when x"7354",
			x"0000" when x"7355",
			x"0000" when x"7356",
			x"0000" when x"7357",
			x"0000" when x"7358",
			x"0000" when x"7359",
			x"0000" when x"735A",
			x"0000" when x"735B",
			x"0000" when x"735C",
			x"0000" when x"735D",
			x"0000" when x"735E",
			x"0000" when x"735F",
			x"0000" when x"7360",
			x"0000" when x"7361",
			x"0000" when x"7362",
			x"0000" when x"7363",
			x"0000" when x"7364",
			x"0000" when x"7365",
			x"0000" when x"7366",
			x"0000" when x"7367",
			x"0000" when x"7368",
			x"0000" when x"7369",
			x"0000" when x"736A",
			x"0000" when x"736B",
			x"0000" when x"736C",
			x"0000" when x"736D",
			x"0000" when x"736E",
			x"0000" when x"736F",
			x"0000" when x"7370",
			x"0000" when x"7371",
			x"0000" when x"7372",
			x"0000" when x"7373",
			x"0000" when x"7374",
			x"0000" when x"7375",
			x"0000" when x"7376",
			x"0000" when x"7377",
			x"0000" when x"7378",
			x"0000" when x"7379",
			x"0000" when x"737A",
			x"0000" when x"737B",
			x"0000" when x"737C",
			x"0000" when x"737D",
			x"0000" when x"737E",
			x"0000" when x"737F",
			x"0000" when x"7380",
			x"0000" when x"7381",
			x"0000" when x"7382",
			x"0000" when x"7383",
			x"0000" when x"7384",
			x"0000" when x"7385",
			x"0000" when x"7386",
			x"0000" when x"7387",
			x"0000" when x"7388",
			x"0000" when x"7389",
			x"0000" when x"738A",
			x"0000" when x"738B",
			x"0000" when x"738C",
			x"0000" when x"738D",
			x"0000" when x"738E",
			x"0000" when x"738F",
			x"0000" when x"7390",
			x"0000" when x"7391",
			x"0000" when x"7392",
			x"0000" when x"7393",
			x"0000" when x"7394",
			x"0000" when x"7395",
			x"0000" when x"7396",
			x"0000" when x"7397",
			x"0000" when x"7398",
			x"0000" when x"7399",
			x"0000" when x"739A",
			x"0000" when x"739B",
			x"0000" when x"739C",
			x"0000" when x"739D",
			x"0000" when x"739E",
			x"0000" when x"739F",
			x"0000" when x"73A0",
			x"0000" when x"73A1",
			x"0000" when x"73A2",
			x"0000" when x"73A3",
			x"0000" when x"73A4",
			x"0000" when x"73A5",
			x"0000" when x"73A6",
			x"0000" when x"73A7",
			x"0000" when x"73A8",
			x"0000" when x"73A9",
			x"0000" when x"73AA",
			x"0000" when x"73AB",
			x"0000" when x"73AC",
			x"0000" when x"73AD",
			x"0000" when x"73AE",
			x"0000" when x"73AF",
			x"0000" when x"73B0",
			x"0000" when x"73B1",
			x"0000" when x"73B2",
			x"0000" when x"73B3",
			x"0000" when x"73B4",
			x"0000" when x"73B5",
			x"0000" when x"73B6",
			x"0000" when x"73B7",
			x"0000" when x"73B8",
			x"0000" when x"73B9",
			x"0000" when x"73BA",
			x"0000" when x"73BB",
			x"0000" when x"73BC",
			x"0000" when x"73BD",
			x"0000" when x"73BE",
			x"0000" when x"73BF",
			x"0000" when x"73C0",
			x"0000" when x"73C1",
			x"0000" when x"73C2",
			x"0000" when x"73C3",
			x"0000" when x"73C4",
			x"0000" when x"73C5",
			x"0000" when x"73C6",
			x"0000" when x"73C7",
			x"0000" when x"73C8",
			x"0000" when x"73C9",
			x"0000" when x"73CA",
			x"0000" when x"73CB",
			x"0000" when x"73CC",
			x"0000" when x"73CD",
			x"0000" when x"73CE",
			x"0000" when x"73CF",
			x"0000" when x"73D0",
			x"0000" when x"73D1",
			x"0000" when x"73D2",
			x"0000" when x"73D3",
			x"0000" when x"73D4",
			x"0000" when x"73D5",
			x"0000" when x"73D6",
			x"0000" when x"73D7",
			x"0000" when x"73D8",
			x"0000" when x"73D9",
			x"0000" when x"73DA",
			x"0000" when x"73DB",
			x"0000" when x"73DC",
			x"0000" when x"73DD",
			x"0000" when x"73DE",
			x"0000" when x"73DF",
			x"0000" when x"73E0",
			x"0000" when x"73E1",
			x"0000" when x"73E2",
			x"0000" when x"73E3",
			x"0000" when x"73E4",
			x"0000" when x"73E5",
			x"0000" when x"73E6",
			x"0000" when x"73E7",
			x"0000" when x"73E8",
			x"0000" when x"73E9",
			x"0000" when x"73EA",
			x"0000" when x"73EB",
			x"0000" when x"73EC",
			x"0000" when x"73ED",
			x"0000" when x"73EE",
			x"0000" when x"73EF",
			x"0000" when x"73F0",
			x"0000" when x"73F1",
			x"0000" when x"73F2",
			x"0000" when x"73F3",
			x"0000" when x"73F4",
			x"0000" when x"73F5",
			x"0000" when x"73F6",
			x"0000" when x"73F7",
			x"0000" when x"73F8",
			x"0000" when x"73F9",
			x"0000" when x"73FA",
			x"0000" when x"73FB",
			x"0000" when x"73FC",
			x"0000" when x"73FD",
			x"0000" when x"73FE",
			x"0000" when x"73FF",
			x"0000" when x"7400",
			x"0000" when x"7401",
			x"0000" when x"7402",
			x"0000" when x"7403",
			x"0000" when x"7404",
			x"0000" when x"7405",
			x"0000" when x"7406",
			x"0000" when x"7407",
			x"0000" when x"7408",
			x"0000" when x"7409",
			x"0000" when x"740A",
			x"0000" when x"740B",
			x"0000" when x"740C",
			x"0000" when x"740D",
			x"0000" when x"740E",
			x"0000" when x"740F",
			x"0000" when x"7410",
			x"0000" when x"7411",
			x"0000" when x"7412",
			x"0000" when x"7413",
			x"0000" when x"7414",
			x"0000" when x"7415",
			x"0000" when x"7416",
			x"0000" when x"7417",
			x"0000" when x"7418",
			x"0000" when x"7419",
			x"0000" when x"741A",
			x"0000" when x"741B",
			x"0000" when x"741C",
			x"0000" when x"741D",
			x"0000" when x"741E",
			x"0000" when x"741F",
			x"0000" when x"7420",
			x"0000" when x"7421",
			x"0000" when x"7422",
			x"0000" when x"7423",
			x"0000" when x"7424",
			x"0000" when x"7425",
			x"0000" when x"7426",
			x"0000" when x"7427",
			x"0000" when x"7428",
			x"0000" when x"7429",
			x"0000" when x"742A",
			x"0000" when x"742B",
			x"0000" when x"742C",
			x"0000" when x"742D",
			x"0000" when x"742E",
			x"0000" when x"742F",
			x"0000" when x"7430",
			x"0000" when x"7431",
			x"0000" when x"7432",
			x"0000" when x"7433",
			x"0000" when x"7434",
			x"0000" when x"7435",
			x"0000" when x"7436",
			x"0000" when x"7437",
			x"0000" when x"7438",
			x"0000" when x"7439",
			x"0000" when x"743A",
			x"0000" when x"743B",
			x"0000" when x"743C",
			x"0000" when x"743D",
			x"0000" when x"743E",
			x"0000" when x"743F",
			x"0000" when x"7440",
			x"0000" when x"7441",
			x"0000" when x"7442",
			x"0000" when x"7443",
			x"0000" when x"7444",
			x"0000" when x"7445",
			x"0000" when x"7446",
			x"0000" when x"7447",
			x"0000" when x"7448",
			x"0000" when x"7449",
			x"0000" when x"744A",
			x"0000" when x"744B",
			x"0000" when x"744C",
			x"0000" when x"744D",
			x"0000" when x"744E",
			x"0000" when x"744F",
			x"0000" when x"7450",
			x"0000" when x"7451",
			x"0000" when x"7452",
			x"0000" when x"7453",
			x"0000" when x"7454",
			x"0000" when x"7455",
			x"0000" when x"7456",
			x"0000" when x"7457",
			x"0000" when x"7458",
			x"0000" when x"7459",
			x"0000" when x"745A",
			x"0000" when x"745B",
			x"0000" when x"745C",
			x"0000" when x"745D",
			x"0000" when x"745E",
			x"0000" when x"745F",
			x"0000" when x"7460",
			x"0000" when x"7461",
			x"0000" when x"7462",
			x"0000" when x"7463",
			x"0000" when x"7464",
			x"0000" when x"7465",
			x"0000" when x"7466",
			x"0000" when x"7467",
			x"0000" when x"7468",
			x"0000" when x"7469",
			x"0000" when x"746A",
			x"0000" when x"746B",
			x"0000" when x"746C",
			x"0000" when x"746D",
			x"0000" when x"746E",
			x"0000" when x"746F",
			x"0000" when x"7470",
			x"0000" when x"7471",
			x"0000" when x"7472",
			x"0000" when x"7473",
			x"0000" when x"7474",
			x"0000" when x"7475",
			x"0000" when x"7476",
			x"0000" when x"7477",
			x"0000" when x"7478",
			x"0000" when x"7479",
			x"0000" when x"747A",
			x"0000" when x"747B",
			x"0000" when x"747C",
			x"0000" when x"747D",
			x"0000" when x"747E",
			x"0000" when x"747F",
			x"0000" when x"7480",
			x"0000" when x"7481",
			x"0000" when x"7482",
			x"0000" when x"7483",
			x"0000" when x"7484",
			x"0000" when x"7485",
			x"0000" when x"7486",
			x"0000" when x"7487",
			x"0000" when x"7488",
			x"0000" when x"7489",
			x"0000" when x"748A",
			x"0000" when x"748B",
			x"0000" when x"748C",
			x"0000" when x"748D",
			x"0000" when x"748E",
			x"0000" when x"748F",
			x"0000" when x"7490",
			x"0000" when x"7491",
			x"0000" when x"7492",
			x"0000" when x"7493",
			x"0000" when x"7494",
			x"0000" when x"7495",
			x"0000" when x"7496",
			x"0000" when x"7497",
			x"0000" when x"7498",
			x"0000" when x"7499",
			x"0000" when x"749A",
			x"0000" when x"749B",
			x"0000" when x"749C",
			x"0000" when x"749D",
			x"0000" when x"749E",
			x"0000" when x"749F",
			x"0000" when x"74A0",
			x"0000" when x"74A1",
			x"0000" when x"74A2",
			x"0000" when x"74A3",
			x"0000" when x"74A4",
			x"0000" when x"74A5",
			x"0000" when x"74A6",
			x"0000" when x"74A7",
			x"0000" when x"74A8",
			x"0000" when x"74A9",
			x"0000" when x"74AA",
			x"0000" when x"74AB",
			x"0000" when x"74AC",
			x"0000" when x"74AD",
			x"0000" when x"74AE",
			x"0000" when x"74AF",
			x"0000" when x"74B0",
			x"0000" when x"74B1",
			x"0000" when x"74B2",
			x"0000" when x"74B3",
			x"0000" when x"74B4",
			x"0000" when x"74B5",
			x"0000" when x"74B6",
			x"0000" when x"74B7",
			x"0000" when x"74B8",
			x"0000" when x"74B9",
			x"0000" when x"74BA",
			x"0000" when x"74BB",
			x"0000" when x"74BC",
			x"0000" when x"74BD",
			x"0000" when x"74BE",
			x"0000" when x"74BF",
			x"0000" when x"74C0",
			x"0000" when x"74C1",
			x"0000" when x"74C2",
			x"0000" when x"74C3",
			x"0000" when x"74C4",
			x"0000" when x"74C5",
			x"0000" when x"74C6",
			x"0000" when x"74C7",
			x"0000" when x"74C8",
			x"0000" when x"74C9",
			x"0000" when x"74CA",
			x"0000" when x"74CB",
			x"0000" when x"74CC",
			x"0000" when x"74CD",
			x"0000" when x"74CE",
			x"0000" when x"74CF",
			x"0000" when x"74D0",
			x"0000" when x"74D1",
			x"0000" when x"74D2",
			x"0000" when x"74D3",
			x"0000" when x"74D4",
			x"0000" when x"74D5",
			x"0000" when x"74D6",
			x"0000" when x"74D7",
			x"0000" when x"74D8",
			x"0000" when x"74D9",
			x"0000" when x"74DA",
			x"0000" when x"74DB",
			x"0000" when x"74DC",
			x"0000" when x"74DD",
			x"0000" when x"74DE",
			x"0000" when x"74DF",
			x"0000" when x"74E0",
			x"0000" when x"74E1",
			x"0000" when x"74E2",
			x"0000" when x"74E3",
			x"0000" when x"74E4",
			x"0000" when x"74E5",
			x"0000" when x"74E6",
			x"0000" when x"74E7",
			x"0000" when x"74E8",
			x"0000" when x"74E9",
			x"0000" when x"74EA",
			x"0000" when x"74EB",
			x"0000" when x"74EC",
			x"0000" when x"74ED",
			x"0000" when x"74EE",
			x"0000" when x"74EF",
			x"0000" when x"74F0",
			x"0000" when x"74F1",
			x"0000" when x"74F2",
			x"0000" when x"74F3",
			x"0000" when x"74F4",
			x"0000" when x"74F5",
			x"0000" when x"74F6",
			x"0000" when x"74F7",
			x"0000" when x"74F8",
			x"0000" when x"74F9",
			x"0000" when x"74FA",
			x"0000" when x"74FB",
			x"0000" when x"74FC",
			x"0000" when x"74FD",
			x"0000" when x"74FE",
			x"0000" when x"74FF",
			x"0000" when x"7500",
			x"0000" when x"7501",
			x"0000" when x"7502",
			x"0000" when x"7503",
			x"0000" when x"7504",
			x"0000" when x"7505",
			x"0000" when x"7506",
			x"0000" when x"7507",
			x"0000" when x"7508",
			x"0000" when x"7509",
			x"0000" when x"750A",
			x"0000" when x"750B",
			x"0000" when x"750C",
			x"0000" when x"750D",
			x"0000" when x"750E",
			x"0000" when x"750F",
			x"0000" when x"7510",
			x"0000" when x"7511",
			x"0000" when x"7512",
			x"0000" when x"7513",
			x"0000" when x"7514",
			x"0000" when x"7515",
			x"0000" when x"7516",
			x"0000" when x"7517",
			x"0000" when x"7518",
			x"0000" when x"7519",
			x"0000" when x"751A",
			x"0000" when x"751B",
			x"0000" when x"751C",
			x"0000" when x"751D",
			x"0000" when x"751E",
			x"0000" when x"751F",
			x"0000" when x"7520",
			x"0000" when x"7521",
			x"0000" when x"7522",
			x"0000" when x"7523",
			x"0000" when x"7524",
			x"0000" when x"7525",
			x"0000" when x"7526",
			x"0000" when x"7527",
			x"0000" when x"7528",
			x"0000" when x"7529",
			x"0000" when x"752A",
			x"0000" when x"752B",
			x"0000" when x"752C",
			x"0000" when x"752D",
			x"0000" when x"752E",
			x"0000" when x"752F",
			x"0000" when x"7530",
			x"0000" when x"7531",
			x"0000" when x"7532",
			x"0000" when x"7533",
			x"0000" when x"7534",
			x"0000" when x"7535",
			x"0000" when x"7536",
			x"0000" when x"7537",
			x"0000" when x"7538",
			x"0000" when x"7539",
			x"0000" when x"753A",
			x"0000" when x"753B",
			x"0000" when x"753C",
			x"0000" when x"753D",
			x"0000" when x"753E",
			x"0000" when x"753F",
			x"0000" when x"7540",
			x"0000" when x"7541",
			x"0000" when x"7542",
			x"0000" when x"7543",
			x"0000" when x"7544",
			x"0000" when x"7545",
			x"0000" when x"7546",
			x"0000" when x"7547",
			x"0000" when x"7548",
			x"0000" when x"7549",
			x"0000" when x"754A",
			x"0000" when x"754B",
			x"0000" when x"754C",
			x"0000" when x"754D",
			x"0000" when x"754E",
			x"0000" when x"754F",
			x"0000" when x"7550",
			x"0000" when x"7551",
			x"0000" when x"7552",
			x"0000" when x"7553",
			x"0000" when x"7554",
			x"0000" when x"7555",
			x"0000" when x"7556",
			x"0000" when x"7557",
			x"0000" when x"7558",
			x"0000" when x"7559",
			x"0000" when x"755A",
			x"0000" when x"755B",
			x"0000" when x"755C",
			x"0000" when x"755D",
			x"0000" when x"755E",
			x"0000" when x"755F",
			x"0000" when x"7560",
			x"0000" when x"7561",
			x"0000" when x"7562",
			x"0000" when x"7563",
			x"0000" when x"7564",
			x"0000" when x"7565",
			x"0000" when x"7566",
			x"0000" when x"7567",
			x"0000" when x"7568",
			x"0000" when x"7569",
			x"0000" when x"756A",
			x"0000" when x"756B",
			x"0000" when x"756C",
			x"0000" when x"756D",
			x"0000" when x"756E",
			x"0000" when x"756F",
			x"0000" when x"7570",
			x"0000" when x"7571",
			x"0000" when x"7572",
			x"0000" when x"7573",
			x"0000" when x"7574",
			x"0000" when x"7575",
			x"0000" when x"7576",
			x"0000" when x"7577",
			x"0000" when x"7578",
			x"0000" when x"7579",
			x"0000" when x"757A",
			x"0000" when x"757B",
			x"0000" when x"757C",
			x"0000" when x"757D",
			x"0000" when x"757E",
			x"0000" when x"757F",
			x"0000" when x"7580",
			x"0000" when x"7581",
			x"0000" when x"7582",
			x"0000" when x"7583",
			x"0000" when x"7584",
			x"0000" when x"7585",
			x"0000" when x"7586",
			x"0000" when x"7587",
			x"0000" when x"7588",
			x"0000" when x"7589",
			x"0000" when x"758A",
			x"0000" when x"758B",
			x"0000" when x"758C",
			x"0000" when x"758D",
			x"0000" when x"758E",
			x"0000" when x"758F",
			x"0000" when x"7590",
			x"0000" when x"7591",
			x"0000" when x"7592",
			x"0000" when x"7593",
			x"0000" when x"7594",
			x"0000" when x"7595",
			x"0000" when x"7596",
			x"0000" when x"7597",
			x"0000" when x"7598",
			x"0000" when x"7599",
			x"0000" when x"759A",
			x"0000" when x"759B",
			x"0000" when x"759C",
			x"0000" when x"759D",
			x"0000" when x"759E",
			x"0000" when x"759F",
			x"0000" when x"75A0",
			x"0000" when x"75A1",
			x"0000" when x"75A2",
			x"0000" when x"75A3",
			x"0000" when x"75A4",
			x"0000" when x"75A5",
			x"0000" when x"75A6",
			x"0000" when x"75A7",
			x"0000" when x"75A8",
			x"0000" when x"75A9",
			x"0000" when x"75AA",
			x"0000" when x"75AB",
			x"0000" when x"75AC",
			x"0000" when x"75AD",
			x"0000" when x"75AE",
			x"0000" when x"75AF",
			x"0000" when x"75B0",
			x"0000" when x"75B1",
			x"0000" when x"75B2",
			x"0000" when x"75B3",
			x"0000" when x"75B4",
			x"0000" when x"75B5",
			x"0000" when x"75B6",
			x"0000" when x"75B7",
			x"0000" when x"75B8",
			x"0000" when x"75B9",
			x"0000" when x"75BA",
			x"0000" when x"75BB",
			x"0000" when x"75BC",
			x"0000" when x"75BD",
			x"0000" when x"75BE",
			x"0000" when x"75BF",
			x"0000" when x"75C0",
			x"0000" when x"75C1",
			x"0000" when x"75C2",
			x"0000" when x"75C3",
			x"0000" when x"75C4",
			x"0000" when x"75C5",
			x"0000" when x"75C6",
			x"0000" when x"75C7",
			x"0000" when x"75C8",
			x"0000" when x"75C9",
			x"0000" when x"75CA",
			x"0000" when x"75CB",
			x"0000" when x"75CC",
			x"0000" when x"75CD",
			x"0000" when x"75CE",
			x"0000" when x"75CF",
			x"0000" when x"75D0",
			x"0000" when x"75D1",
			x"0000" when x"75D2",
			x"0000" when x"75D3",
			x"0000" when x"75D4",
			x"0000" when x"75D5",
			x"0000" when x"75D6",
			x"0000" when x"75D7",
			x"0000" when x"75D8",
			x"0000" when x"75D9",
			x"0000" when x"75DA",
			x"0000" when x"75DB",
			x"0000" when x"75DC",
			x"0000" when x"75DD",
			x"0000" when x"75DE",
			x"0000" when x"75DF",
			x"0000" when x"75E0",
			x"0000" when x"75E1",
			x"0000" when x"75E2",
			x"0000" when x"75E3",
			x"0000" when x"75E4",
			x"0000" when x"75E5",
			x"0000" when x"75E6",
			x"0000" when x"75E7",
			x"0000" when x"75E8",
			x"0000" when x"75E9",
			x"0000" when x"75EA",
			x"0000" when x"75EB",
			x"0000" when x"75EC",
			x"0000" when x"75ED",
			x"0000" when x"75EE",
			x"0000" when x"75EF",
			x"0000" when x"75F0",
			x"0000" when x"75F1",
			x"0000" when x"75F2",
			x"0000" when x"75F3",
			x"0000" when x"75F4",
			x"0000" when x"75F5",
			x"0000" when x"75F6",
			x"0000" when x"75F7",
			x"0000" when x"75F8",
			x"0000" when x"75F9",
			x"0000" when x"75FA",
			x"0000" when x"75FB",
			x"0000" when x"75FC",
			x"0000" when x"75FD",
			x"0000" when x"75FE",
			x"0000" when x"75FF",
			x"0000" when x"7600",
			x"0000" when x"7601",
			x"0000" when x"7602",
			x"0000" when x"7603",
			x"0000" when x"7604",
			x"0000" when x"7605",
			x"0000" when x"7606",
			x"0000" when x"7607",
			x"0000" when x"7608",
			x"0000" when x"7609",
			x"0000" when x"760A",
			x"0000" when x"760B",
			x"0000" when x"760C",
			x"0000" when x"760D",
			x"0000" when x"760E",
			x"0000" when x"760F",
			x"0000" when x"7610",
			x"0000" when x"7611",
			x"0000" when x"7612",
			x"0000" when x"7613",
			x"0000" when x"7614",
			x"0000" when x"7615",
			x"0000" when x"7616",
			x"0000" when x"7617",
			x"0000" when x"7618",
			x"0000" when x"7619",
			x"0000" when x"761A",
			x"0000" when x"761B",
			x"0000" when x"761C",
			x"0000" when x"761D",
			x"0000" when x"761E",
			x"0000" when x"761F",
			x"0000" when x"7620",
			x"0000" when x"7621",
			x"0000" when x"7622",
			x"0000" when x"7623",
			x"0000" when x"7624",
			x"0000" when x"7625",
			x"0000" when x"7626",
			x"0000" when x"7627",
			x"0000" when x"7628",
			x"0000" when x"7629",
			x"0000" when x"762A",
			x"0000" when x"762B",
			x"0000" when x"762C",
			x"0000" when x"762D",
			x"0000" when x"762E",
			x"0000" when x"762F",
			x"0000" when x"7630",
			x"0000" when x"7631",
			x"0000" when x"7632",
			x"0000" when x"7633",
			x"0000" when x"7634",
			x"0000" when x"7635",
			x"0000" when x"7636",
			x"0000" when x"7637",
			x"0000" when x"7638",
			x"0000" when x"7639",
			x"0000" when x"763A",
			x"0000" when x"763B",
			x"0000" when x"763C",
			x"0000" when x"763D",
			x"0000" when x"763E",
			x"0000" when x"763F",
			x"0000" when x"7640",
			x"0000" when x"7641",
			x"0000" when x"7642",
			x"0000" when x"7643",
			x"0000" when x"7644",
			x"0000" when x"7645",
			x"0000" when x"7646",
			x"0000" when x"7647",
			x"0000" when x"7648",
			x"0000" when x"7649",
			x"0000" when x"764A",
			x"0000" when x"764B",
			x"0000" when x"764C",
			x"0000" when x"764D",
			x"0000" when x"764E",
			x"0000" when x"764F",
			x"0000" when x"7650",
			x"0000" when x"7651",
			x"0000" when x"7652",
			x"0000" when x"7653",
			x"0000" when x"7654",
			x"0000" when x"7655",
			x"0000" when x"7656",
			x"0000" when x"7657",
			x"0000" when x"7658",
			x"0000" when x"7659",
			x"0000" when x"765A",
			x"0000" when x"765B",
			x"0000" when x"765C",
			x"0000" when x"765D",
			x"0000" when x"765E",
			x"0000" when x"765F",
			x"0000" when x"7660",
			x"0000" when x"7661",
			x"0000" when x"7662",
			x"0000" when x"7663",
			x"0000" when x"7664",
			x"0000" when x"7665",
			x"0000" when x"7666",
			x"0000" when x"7667",
			x"0000" when x"7668",
			x"0000" when x"7669",
			x"0000" when x"766A",
			x"0000" when x"766B",
			x"0000" when x"766C",
			x"0000" when x"766D",
			x"0000" when x"766E",
			x"0000" when x"766F",
			x"0000" when x"7670",
			x"0000" when x"7671",
			x"0000" when x"7672",
			x"0000" when x"7673",
			x"0000" when x"7674",
			x"0000" when x"7675",
			x"0000" when x"7676",
			x"0000" when x"7677",
			x"0000" when x"7678",
			x"0000" when x"7679",
			x"0000" when x"767A",
			x"0000" when x"767B",
			x"0000" when x"767C",
			x"0000" when x"767D",
			x"0000" when x"767E",
			x"0000" when x"767F",
			x"0000" when x"7680",
			x"0000" when x"7681",
			x"0000" when x"7682",
			x"0000" when x"7683",
			x"0000" when x"7684",
			x"0000" when x"7685",
			x"0000" when x"7686",
			x"0000" when x"7687",
			x"0000" when x"7688",
			x"0000" when x"7689",
			x"0000" when x"768A",
			x"0000" when x"768B",
			x"0000" when x"768C",
			x"0000" when x"768D",
			x"0000" when x"768E",
			x"0000" when x"768F",
			x"0000" when x"7690",
			x"0000" when x"7691",
			x"0000" when x"7692",
			x"0000" when x"7693",
			x"0000" when x"7694",
			x"0000" when x"7695",
			x"0000" when x"7696",
			x"0000" when x"7697",
			x"0000" when x"7698",
			x"0000" when x"7699",
			x"0000" when x"769A",
			x"0000" when x"769B",
			x"0000" when x"769C",
			x"0000" when x"769D",
			x"0000" when x"769E",
			x"0000" when x"769F",
			x"0000" when x"76A0",
			x"0000" when x"76A1",
			x"0000" when x"76A2",
			x"0000" when x"76A3",
			x"0000" when x"76A4",
			x"0000" when x"76A5",
			x"0000" when x"76A6",
			x"0000" when x"76A7",
			x"0000" when x"76A8",
			x"0000" when x"76A9",
			x"0000" when x"76AA",
			x"0000" when x"76AB",
			x"0000" when x"76AC",
			x"0000" when x"76AD",
			x"0000" when x"76AE",
			x"0000" when x"76AF",
			x"0000" when x"76B0",
			x"0000" when x"76B1",
			x"0000" when x"76B2",
			x"0000" when x"76B3",
			x"0000" when x"76B4",
			x"0000" when x"76B5",
			x"0000" when x"76B6",
			x"0000" when x"76B7",
			x"0000" when x"76B8",
			x"0000" when x"76B9",
			x"0000" when x"76BA",
			x"0000" when x"76BB",
			x"0000" when x"76BC",
			x"0000" when x"76BD",
			x"0000" when x"76BE",
			x"0000" when x"76BF",
			x"0000" when x"76C0",
			x"0000" when x"76C1",
			x"0000" when x"76C2",
			x"0000" when x"76C3",
			x"0000" when x"76C4",
			x"0000" when x"76C5",
			x"0000" when x"76C6",
			x"0000" when x"76C7",
			x"0000" when x"76C8",
			x"0000" when x"76C9",
			x"0000" when x"76CA",
			x"0000" when x"76CB",
			x"0000" when x"76CC",
			x"0000" when x"76CD",
			x"0000" when x"76CE",
			x"0000" when x"76CF",
			x"0000" when x"76D0",
			x"0000" when x"76D1",
			x"0000" when x"76D2",
			x"0000" when x"76D3",
			x"0000" when x"76D4",
			x"0000" when x"76D5",
			x"0000" when x"76D6",
			x"0000" when x"76D7",
			x"0000" when x"76D8",
			x"0000" when x"76D9",
			x"0000" when x"76DA",
			x"0000" when x"76DB",
			x"0000" when x"76DC",
			x"0000" when x"76DD",
			x"0000" when x"76DE",
			x"0000" when x"76DF",
			x"0000" when x"76E0",
			x"0000" when x"76E1",
			x"0000" when x"76E2",
			x"0000" when x"76E3",
			x"0000" when x"76E4",
			x"0000" when x"76E5",
			x"0000" when x"76E6",
			x"0000" when x"76E7",
			x"0000" when x"76E8",
			x"0000" when x"76E9",
			x"0000" when x"76EA",
			x"0000" when x"76EB",
			x"0000" when x"76EC",
			x"0000" when x"76ED",
			x"0000" when x"76EE",
			x"0000" when x"76EF",
			x"0000" when x"76F0",
			x"0000" when x"76F1",
			x"0000" when x"76F2",
			x"0000" when x"76F3",
			x"0000" when x"76F4",
			x"0000" when x"76F5",
			x"0000" when x"76F6",
			x"0000" when x"76F7",
			x"0000" when x"76F8",
			x"0000" when x"76F9",
			x"0000" when x"76FA",
			x"0000" when x"76FB",
			x"0000" when x"76FC",
			x"0000" when x"76FD",
			x"0000" when x"76FE",
			x"0000" when x"76FF",
			x"0000" when x"7700",
			x"0000" when x"7701",
			x"0000" when x"7702",
			x"0000" when x"7703",
			x"0000" when x"7704",
			x"0000" when x"7705",
			x"0000" when x"7706",
			x"0000" when x"7707",
			x"0000" when x"7708",
			x"0000" when x"7709",
			x"0000" when x"770A",
			x"0000" when x"770B",
			x"0000" when x"770C",
			x"0000" when x"770D",
			x"0000" when x"770E",
			x"0000" when x"770F",
			x"0000" when x"7710",
			x"0000" when x"7711",
			x"0000" when x"7712",
			x"0000" when x"7713",
			x"0000" when x"7714",
			x"0000" when x"7715",
			x"0000" when x"7716",
			x"0000" when x"7717",
			x"0000" when x"7718",
			x"0000" when x"7719",
			x"0000" when x"771A",
			x"0000" when x"771B",
			x"0000" when x"771C",
			x"0000" when x"771D",
			x"0000" when x"771E",
			x"0000" when x"771F",
			x"0000" when x"7720",
			x"0000" when x"7721",
			x"0000" when x"7722",
			x"0000" when x"7723",
			x"0000" when x"7724",
			x"0000" when x"7725",
			x"0000" when x"7726",
			x"0000" when x"7727",
			x"0000" when x"7728",
			x"0000" when x"7729",
			x"0000" when x"772A",
			x"0000" when x"772B",
			x"0000" when x"772C",
			x"0000" when x"772D",
			x"0000" when x"772E",
			x"0000" when x"772F",
			x"0000" when x"7730",
			x"0000" when x"7731",
			x"0000" when x"7732",
			x"0000" when x"7733",
			x"0000" when x"7734",
			x"0000" when x"7735",
			x"0000" when x"7736",
			x"0000" when x"7737",
			x"0000" when x"7738",
			x"0000" when x"7739",
			x"0000" when x"773A",
			x"0000" when x"773B",
			x"0000" when x"773C",
			x"0000" when x"773D",
			x"0000" when x"773E",
			x"0000" when x"773F",
			x"0000" when x"7740",
			x"0000" when x"7741",
			x"0000" when x"7742",
			x"0000" when x"7743",
			x"0000" when x"7744",
			x"0000" when x"7745",
			x"0000" when x"7746",
			x"0000" when x"7747",
			x"0000" when x"7748",
			x"0000" when x"7749",
			x"0000" when x"774A",
			x"0000" when x"774B",
			x"0000" when x"774C",
			x"0000" when x"774D",
			x"0000" when x"774E",
			x"0000" when x"774F",
			x"0000" when x"7750",
			x"0000" when x"7751",
			x"0000" when x"7752",
			x"0000" when x"7753",
			x"0000" when x"7754",
			x"0000" when x"7755",
			x"0000" when x"7756",
			x"0000" when x"7757",
			x"0000" when x"7758",
			x"0000" when x"7759",
			x"0000" when x"775A",
			x"0000" when x"775B",
			x"0000" when x"775C",
			x"0000" when x"775D",
			x"0000" when x"775E",
			x"0000" when x"775F",
			x"0000" when x"7760",
			x"0000" when x"7761",
			x"0000" when x"7762",
			x"0000" when x"7763",
			x"0000" when x"7764",
			x"0000" when x"7765",
			x"0000" when x"7766",
			x"0000" when x"7767",
			x"0000" when x"7768",
			x"0000" when x"7769",
			x"0000" when x"776A",
			x"0000" when x"776B",
			x"0000" when x"776C",
			x"0000" when x"776D",
			x"0000" when x"776E",
			x"0000" when x"776F",
			x"0000" when x"7770",
			x"0000" when x"7771",
			x"0000" when x"7772",
			x"0000" when x"7773",
			x"0000" when x"7774",
			x"0000" when x"7775",
			x"0000" when x"7776",
			x"0000" when x"7777",
			x"0000" when x"7778",
			x"0000" when x"7779",
			x"0000" when x"777A",
			x"0000" when x"777B",
			x"0000" when x"777C",
			x"0000" when x"777D",
			x"0000" when x"777E",
			x"0000" when x"777F",
			x"0000" when x"7780",
			x"0000" when x"7781",
			x"0000" when x"7782",
			x"0000" when x"7783",
			x"0000" when x"7784",
			x"0000" when x"7785",
			x"0000" when x"7786",
			x"0000" when x"7787",
			x"0000" when x"7788",
			x"0000" when x"7789",
			x"0000" when x"778A",
			x"0000" when x"778B",
			x"0000" when x"778C",
			x"0000" when x"778D",
			x"0000" when x"778E",
			x"0000" when x"778F",
			x"0000" when x"7790",
			x"0000" when x"7791",
			x"0000" when x"7792",
			x"0000" when x"7793",
			x"0000" when x"7794",
			x"0000" when x"7795",
			x"0000" when x"7796",
			x"0000" when x"7797",
			x"0000" when x"7798",
			x"0000" when x"7799",
			x"0000" when x"779A",
			x"0000" when x"779B",
			x"0000" when x"779C",
			x"0000" when x"779D",
			x"0000" when x"779E",
			x"0000" when x"779F",
			x"0000" when x"77A0",
			x"0000" when x"77A1",
			x"0000" when x"77A2",
			x"0000" when x"77A3",
			x"0000" when x"77A4",
			x"0000" when x"77A5",
			x"0000" when x"77A6",
			x"0000" when x"77A7",
			x"0000" when x"77A8",
			x"0000" when x"77A9",
			x"0000" when x"77AA",
			x"0000" when x"77AB",
			x"0000" when x"77AC",
			x"0000" when x"77AD",
			x"0000" when x"77AE",
			x"0000" when x"77AF",
			x"0000" when x"77B0",
			x"0000" when x"77B1",
			x"0000" when x"77B2",
			x"0000" when x"77B3",
			x"0000" when x"77B4",
			x"0000" when x"77B5",
			x"0000" when x"77B6",
			x"0000" when x"77B7",
			x"0000" when x"77B8",
			x"0000" when x"77B9",
			x"0000" when x"77BA",
			x"0000" when x"77BB",
			x"0000" when x"77BC",
			x"0000" when x"77BD",
			x"0000" when x"77BE",
			x"0000" when x"77BF",
			x"0000" when x"77C0",
			x"0000" when x"77C1",
			x"0000" when x"77C2",
			x"0000" when x"77C3",
			x"0000" when x"77C4",
			x"0000" when x"77C5",
			x"0000" when x"77C6",
			x"0000" when x"77C7",
			x"0000" when x"77C8",
			x"0000" when x"77C9",
			x"0000" when x"77CA",
			x"0000" when x"77CB",
			x"0000" when x"77CC",
			x"0000" when x"77CD",
			x"0000" when x"77CE",
			x"0000" when x"77CF",
			x"0000" when x"77D0",
			x"0000" when x"77D1",
			x"0000" when x"77D2",
			x"0000" when x"77D3",
			x"0000" when x"77D4",
			x"0000" when x"77D5",
			x"0000" when x"77D6",
			x"0000" when x"77D7",
			x"0000" when x"77D8",
			x"0000" when x"77D9",
			x"0000" when x"77DA",
			x"0000" when x"77DB",
			x"0000" when x"77DC",
			x"0000" when x"77DD",
			x"0000" when x"77DE",
			x"0000" when x"77DF",
			x"0000" when x"77E0",
			x"0000" when x"77E1",
			x"0000" when x"77E2",
			x"0000" when x"77E3",
			x"0000" when x"77E4",
			x"0000" when x"77E5",
			x"0000" when x"77E6",
			x"0000" when x"77E7",
			x"0000" when x"77E8",
			x"0000" when x"77E9",
			x"0000" when x"77EA",
			x"0000" when x"77EB",
			x"0000" when x"77EC",
			x"0000" when x"77ED",
			x"0000" when x"77EE",
			x"0000" when x"77EF",
			x"0000" when x"77F0",
			x"0000" when x"77F1",
			x"0000" when x"77F2",
			x"0000" when x"77F3",
			x"0000" when x"77F4",
			x"0000" when x"77F5",
			x"0000" when x"77F6",
			x"0000" when x"77F7",
			x"0000" when x"77F8",
			x"0000" when x"77F9",
			x"0000" when x"77FA",
			x"0000" when x"77FB",
			x"0000" when x"77FC",
			x"0000" when x"77FD",
			x"0000" when x"77FE",
			x"0000" when x"77FF",
			x"0000" when x"7800",
			x"0000" when x"7801",
			x"0000" when x"7802",
			x"0000" when x"7803",
			x"0000" when x"7804",
			x"0000" when x"7805",
			x"0000" when x"7806",
			x"0000" when x"7807",
			x"0000" when x"7808",
			x"0000" when x"7809",
			x"0000" when x"780A",
			x"0000" when x"780B",
			x"0000" when x"780C",
			x"0000" when x"780D",
			x"0000" when x"780E",
			x"0000" when x"780F",
			x"0000" when x"7810",
			x"0000" when x"7811",
			x"0000" when x"7812",
			x"0000" when x"7813",
			x"0000" when x"7814",
			x"0000" when x"7815",
			x"0000" when x"7816",
			x"0000" when x"7817",
			x"0000" when x"7818",
			x"0000" when x"7819",
			x"0000" when x"781A",
			x"0000" when x"781B",
			x"0000" when x"781C",
			x"0000" when x"781D",
			x"0000" when x"781E",
			x"0000" when x"781F",
			x"0000" when x"7820",
			x"0000" when x"7821",
			x"0000" when x"7822",
			x"0000" when x"7823",
			x"0000" when x"7824",
			x"0000" when x"7825",
			x"0000" when x"7826",
			x"0000" when x"7827",
			x"0000" when x"7828",
			x"0000" when x"7829",
			x"0000" when x"782A",
			x"0000" when x"782B",
			x"0000" when x"782C",
			x"0000" when x"782D",
			x"0000" when x"782E",
			x"0000" when x"782F",
			x"0000" when x"7830",
			x"0000" when x"7831",
			x"0000" when x"7832",
			x"0000" when x"7833",
			x"0000" when x"7834",
			x"0000" when x"7835",
			x"0000" when x"7836",
			x"0000" when x"7837",
			x"0000" when x"7838",
			x"0000" when x"7839",
			x"0000" when x"783A",
			x"0000" when x"783B",
			x"0000" when x"783C",
			x"0000" when x"783D",
			x"0000" when x"783E",
			x"0000" when x"783F",
			x"0000" when x"7840",
			x"0000" when x"7841",
			x"0000" when x"7842",
			x"0000" when x"7843",
			x"0000" when x"7844",
			x"0000" when x"7845",
			x"0000" when x"7846",
			x"0000" when x"7847",
			x"0000" when x"7848",
			x"0000" when x"7849",
			x"0000" when x"784A",
			x"0000" when x"784B",
			x"0000" when x"784C",
			x"0000" when x"784D",
			x"0000" when x"784E",
			x"0000" when x"784F",
			x"0000" when x"7850",
			x"0000" when x"7851",
			x"0000" when x"7852",
			x"0000" when x"7853",
			x"0000" when x"7854",
			x"0000" when x"7855",
			x"0000" when x"7856",
			x"0000" when x"7857",
			x"0000" when x"7858",
			x"0000" when x"7859",
			x"0000" when x"785A",
			x"0000" when x"785B",
			x"0000" when x"785C",
			x"0000" when x"785D",
			x"0000" when x"785E",
			x"0000" when x"785F",
			x"0000" when x"7860",
			x"0000" when x"7861",
			x"0000" when x"7862",
			x"0000" when x"7863",
			x"0000" when x"7864",
			x"0000" when x"7865",
			x"0000" when x"7866",
			x"0000" when x"7867",
			x"0000" when x"7868",
			x"0000" when x"7869",
			x"0000" when x"786A",
			x"0000" when x"786B",
			x"0000" when x"786C",
			x"0000" when x"786D",
			x"0000" when x"786E",
			x"0000" when x"786F",
			x"0000" when x"7870",
			x"0000" when x"7871",
			x"0000" when x"7872",
			x"0000" when x"7873",
			x"0000" when x"7874",
			x"0000" when x"7875",
			x"0000" when x"7876",
			x"0000" when x"7877",
			x"0000" when x"7878",
			x"0000" when x"7879",
			x"0000" when x"787A",
			x"0000" when x"787B",
			x"0000" when x"787C",
			x"0000" when x"787D",
			x"0000" when x"787E",
			x"0000" when x"787F",
			x"0000" when x"7880",
			x"0000" when x"7881",
			x"0000" when x"7882",
			x"0000" when x"7883",
			x"0000" when x"7884",
			x"0000" when x"7885",
			x"0000" when x"7886",
			x"0000" when x"7887",
			x"0000" when x"7888",
			x"0000" when x"7889",
			x"0000" when x"788A",
			x"0000" when x"788B",
			x"0000" when x"788C",
			x"0000" when x"788D",
			x"0000" when x"788E",
			x"0000" when x"788F",
			x"0000" when x"7890",
			x"0000" when x"7891",
			x"0000" when x"7892",
			x"0000" when x"7893",
			x"0000" when x"7894",
			x"0000" when x"7895",
			x"0000" when x"7896",
			x"0000" when x"7897",
			x"0000" when x"7898",
			x"0000" when x"7899",
			x"0000" when x"789A",
			x"0000" when x"789B",
			x"0000" when x"789C",
			x"0000" when x"789D",
			x"0000" when x"789E",
			x"0000" when x"789F",
			x"0000" when x"78A0",
			x"0000" when x"78A1",
			x"0000" when x"78A2",
			x"0000" when x"78A3",
			x"0000" when x"78A4",
			x"0000" when x"78A5",
			x"0000" when x"78A6",
			x"0000" when x"78A7",
			x"0000" when x"78A8",
			x"0000" when x"78A9",
			x"0000" when x"78AA",
			x"0000" when x"78AB",
			x"0000" when x"78AC",
			x"0000" when x"78AD",
			x"0000" when x"78AE",
			x"0000" when x"78AF",
			x"0000" when x"78B0",
			x"0000" when x"78B1",
			x"0000" when x"78B2",
			x"0000" when x"78B3",
			x"0000" when x"78B4",
			x"0000" when x"78B5",
			x"0000" when x"78B6",
			x"0000" when x"78B7",
			x"0000" when x"78B8",
			x"0000" when x"78B9",
			x"0000" when x"78BA",
			x"0000" when x"78BB",
			x"0000" when x"78BC",
			x"0000" when x"78BD",
			x"0000" when x"78BE",
			x"0000" when x"78BF",
			x"0000" when x"78C0",
			x"0000" when x"78C1",
			x"0000" when x"78C2",
			x"0000" when x"78C3",
			x"0000" when x"78C4",
			x"0000" when x"78C5",
			x"0000" when x"78C6",
			x"0000" when x"78C7",
			x"0000" when x"78C8",
			x"0000" when x"78C9",
			x"0000" when x"78CA",
			x"0000" when x"78CB",
			x"0000" when x"78CC",
			x"0000" when x"78CD",
			x"0000" when x"78CE",
			x"0000" when x"78CF",
			x"0000" when x"78D0",
			x"0000" when x"78D1",
			x"0000" when x"78D2",
			x"0000" when x"78D3",
			x"0000" when x"78D4",
			x"0000" when x"78D5",
			x"0000" when x"78D6",
			x"0000" when x"78D7",
			x"0000" when x"78D8",
			x"0000" when x"78D9",
			x"0000" when x"78DA",
			x"0000" when x"78DB",
			x"0000" when x"78DC",
			x"0000" when x"78DD",
			x"0000" when x"78DE",
			x"0000" when x"78DF",
			x"0000" when x"78E0",
			x"0000" when x"78E1",
			x"0000" when x"78E2",
			x"0000" when x"78E3",
			x"0000" when x"78E4",
			x"0000" when x"78E5",
			x"0000" when x"78E6",
			x"0000" when x"78E7",
			x"0000" when x"78E8",
			x"0000" when x"78E9",
			x"0000" when x"78EA",
			x"0000" when x"78EB",
			x"0000" when x"78EC",
			x"0000" when x"78ED",
			x"0000" when x"78EE",
			x"0000" when x"78EF",
			x"0000" when x"78F0",
			x"0000" when x"78F1",
			x"0000" when x"78F2",
			x"0000" when x"78F3",
			x"0000" when x"78F4",
			x"0000" when x"78F5",
			x"0000" when x"78F6",
			x"0000" when x"78F7",
			x"0000" when x"78F8",
			x"0000" when x"78F9",
			x"0000" when x"78FA",
			x"0000" when x"78FB",
			x"0000" when x"78FC",
			x"0000" when x"78FD",
			x"0000" when x"78FE",
			x"0000" when x"78FF",
			x"0000" when x"7900",
			x"0000" when x"7901",
			x"0000" when x"7902",
			x"0000" when x"7903",
			x"0000" when x"7904",
			x"0000" when x"7905",
			x"0000" when x"7906",
			x"0000" when x"7907",
			x"0000" when x"7908",
			x"0000" when x"7909",
			x"0000" when x"790A",
			x"0000" when x"790B",
			x"0000" when x"790C",
			x"0000" when x"790D",
			x"0000" when x"790E",
			x"0000" when x"790F",
			x"0000" when x"7910",
			x"0000" when x"7911",
			x"0000" when x"7912",
			x"0000" when x"7913",
			x"0000" when x"7914",
			x"0000" when x"7915",
			x"0000" when x"7916",
			x"0000" when x"7917",
			x"0000" when x"7918",
			x"0000" when x"7919",
			x"0000" when x"791A",
			x"0000" when x"791B",
			x"0000" when x"791C",
			x"0000" when x"791D",
			x"0000" when x"791E",
			x"0000" when x"791F",
			x"0000" when x"7920",
			x"0000" when x"7921",
			x"0000" when x"7922",
			x"0000" when x"7923",
			x"0000" when x"7924",
			x"0000" when x"7925",
			x"0000" when x"7926",
			x"0000" when x"7927",
			x"0000" when x"7928",
			x"0000" when x"7929",
			x"0000" when x"792A",
			x"0000" when x"792B",
			x"0000" when x"792C",
			x"0000" when x"792D",
			x"0000" when x"792E",
			x"0000" when x"792F",
			x"0000" when x"7930",
			x"0000" when x"7931",
			x"0000" when x"7932",
			x"0000" when x"7933",
			x"0000" when x"7934",
			x"0000" when x"7935",
			x"0000" when x"7936",
			x"0000" when x"7937",
			x"0000" when x"7938",
			x"0000" when x"7939",
			x"0000" when x"793A",
			x"0000" when x"793B",
			x"0000" when x"793C",
			x"0000" when x"793D",
			x"0000" when x"793E",
			x"0000" when x"793F",
			x"0000" when x"7940",
			x"0000" when x"7941",
			x"0000" when x"7942",
			x"0000" when x"7943",
			x"0000" when x"7944",
			x"0000" when x"7945",
			x"0000" when x"7946",
			x"0000" when x"7947",
			x"0000" when x"7948",
			x"0000" when x"7949",
			x"0000" when x"794A",
			x"0000" when x"794B",
			x"0000" when x"794C",
			x"0000" when x"794D",
			x"0000" when x"794E",
			x"0000" when x"794F",
			x"0000" when x"7950",
			x"0000" when x"7951",
			x"0000" when x"7952",
			x"0000" when x"7953",
			x"0000" when x"7954",
			x"0000" when x"7955",
			x"0000" when x"7956",
			x"0000" when x"7957",
			x"0000" when x"7958",
			x"0000" when x"7959",
			x"0000" when x"795A",
			x"0000" when x"795B",
			x"0000" when x"795C",
			x"0000" when x"795D",
			x"0000" when x"795E",
			x"0000" when x"795F",
			x"0000" when x"7960",
			x"0000" when x"7961",
			x"0000" when x"7962",
			x"0000" when x"7963",
			x"0000" when x"7964",
			x"0000" when x"7965",
			x"0000" when x"7966",
			x"0000" when x"7967",
			x"0000" when x"7968",
			x"0000" when x"7969",
			x"0000" when x"796A",
			x"0000" when x"796B",
			x"0000" when x"796C",
			x"0000" when x"796D",
			x"0000" when x"796E",
			x"0000" when x"796F",
			x"0000" when x"7970",
			x"0000" when x"7971",
			x"0000" when x"7972",
			x"0000" when x"7973",
			x"0000" when x"7974",
			x"0000" when x"7975",
			x"0000" when x"7976",
			x"0000" when x"7977",
			x"0000" when x"7978",
			x"0000" when x"7979",
			x"0000" when x"797A",
			x"0000" when x"797B",
			x"0000" when x"797C",
			x"0000" when x"797D",
			x"0000" when x"797E",
			x"0000" when x"797F",
			x"0000" when x"7980",
			x"0000" when x"7981",
			x"0000" when x"7982",
			x"0000" when x"7983",
			x"0000" when x"7984",
			x"0000" when x"7985",
			x"0000" when x"7986",
			x"0000" when x"7987",
			x"0000" when x"7988",
			x"0000" when x"7989",
			x"0000" when x"798A",
			x"0000" when x"798B",
			x"0000" when x"798C",
			x"0000" when x"798D",
			x"0000" when x"798E",
			x"0000" when x"798F",
			x"0000" when x"7990",
			x"0000" when x"7991",
			x"0000" when x"7992",
			x"0000" when x"7993",
			x"0000" when x"7994",
			x"0000" when x"7995",
			x"0000" when x"7996",
			x"0000" when x"7997",
			x"0000" when x"7998",
			x"0000" when x"7999",
			x"0000" when x"799A",
			x"0000" when x"799B",
			x"0000" when x"799C",
			x"0000" when x"799D",
			x"0000" when x"799E",
			x"0000" when x"799F",
			x"0000" when x"79A0",
			x"0000" when x"79A1",
			x"0000" when x"79A2",
			x"0000" when x"79A3",
			x"0000" when x"79A4",
			x"0000" when x"79A5",
			x"0000" when x"79A6",
			x"0000" when x"79A7",
			x"0000" when x"79A8",
			x"0000" when x"79A9",
			x"0000" when x"79AA",
			x"0000" when x"79AB",
			x"0000" when x"79AC",
			x"0000" when x"79AD",
			x"0000" when x"79AE",
			x"0000" when x"79AF",
			x"0000" when x"79B0",
			x"0000" when x"79B1",
			x"0000" when x"79B2",
			x"0000" when x"79B3",
			x"0000" when x"79B4",
			x"0000" when x"79B5",
			x"0000" when x"79B6",
			x"0000" when x"79B7",
			x"0000" when x"79B8",
			x"0000" when x"79B9",
			x"0000" when x"79BA",
			x"0000" when x"79BB",
			x"0000" when x"79BC",
			x"0000" when x"79BD",
			x"0000" when x"79BE",
			x"0000" when x"79BF",
			x"0000" when x"79C0",
			x"0000" when x"79C1",
			x"0000" when x"79C2",
			x"0000" when x"79C3",
			x"0000" when x"79C4",
			x"0000" when x"79C5",
			x"0000" when x"79C6",
			x"0000" when x"79C7",
			x"0000" when x"79C8",
			x"0000" when x"79C9",
			x"0000" when x"79CA",
			x"0000" when x"79CB",
			x"0000" when x"79CC",
			x"0000" when x"79CD",
			x"0000" when x"79CE",
			x"0000" when x"79CF",
			x"0000" when x"79D0",
			x"0000" when x"79D1",
			x"0000" when x"79D2",
			x"0000" when x"79D3",
			x"0000" when x"79D4",
			x"0000" when x"79D5",
			x"0000" when x"79D6",
			x"0000" when x"79D7",
			x"0000" when x"79D8",
			x"0000" when x"79D9",
			x"0000" when x"79DA",
			x"0000" when x"79DB",
			x"0000" when x"79DC",
			x"0000" when x"79DD",
			x"0000" when x"79DE",
			x"0000" when x"79DF",
			x"0000" when x"79E0",
			x"0000" when x"79E1",
			x"0000" when x"79E2",
			x"0000" when x"79E3",
			x"0000" when x"79E4",
			x"0000" when x"79E5",
			x"0000" when x"79E6",
			x"0000" when x"79E7",
			x"0000" when x"79E8",
			x"0000" when x"79E9",
			x"0000" when x"79EA",
			x"0000" when x"79EB",
			x"0000" when x"79EC",
			x"0000" when x"79ED",
			x"0000" when x"79EE",
			x"0000" when x"79EF",
			x"0000" when x"79F0",
			x"0000" when x"79F1",
			x"0000" when x"79F2",
			x"0000" when x"79F3",
			x"0000" when x"79F4",
			x"0000" when x"79F5",
			x"0000" when x"79F6",
			x"0000" when x"79F7",
			x"0000" when x"79F8",
			x"0000" when x"79F9",
			x"0000" when x"79FA",
			x"0000" when x"79FB",
			x"0000" when x"79FC",
			x"0000" when x"79FD",
			x"0000" when x"79FE",
			x"0000" when x"79FF",
			x"0000" when x"7A00",
			x"0000" when x"7A01",
			x"0000" when x"7A02",
			x"0000" when x"7A03",
			x"0000" when x"7A04",
			x"0000" when x"7A05",
			x"0000" when x"7A06",
			x"0000" when x"7A07",
			x"0000" when x"7A08",
			x"0000" when x"7A09",
			x"0000" when x"7A0A",
			x"0000" when x"7A0B",
			x"0000" when x"7A0C",
			x"0000" when x"7A0D",
			x"0000" when x"7A0E",
			x"0000" when x"7A0F",
			x"0000" when x"7A10",
			x"0000" when x"7A11",
			x"0000" when x"7A12",
			x"0000" when x"7A13",
			x"0000" when x"7A14",
			x"0000" when x"7A15",
			x"0000" when x"7A16",
			x"0000" when x"7A17",
			x"0000" when x"7A18",
			x"0000" when x"7A19",
			x"0000" when x"7A1A",
			x"0000" when x"7A1B",
			x"0000" when x"7A1C",
			x"0000" when x"7A1D",
			x"0000" when x"7A1E",
			x"0000" when x"7A1F",
			x"0000" when x"7A20",
			x"0000" when x"7A21",
			x"0000" when x"7A22",
			x"0000" when x"7A23",
			x"0000" when x"7A24",
			x"0000" when x"7A25",
			x"0000" when x"7A26",
			x"0000" when x"7A27",
			x"0000" when x"7A28",
			x"0000" when x"7A29",
			x"0000" when x"7A2A",
			x"0000" when x"7A2B",
			x"0000" when x"7A2C",
			x"0000" when x"7A2D",
			x"0000" when x"7A2E",
			x"0000" when x"7A2F",
			x"0000" when x"7A30",
			x"0000" when x"7A31",
			x"0000" when x"7A32",
			x"0000" when x"7A33",
			x"0000" when x"7A34",
			x"0000" when x"7A35",
			x"0000" when x"7A36",
			x"0000" when x"7A37",
			x"0000" when x"7A38",
			x"0000" when x"7A39",
			x"0000" when x"7A3A",
			x"0000" when x"7A3B",
			x"0000" when x"7A3C",
			x"0000" when x"7A3D",
			x"0000" when x"7A3E",
			x"0000" when x"7A3F",
			x"0000" when x"7A40",
			x"0000" when x"7A41",
			x"0000" when x"7A42",
			x"0000" when x"7A43",
			x"0000" when x"7A44",
			x"0000" when x"7A45",
			x"0000" when x"7A46",
			x"0000" when x"7A47",
			x"0000" when x"7A48",
			x"0000" when x"7A49",
			x"0000" when x"7A4A",
			x"0000" when x"7A4B",
			x"0000" when x"7A4C",
			x"0000" when x"7A4D",
			x"0000" when x"7A4E",
			x"0000" when x"7A4F",
			x"0000" when x"7A50",
			x"0000" when x"7A51",
			x"0000" when x"7A52",
			x"0000" when x"7A53",
			x"0000" when x"7A54",
			x"0000" when x"7A55",
			x"0000" when x"7A56",
			x"0000" when x"7A57",
			x"0000" when x"7A58",
			x"0000" when x"7A59",
			x"0000" when x"7A5A",
			x"0000" when x"7A5B",
			x"0000" when x"7A5C",
			x"0000" when x"7A5D",
			x"0000" when x"7A5E",
			x"0000" when x"7A5F",
			x"0000" when x"7A60",
			x"0000" when x"7A61",
			x"0000" when x"7A62",
			x"0000" when x"7A63",
			x"0000" when x"7A64",
			x"0000" when x"7A65",
			x"0000" when x"7A66",
			x"0000" when x"7A67",
			x"0000" when x"7A68",
			x"0000" when x"7A69",
			x"0000" when x"7A6A",
			x"0000" when x"7A6B",
			x"0000" when x"7A6C",
			x"0000" when x"7A6D",
			x"0000" when x"7A6E",
			x"0000" when x"7A6F",
			x"0000" when x"7A70",
			x"0000" when x"7A71",
			x"0000" when x"7A72",
			x"0000" when x"7A73",
			x"0000" when x"7A74",
			x"0000" when x"7A75",
			x"0000" when x"7A76",
			x"0000" when x"7A77",
			x"0000" when x"7A78",
			x"0000" when x"7A79",
			x"0000" when x"7A7A",
			x"0000" when x"7A7B",
			x"0000" when x"7A7C",
			x"0000" when x"7A7D",
			x"0000" when x"7A7E",
			x"0000" when x"7A7F",
			x"0000" when x"7A80",
			x"0000" when x"7A81",
			x"0000" when x"7A82",
			x"0000" when x"7A83",
			x"0000" when x"7A84",
			x"0000" when x"7A85",
			x"0000" when x"7A86",
			x"0000" when x"7A87",
			x"0000" when x"7A88",
			x"0000" when x"7A89",
			x"0000" when x"7A8A",
			x"0000" when x"7A8B",
			x"0000" when x"7A8C",
			x"0000" when x"7A8D",
			x"0000" when x"7A8E",
			x"0000" when x"7A8F",
			x"0000" when x"7A90",
			x"0000" when x"7A91",
			x"0000" when x"7A92",
			x"0000" when x"7A93",
			x"0000" when x"7A94",
			x"0000" when x"7A95",
			x"0000" when x"7A96",
			x"0000" when x"7A97",
			x"0000" when x"7A98",
			x"0000" when x"7A99",
			x"0000" when x"7A9A",
			x"0000" when x"7A9B",
			x"0000" when x"7A9C",
			x"0000" when x"7A9D",
			x"0000" when x"7A9E",
			x"0000" when x"7A9F",
			x"0000" when x"7AA0",
			x"0000" when x"7AA1",
			x"0000" when x"7AA2",
			x"0000" when x"7AA3",
			x"0000" when x"7AA4",
			x"0000" when x"7AA5",
			x"0000" when x"7AA6",
			x"0000" when x"7AA7",
			x"0000" when x"7AA8",
			x"0000" when x"7AA9",
			x"0000" when x"7AAA",
			x"0000" when x"7AAB",
			x"0000" when x"7AAC",
			x"0000" when x"7AAD",
			x"0000" when x"7AAE",
			x"0000" when x"7AAF",
			x"0000" when x"7AB0",
			x"0000" when x"7AB1",
			x"0000" when x"7AB2",
			x"0000" when x"7AB3",
			x"0000" when x"7AB4",
			x"0000" when x"7AB5",
			x"0000" when x"7AB6",
			x"0000" when x"7AB7",
			x"0000" when x"7AB8",
			x"0000" when x"7AB9",
			x"0000" when x"7ABA",
			x"0000" when x"7ABB",
			x"0000" when x"7ABC",
			x"0000" when x"7ABD",
			x"0000" when x"7ABE",
			x"0000" when x"7ABF",
			x"0000" when x"7AC0",
			x"0000" when x"7AC1",
			x"0000" when x"7AC2",
			x"0000" when x"7AC3",
			x"0000" when x"7AC4",
			x"0000" when x"7AC5",
			x"0000" when x"7AC6",
			x"0000" when x"7AC7",
			x"0000" when x"7AC8",
			x"0000" when x"7AC9",
			x"0000" when x"7ACA",
			x"0000" when x"7ACB",
			x"0000" when x"7ACC",
			x"0000" when x"7ACD",
			x"0000" when x"7ACE",
			x"0000" when x"7ACF",
			x"0000" when x"7AD0",
			x"0000" when x"7AD1",
			x"0000" when x"7AD2",
			x"0000" when x"7AD3",
			x"0000" when x"7AD4",
			x"0000" when x"7AD5",
			x"0000" when x"7AD6",
			x"0000" when x"7AD7",
			x"0000" when x"7AD8",
			x"0000" when x"7AD9",
			x"0000" when x"7ADA",
			x"0000" when x"7ADB",
			x"0000" when x"7ADC",
			x"0000" when x"7ADD",
			x"0000" when x"7ADE",
			x"0000" when x"7ADF",
			x"0000" when x"7AE0",
			x"0000" when x"7AE1",
			x"0000" when x"7AE2",
			x"0000" when x"7AE3",
			x"0000" when x"7AE4",
			x"0000" when x"7AE5",
			x"0000" when x"7AE6",
			x"0000" when x"7AE7",
			x"0000" when x"7AE8",
			x"0000" when x"7AE9",
			x"0000" when x"7AEA",
			x"0000" when x"7AEB",
			x"0000" when x"7AEC",
			x"0000" when x"7AED",
			x"0000" when x"7AEE",
			x"0000" when x"7AEF",
			x"0000" when x"7AF0",
			x"0000" when x"7AF1",
			x"0000" when x"7AF2",
			x"0000" when x"7AF3",
			x"0000" when x"7AF4",
			x"0000" when x"7AF5",
			x"0000" when x"7AF6",
			x"0000" when x"7AF7",
			x"0000" when x"7AF8",
			x"0000" when x"7AF9",
			x"0000" when x"7AFA",
			x"0000" when x"7AFB",
			x"0000" when x"7AFC",
			x"0000" when x"7AFD",
			x"0000" when x"7AFE",
			x"0000" when x"7AFF",
			x"0000" when x"7B00",
			x"0000" when x"7B01",
			x"0000" when x"7B02",
			x"0000" when x"7B03",
			x"0000" when x"7B04",
			x"0000" when x"7B05",
			x"0000" when x"7B06",
			x"0000" when x"7B07",
			x"0000" when x"7B08",
			x"0000" when x"7B09",
			x"0000" when x"7B0A",
			x"0000" when x"7B0B",
			x"0000" when x"7B0C",
			x"0000" when x"7B0D",
			x"0000" when x"7B0E",
			x"0000" when x"7B0F",
			x"0000" when x"7B10",
			x"0000" when x"7B11",
			x"0000" when x"7B12",
			x"0000" when x"7B13",
			x"0000" when x"7B14",
			x"0000" when x"7B15",
			x"0000" when x"7B16",
			x"0000" when x"7B17",
			x"0000" when x"7B18",
			x"0000" when x"7B19",
			x"0000" when x"7B1A",
			x"0000" when x"7B1B",
			x"0000" when x"7B1C",
			x"0000" when x"7B1D",
			x"0000" when x"7B1E",
			x"0000" when x"7B1F",
			x"0000" when x"7B20",
			x"0000" when x"7B21",
			x"0000" when x"7B22",
			x"0000" when x"7B23",
			x"0000" when x"7B24",
			x"0000" when x"7B25",
			x"0000" when x"7B26",
			x"0000" when x"7B27",
			x"0000" when x"7B28",
			x"0000" when x"7B29",
			x"0000" when x"7B2A",
			x"0000" when x"7B2B",
			x"0000" when x"7B2C",
			x"0000" when x"7B2D",
			x"0000" when x"7B2E",
			x"0000" when x"7B2F",
			x"0000" when x"7B30",
			x"0000" when x"7B31",
			x"0000" when x"7B32",
			x"0000" when x"7B33",
			x"0000" when x"7B34",
			x"0000" when x"7B35",
			x"0000" when x"7B36",
			x"0000" when x"7B37",
			x"0000" when x"7B38",
			x"0000" when x"7B39",
			x"0000" when x"7B3A",
			x"0000" when x"7B3B",
			x"0000" when x"7B3C",
			x"0000" when x"7B3D",
			x"0000" when x"7B3E",
			x"0000" when x"7B3F",
			x"0000" when x"7B40",
			x"0000" when x"7B41",
			x"0000" when x"7B42",
			x"0000" when x"7B43",
			x"0000" when x"7B44",
			x"0000" when x"7B45",
			x"0000" when x"7B46",
			x"0000" when x"7B47",
			x"0000" when x"7B48",
			x"0000" when x"7B49",
			x"0000" when x"7B4A",
			x"0000" when x"7B4B",
			x"0000" when x"7B4C",
			x"0000" when x"7B4D",
			x"0000" when x"7B4E",
			x"0000" when x"7B4F",
			x"0000" when x"7B50",
			x"0000" when x"7B51",
			x"0000" when x"7B52",
			x"0000" when x"7B53",
			x"0000" when x"7B54",
			x"0000" when x"7B55",
			x"0000" when x"7B56",
			x"0000" when x"7B57",
			x"0000" when x"7B58",
			x"0000" when x"7B59",
			x"0000" when x"7B5A",
			x"0000" when x"7B5B",
			x"0000" when x"7B5C",
			x"0000" when x"7B5D",
			x"0000" when x"7B5E",
			x"0000" when x"7B5F",
			x"0000" when x"7B60",
			x"0000" when x"7B61",
			x"0000" when x"7B62",
			x"0000" when x"7B63",
			x"0000" when x"7B64",
			x"0000" when x"7B65",
			x"0000" when x"7B66",
			x"0000" when x"7B67",
			x"0000" when x"7B68",
			x"0000" when x"7B69",
			x"0000" when x"7B6A",
			x"0000" when x"7B6B",
			x"0000" when x"7B6C",
			x"0000" when x"7B6D",
			x"0000" when x"7B6E",
			x"0000" when x"7B6F",
			x"0000" when x"7B70",
			x"0000" when x"7B71",
			x"0000" when x"7B72",
			x"0000" when x"7B73",
			x"0000" when x"7B74",
			x"0000" when x"7B75",
			x"0000" when x"7B76",
			x"0000" when x"7B77",
			x"0000" when x"7B78",
			x"0000" when x"7B79",
			x"0000" when x"7B7A",
			x"0000" when x"7B7B",
			x"0000" when x"7B7C",
			x"0000" when x"7B7D",
			x"0000" when x"7B7E",
			x"0000" when x"7B7F",
			x"0000" when x"7B80",
			x"0000" when x"7B81",
			x"0000" when x"7B82",
			x"0000" when x"7B83",
			x"0000" when x"7B84",
			x"0000" when x"7B85",
			x"0000" when x"7B86",
			x"0000" when x"7B87",
			x"0000" when x"7B88",
			x"0000" when x"7B89",
			x"0000" when x"7B8A",
			x"0000" when x"7B8B",
			x"0000" when x"7B8C",
			x"0000" when x"7B8D",
			x"0000" when x"7B8E",
			x"0000" when x"7B8F",
			x"0000" when x"7B90",
			x"0000" when x"7B91",
			x"0000" when x"7B92",
			x"0000" when x"7B93",
			x"0000" when x"7B94",
			x"0000" when x"7B95",
			x"0000" when x"7B96",
			x"0000" when x"7B97",
			x"0000" when x"7B98",
			x"0000" when x"7B99",
			x"0000" when x"7B9A",
			x"0000" when x"7B9B",
			x"0000" when x"7B9C",
			x"0000" when x"7B9D",
			x"0000" when x"7B9E",
			x"0000" when x"7B9F",
			x"0000" when x"7BA0",
			x"0000" when x"7BA1",
			x"0000" when x"7BA2",
			x"0000" when x"7BA3",
			x"0000" when x"7BA4",
			x"0000" when x"7BA5",
			x"0000" when x"7BA6",
			x"0000" when x"7BA7",
			x"0000" when x"7BA8",
			x"0000" when x"7BA9",
			x"0000" when x"7BAA",
			x"0000" when x"7BAB",
			x"0000" when x"7BAC",
			x"0000" when x"7BAD",
			x"0000" when x"7BAE",
			x"0000" when x"7BAF",
			x"0000" when x"7BB0",
			x"0000" when x"7BB1",
			x"0000" when x"7BB2",
			x"0000" when x"7BB3",
			x"0000" when x"7BB4",
			x"0000" when x"7BB5",
			x"0000" when x"7BB6",
			x"0000" when x"7BB7",
			x"0000" when x"7BB8",
			x"0000" when x"7BB9",
			x"0000" when x"7BBA",
			x"0000" when x"7BBB",
			x"0000" when x"7BBC",
			x"0000" when x"7BBD",
			x"0000" when x"7BBE",
			x"0000" when x"7BBF",
			x"0000" when x"7BC0",
			x"0000" when x"7BC1",
			x"0000" when x"7BC2",
			x"0000" when x"7BC3",
			x"0000" when x"7BC4",
			x"0000" when x"7BC5",
			x"0000" when x"7BC6",
			x"0000" when x"7BC7",
			x"0000" when x"7BC8",
			x"0000" when x"7BC9",
			x"0000" when x"7BCA",
			x"0000" when x"7BCB",
			x"0000" when x"7BCC",
			x"0000" when x"7BCD",
			x"0000" when x"7BCE",
			x"0000" when x"7BCF",
			x"0000" when x"7BD0",
			x"0000" when x"7BD1",
			x"0000" when x"7BD2",
			x"0000" when x"7BD3",
			x"0000" when x"7BD4",
			x"0000" when x"7BD5",
			x"0000" when x"7BD6",
			x"0000" when x"7BD7",
			x"0000" when x"7BD8",
			x"0000" when x"7BD9",
			x"0000" when x"7BDA",
			x"0000" when x"7BDB",
			x"0000" when x"7BDC",
			x"0000" when x"7BDD",
			x"0000" when x"7BDE",
			x"0000" when x"7BDF",
			x"0000" when x"7BE0",
			x"0000" when x"7BE1",
			x"0000" when x"7BE2",
			x"0000" when x"7BE3",
			x"0000" when x"7BE4",
			x"0000" when x"7BE5",
			x"0000" when x"7BE6",
			x"0000" when x"7BE7",
			x"0000" when x"7BE8",
			x"0000" when x"7BE9",
			x"0000" when x"7BEA",
			x"0000" when x"7BEB",
			x"0000" when x"7BEC",
			x"0000" when x"7BED",
			x"0000" when x"7BEE",
			x"0000" when x"7BEF",
			x"0000" when x"7BF0",
			x"0000" when x"7BF1",
			x"0000" when x"7BF2",
			x"0000" when x"7BF3",
			x"0000" when x"7BF4",
			x"0000" when x"7BF5",
			x"0000" when x"7BF6",
			x"0000" when x"7BF7",
			x"0000" when x"7BF8",
			x"0000" when x"7BF9",
			x"0000" when x"7BFA",
			x"0000" when x"7BFB",
			x"0000" when x"7BFC",
			x"0000" when x"7BFD",
			x"0000" when x"7BFE",
			x"0000" when x"7BFF",
			x"0000" when x"7C00",
			x"0000" when x"7C01",
			x"0000" when x"7C02",
			x"0000" when x"7C03",
			x"0000" when x"7C04",
			x"0000" when x"7C05",
			x"0000" when x"7C06",
			x"0000" when x"7C07",
			x"0000" when x"7C08",
			x"0000" when x"7C09",
			x"0000" when x"7C0A",
			x"0000" when x"7C0B",
			x"0000" when x"7C0C",
			x"0000" when x"7C0D",
			x"0000" when x"7C0E",
			x"0000" when x"7C0F",
			x"0000" when x"7C10",
			x"0000" when x"7C11",
			x"0000" when x"7C12",
			x"0000" when x"7C13",
			x"0000" when x"7C14",
			x"0000" when x"7C15",
			x"0000" when x"7C16",
			x"0000" when x"7C17",
			x"0000" when x"7C18",
			x"0000" when x"7C19",
			x"0000" when x"7C1A",
			x"0000" when x"7C1B",
			x"0000" when x"7C1C",
			x"0000" when x"7C1D",
			x"0000" when x"7C1E",
			x"0000" when x"7C1F",
			x"0000" when x"7C20",
			x"0000" when x"7C21",
			x"0000" when x"7C22",
			x"0000" when x"7C23",
			x"0000" when x"7C24",
			x"0000" when x"7C25",
			x"0000" when x"7C26",
			x"0000" when x"7C27",
			x"0000" when x"7C28",
			x"0000" when x"7C29",
			x"0000" when x"7C2A",
			x"0000" when x"7C2B",
			x"0000" when x"7C2C",
			x"0000" when x"7C2D",
			x"0000" when x"7C2E",
			x"0000" when x"7C2F",
			x"0000" when x"7C30",
			x"0000" when x"7C31",
			x"0000" when x"7C32",
			x"0000" when x"7C33",
			x"0000" when x"7C34",
			x"0000" when x"7C35",
			x"0000" when x"7C36",
			x"0000" when x"7C37",
			x"0000" when x"7C38",
			x"0000" when x"7C39",
			x"0000" when x"7C3A",
			x"0000" when x"7C3B",
			x"0000" when x"7C3C",
			x"0000" when x"7C3D",
			x"0000" when x"7C3E",
			x"0000" when x"7C3F",
			x"0000" when x"7C40",
			x"0000" when x"7C41",
			x"0000" when x"7C42",
			x"0000" when x"7C43",
			x"0000" when x"7C44",
			x"0000" when x"7C45",
			x"0000" when x"7C46",
			x"0000" when x"7C47",
			x"0000" when x"7C48",
			x"0000" when x"7C49",
			x"0000" when x"7C4A",
			x"0000" when x"7C4B",
			x"0000" when x"7C4C",
			x"0000" when x"7C4D",
			x"0000" when x"7C4E",
			x"0000" when x"7C4F",
			x"0000" when x"7C50",
			x"0000" when x"7C51",
			x"0000" when x"7C52",
			x"0000" when x"7C53",
			x"0000" when x"7C54",
			x"0000" when x"7C55",
			x"0000" when x"7C56",
			x"0000" when x"7C57",
			x"0000" when x"7C58",
			x"0000" when x"7C59",
			x"0000" when x"7C5A",
			x"0000" when x"7C5B",
			x"0000" when x"7C5C",
			x"0000" when x"7C5D",
			x"0000" when x"7C5E",
			x"0000" when x"7C5F",
			x"0000" when x"7C60",
			x"0000" when x"7C61",
			x"0000" when x"7C62",
			x"0000" when x"7C63",
			x"0000" when x"7C64",
			x"0000" when x"7C65",
			x"0000" when x"7C66",
			x"0000" when x"7C67",
			x"0000" when x"7C68",
			x"0000" when x"7C69",
			x"0000" when x"7C6A",
			x"0000" when x"7C6B",
			x"0000" when x"7C6C",
			x"0000" when x"7C6D",
			x"0000" when x"7C6E",
			x"0000" when x"7C6F",
			x"0000" when x"7C70",
			x"0000" when x"7C71",
			x"0000" when x"7C72",
			x"0000" when x"7C73",
			x"0000" when x"7C74",
			x"0000" when x"7C75",
			x"0000" when x"7C76",
			x"0000" when x"7C77",
			x"0000" when x"7C78",
			x"0000" when x"7C79",
			x"0000" when x"7C7A",
			x"0000" when x"7C7B",
			x"0000" when x"7C7C",
			x"0000" when x"7C7D",
			x"0000" when x"7C7E",
			x"0000" when x"7C7F",
			x"0000" when x"7C80",
			x"0000" when x"7C81",
			x"0000" when x"7C82",
			x"0000" when x"7C83",
			x"0000" when x"7C84",
			x"0000" when x"7C85",
			x"0000" when x"7C86",
			x"0000" when x"7C87",
			x"0000" when x"7C88",
			x"0000" when x"7C89",
			x"0000" when x"7C8A",
			x"0000" when x"7C8B",
			x"0000" when x"7C8C",
			x"0000" when x"7C8D",
			x"0000" when x"7C8E",
			x"0000" when x"7C8F",
			x"0000" when x"7C90",
			x"0000" when x"7C91",
			x"0000" when x"7C92",
			x"0000" when x"7C93",
			x"0000" when x"7C94",
			x"0000" when x"7C95",
			x"0000" when x"7C96",
			x"0000" when x"7C97",
			x"0000" when x"7C98",
			x"0000" when x"7C99",
			x"0000" when x"7C9A",
			x"0000" when x"7C9B",
			x"0000" when x"7C9C",
			x"0000" when x"7C9D",
			x"0000" when x"7C9E",
			x"0000" when x"7C9F",
			x"0000" when x"7CA0",
			x"0000" when x"7CA1",
			x"0000" when x"7CA2",
			x"0000" when x"7CA3",
			x"0000" when x"7CA4",
			x"0000" when x"7CA5",
			x"0000" when x"7CA6",
			x"0000" when x"7CA7",
			x"0000" when x"7CA8",
			x"0000" when x"7CA9",
			x"0000" when x"7CAA",
			x"0000" when x"7CAB",
			x"0000" when x"7CAC",
			x"0000" when x"7CAD",
			x"0000" when x"7CAE",
			x"0000" when x"7CAF",
			x"0000" when x"7CB0",
			x"0000" when x"7CB1",
			x"0000" when x"7CB2",
			x"0000" when x"7CB3",
			x"0000" when x"7CB4",
			x"0000" when x"7CB5",
			x"0000" when x"7CB6",
			x"0000" when x"7CB7",
			x"0000" when x"7CB8",
			x"0000" when x"7CB9",
			x"0000" when x"7CBA",
			x"0000" when x"7CBB",
			x"0000" when x"7CBC",
			x"0000" when x"7CBD",
			x"0000" when x"7CBE",
			x"0000" when x"7CBF",
			x"0000" when x"7CC0",
			x"0000" when x"7CC1",
			x"0000" when x"7CC2",
			x"0000" when x"7CC3",
			x"0000" when x"7CC4",
			x"0000" when x"7CC5",
			x"0000" when x"7CC6",
			x"0000" when x"7CC7",
			x"0000" when x"7CC8",
			x"0000" when x"7CC9",
			x"0000" when x"7CCA",
			x"0000" when x"7CCB",
			x"0000" when x"7CCC",
			x"0000" when x"7CCD",
			x"0000" when x"7CCE",
			x"0000" when x"7CCF",
			x"0000" when x"7CD0",
			x"0000" when x"7CD1",
			x"0000" when x"7CD2",
			x"0000" when x"7CD3",
			x"0000" when x"7CD4",
			x"0000" when x"7CD5",
			x"0000" when x"7CD6",
			x"0000" when x"7CD7",
			x"0000" when x"7CD8",
			x"0000" when x"7CD9",
			x"0000" when x"7CDA",
			x"0000" when x"7CDB",
			x"0000" when x"7CDC",
			x"0000" when x"7CDD",
			x"0000" when x"7CDE",
			x"0000" when x"7CDF",
			x"0000" when x"7CE0",
			x"0000" when x"7CE1",
			x"0000" when x"7CE2",
			x"0000" when x"7CE3",
			x"0000" when x"7CE4",
			x"0000" when x"7CE5",
			x"0000" when x"7CE6",
			x"0000" when x"7CE7",
			x"0000" when x"7CE8",
			x"0000" when x"7CE9",
			x"0000" when x"7CEA",
			x"0000" when x"7CEB",
			x"0000" when x"7CEC",
			x"0000" when x"7CED",
			x"0000" when x"7CEE",
			x"0000" when x"7CEF",
			x"0000" when x"7CF0",
			x"0000" when x"7CF1",
			x"0000" when x"7CF2",
			x"0000" when x"7CF3",
			x"0000" when x"7CF4",
			x"0000" when x"7CF5",
			x"0000" when x"7CF6",
			x"0000" when x"7CF7",
			x"0000" when x"7CF8",
			x"0000" when x"7CF9",
			x"0000" when x"7CFA",
			x"0000" when x"7CFB",
			x"0000" when x"7CFC",
			x"0000" when x"7CFD",
			x"0000" when x"7CFE",
			x"0000" when x"7CFF",
			x"0000" when x"7D00",
			x"0000" when x"7D01",
			x"0000" when x"7D02",
			x"0000" when x"7D03",
			x"0000" when x"7D04",
			x"0000" when x"7D05",
			x"0000" when x"7D06",
			x"0000" when x"7D07",
			x"0000" when x"7D08",
			x"0000" when x"7D09",
			x"0000" when x"7D0A",
			x"0000" when x"7D0B",
			x"0000" when x"7D0C",
			x"0000" when x"7D0D",
			x"0000" when x"7D0E",
			x"0000" when x"7D0F",
			x"0000" when x"7D10",
			x"0000" when x"7D11",
			x"0000" when x"7D12",
			x"0000" when x"7D13",
			x"0000" when x"7D14",
			x"0000" when x"7D15",
			x"0000" when x"7D16",
			x"0000" when x"7D17",
			x"0000" when x"7D18",
			x"0000" when x"7D19",
			x"0000" when x"7D1A",
			x"0000" when x"7D1B",
			x"0000" when x"7D1C",
			x"0000" when x"7D1D",
			x"0000" when x"7D1E",
			x"0000" when x"7D1F",
			x"0000" when x"7D20",
			x"0000" when x"7D21",
			x"0000" when x"7D22",
			x"0000" when x"7D23",
			x"0000" when x"7D24",
			x"0000" when x"7D25",
			x"0000" when x"7D26",
			x"0000" when x"7D27",
			x"0000" when x"7D28",
			x"0000" when x"7D29",
			x"0000" when x"7D2A",
			x"0000" when x"7D2B",
			x"0000" when x"7D2C",
			x"0000" when x"7D2D",
			x"0000" when x"7D2E",
			x"0000" when x"7D2F",
			x"0000" when x"7D30",
			x"0000" when x"7D31",
			x"0000" when x"7D32",
			x"0000" when x"7D33",
			x"0000" when x"7D34",
			x"0000" when x"7D35",
			x"0000" when x"7D36",
			x"0000" when x"7D37",
			x"0000" when x"7D38",
			x"0000" when x"7D39",
			x"0000" when x"7D3A",
			x"0000" when x"7D3B",
			x"0000" when x"7D3C",
			x"0000" when x"7D3D",
			x"0000" when x"7D3E",
			x"0000" when x"7D3F",
			x"0000" when x"7D40",
			x"0000" when x"7D41",
			x"0000" when x"7D42",
			x"0000" when x"7D43",
			x"0000" when x"7D44",
			x"0000" when x"7D45",
			x"0000" when x"7D46",
			x"0000" when x"7D47",
			x"0000" when x"7D48",
			x"0000" when x"7D49",
			x"0000" when x"7D4A",
			x"0000" when x"7D4B",
			x"0000" when x"7D4C",
			x"0000" when x"7D4D",
			x"0000" when x"7D4E",
			x"0000" when x"7D4F",
			x"0000" when x"7D50",
			x"0000" when x"7D51",
			x"0000" when x"7D52",
			x"0000" when x"7D53",
			x"0000" when x"7D54",
			x"0000" when x"7D55",
			x"0000" when x"7D56",
			x"0000" when x"7D57",
			x"0000" when x"7D58",
			x"0000" when x"7D59",
			x"0000" when x"7D5A",
			x"0000" when x"7D5B",
			x"0000" when x"7D5C",
			x"0000" when x"7D5D",
			x"0000" when x"7D5E",
			x"0000" when x"7D5F",
			x"0000" when x"7D60",
			x"0000" when x"7D61",
			x"0000" when x"7D62",
			x"0000" when x"7D63",
			x"0000" when x"7D64",
			x"0000" when x"7D65",
			x"0000" when x"7D66",
			x"0000" when x"7D67",
			x"0000" when x"7D68",
			x"0000" when x"7D69",
			x"0000" when x"7D6A",
			x"0000" when x"7D6B",
			x"0000" when x"7D6C",
			x"0000" when x"7D6D",
			x"0000" when x"7D6E",
			x"0000" when x"7D6F",
			x"0000" when x"7D70",
			x"0000" when x"7D71",
			x"0000" when x"7D72",
			x"0000" when x"7D73",
			x"0000" when x"7D74",
			x"0000" when x"7D75",
			x"0000" when x"7D76",
			x"0000" when x"7D77",
			x"0000" when x"7D78",
			x"0000" when x"7D79",
			x"0000" when x"7D7A",
			x"0000" when x"7D7B",
			x"0000" when x"7D7C",
			x"0000" when x"7D7D",
			x"0000" when x"7D7E",
			x"0000" when x"7D7F",
			x"0000" when x"7D80",
			x"0000" when x"7D81",
			x"0000" when x"7D82",
			x"0000" when x"7D83",
			x"0000" when x"7D84",
			x"0000" when x"7D85",
			x"0000" when x"7D86",
			x"0000" when x"7D87",
			x"0000" when x"7D88",
			x"0000" when x"7D89",
			x"0000" when x"7D8A",
			x"0000" when x"7D8B",
			x"0000" when x"7D8C",
			x"0000" when x"7D8D",
			x"0000" when x"7D8E",
			x"0000" when x"7D8F",
			x"0000" when x"7D90",
			x"0000" when x"7D91",
			x"0000" when x"7D92",
			x"0000" when x"7D93",
			x"0000" when x"7D94",
			x"0000" when x"7D95",
			x"0000" when x"7D96",
			x"0000" when x"7D97",
			x"0000" when x"7D98",
			x"0000" when x"7D99",
			x"0000" when x"7D9A",
			x"0000" when x"7D9B",
			x"0000" when x"7D9C",
			x"0000" when x"7D9D",
			x"0000" when x"7D9E",
			x"0000" when x"7D9F",
			x"0000" when x"7DA0",
			x"0000" when x"7DA1",
			x"0000" when x"7DA2",
			x"0000" when x"7DA3",
			x"0000" when x"7DA4",
			x"0000" when x"7DA5",
			x"0000" when x"7DA6",
			x"0000" when x"7DA7",
			x"0000" when x"7DA8",
			x"0000" when x"7DA9",
			x"0000" when x"7DAA",
			x"0000" when x"7DAB",
			x"0000" when x"7DAC",
			x"0000" when x"7DAD",
			x"0000" when x"7DAE",
			x"0000" when x"7DAF",
			x"0000" when x"7DB0",
			x"0000" when x"7DB1",
			x"0000" when x"7DB2",
			x"0000" when x"7DB3",
			x"0000" when x"7DB4",
			x"0000" when x"7DB5",
			x"0000" when x"7DB6",
			x"0000" when x"7DB7",
			x"0000" when x"7DB8",
			x"0000" when x"7DB9",
			x"0000" when x"7DBA",
			x"0000" when x"7DBB",
			x"0000" when x"7DBC",
			x"0000" when x"7DBD",
			x"0000" when x"7DBE",
			x"0000" when x"7DBF",
			x"0000" when x"7DC0",
			x"0000" when x"7DC1",
			x"0000" when x"7DC2",
			x"0000" when x"7DC3",
			x"0000" when x"7DC4",
			x"0000" when x"7DC5",
			x"0000" when x"7DC6",
			x"0000" when x"7DC7",
			x"0000" when x"7DC8",
			x"0000" when x"7DC9",
			x"0000" when x"7DCA",
			x"0000" when x"7DCB",
			x"0000" when x"7DCC",
			x"0000" when x"7DCD",
			x"0000" when x"7DCE",
			x"0000" when x"7DCF",
			x"0000" when x"7DD0",
			x"0000" when x"7DD1",
			x"0000" when x"7DD2",
			x"0000" when x"7DD3",
			x"0000" when x"7DD4",
			x"0000" when x"7DD5",
			x"0000" when x"7DD6",
			x"0000" when x"7DD7",
			x"0000" when x"7DD8",
			x"0000" when x"7DD9",
			x"0000" when x"7DDA",
			x"0000" when x"7DDB",
			x"0000" when x"7DDC",
			x"0000" when x"7DDD",
			x"0000" when x"7DDE",
			x"0000" when x"7DDF",
			x"0000" when x"7DE0",
			x"0000" when x"7DE1",
			x"0000" when x"7DE2",
			x"0000" when x"7DE3",
			x"0000" when x"7DE4",
			x"0000" when x"7DE5",
			x"0000" when x"7DE6",
			x"0000" when x"7DE7",
			x"0000" when x"7DE8",
			x"0000" when x"7DE9",
			x"0000" when x"7DEA",
			x"0000" when x"7DEB",
			x"0000" when x"7DEC",
			x"0000" when x"7DED",
			x"0000" when x"7DEE",
			x"0000" when x"7DEF",
			x"0000" when x"7DF0",
			x"0000" when x"7DF1",
			x"0000" when x"7DF2",
			x"0000" when x"7DF3",
			x"0000" when x"7DF4",
			x"0000" when x"7DF5",
			x"0000" when x"7DF6",
			x"0000" when x"7DF7",
			x"0000" when x"7DF8",
			x"0000" when x"7DF9",
			x"0000" when x"7DFA",
			x"0000" when x"7DFB",
			x"0000" when x"7DFC",
			x"0000" when x"7DFD",
			x"0000" when x"7DFE",
			x"0000" when x"7DFF",
			x"0000" when x"7E00",
			x"0000" when x"7E01",
			x"0000" when x"7E02",
			x"0000" when x"7E03",
			x"0000" when x"7E04",
			x"0000" when x"7E05",
			x"0000" when x"7E06",
			x"0000" when x"7E07",
			x"0000" when x"7E08",
			x"0000" when x"7E09",
			x"0000" when x"7E0A",
			x"0000" when x"7E0B",
			x"0000" when x"7E0C",
			x"0000" when x"7E0D",
			x"0000" when x"7E0E",
			x"0000" when x"7E0F",
			x"0000" when x"7E10",
			x"0000" when x"7E11",
			x"0000" when x"7E12",
			x"0000" when x"7E13",
			x"0000" when x"7E14",
			x"0000" when x"7E15",
			x"0000" when x"7E16",
			x"0000" when x"7E17",
			x"0000" when x"7E18",
			x"0000" when x"7E19",
			x"0000" when x"7E1A",
			x"0000" when x"7E1B",
			x"0000" when x"7E1C",
			x"0000" when x"7E1D",
			x"0000" when x"7E1E",
			x"0000" when x"7E1F",
			x"0000" when x"7E20",
			x"0000" when x"7E21",
			x"0000" when x"7E22",
			x"0000" when x"7E23",
			x"0000" when x"7E24",
			x"0000" when x"7E25",
			x"0000" when x"7E26",
			x"0000" when x"7E27",
			x"0000" when x"7E28",
			x"0000" when x"7E29",
			x"0000" when x"7E2A",
			x"0000" when x"7E2B",
			x"0000" when x"7E2C",
			x"0000" when x"7E2D",
			x"0000" when x"7E2E",
			x"0000" when x"7E2F",
			x"0000" when x"7E30",
			x"0000" when x"7E31",
			x"0000" when x"7E32",
			x"0000" when x"7E33",
			x"0000" when x"7E34",
			x"0000" when x"7E35",
			x"0000" when x"7E36",
			x"0000" when x"7E37",
			x"0000" when x"7E38",
			x"0000" when x"7E39",
			x"0000" when x"7E3A",
			x"0000" when x"7E3B",
			x"0000" when x"7E3C",
			x"0000" when x"7E3D",
			x"0000" when x"7E3E",
			x"0000" when x"7E3F",
			x"0000" when x"7E40",
			x"0000" when x"7E41",
			x"0000" when x"7E42",
			x"0000" when x"7E43",
			x"0000" when x"7E44",
			x"0000" when x"7E45",
			x"0000" when x"7E46",
			x"0000" when x"7E47",
			x"0000" when x"7E48",
			x"0000" when x"7E49",
			x"0000" when x"7E4A",
			x"0000" when x"7E4B",
			x"0000" when x"7E4C",
			x"0000" when x"7E4D",
			x"0000" when x"7E4E",
			x"0000" when x"7E4F",
			x"0000" when x"7E50",
			x"0000" when x"7E51",
			x"0000" when x"7E52",
			x"0000" when x"7E53",
			x"0000" when x"7E54",
			x"0000" when x"7E55",
			x"0000" when x"7E56",
			x"0000" when x"7E57",
			x"0000" when x"7E58",
			x"0000" when x"7E59",
			x"0000" when x"7E5A",
			x"0000" when x"7E5B",
			x"0000" when x"7E5C",
			x"0000" when x"7E5D",
			x"0000" when x"7E5E",
			x"0000" when x"7E5F",
			x"0000" when x"7E60",
			x"0000" when x"7E61",
			x"0000" when x"7E62",
			x"0000" when x"7E63",
			x"0000" when x"7E64",
			x"0000" when x"7E65",
			x"0000" when x"7E66",
			x"0000" when x"7E67",
			x"0000" when x"7E68",
			x"0000" when x"7E69",
			x"0000" when x"7E6A",
			x"0000" when x"7E6B",
			x"0000" when x"7E6C",
			x"0000" when x"7E6D",
			x"0000" when x"7E6E",
			x"0000" when x"7E6F",
			x"0000" when x"7E70",
			x"0000" when x"7E71",
			x"0000" when x"7E72",
			x"0000" when x"7E73",
			x"0000" when x"7E74",
			x"0000" when x"7E75",
			x"0000" when x"7E76",
			x"0000" when x"7E77",
			x"0000" when x"7E78",
			x"0000" when x"7E79",
			x"0000" when x"7E7A",
			x"0000" when x"7E7B",
			x"0000" when x"7E7C",
			x"0000" when x"7E7D",
			x"0000" when x"7E7E",
			x"0000" when x"7E7F",
			x"0000" when x"7E80",
			x"0000" when x"7E81",
			x"0000" when x"7E82",
			x"0000" when x"7E83",
			x"0000" when x"7E84",
			x"0000" when x"7E85",
			x"0000" when x"7E86",
			x"0000" when x"7E87",
			x"0000" when x"7E88",
			x"0000" when x"7E89",
			x"0000" when x"7E8A",
			x"0000" when x"7E8B",
			x"0000" when x"7E8C",
			x"0000" when x"7E8D",
			x"0000" when x"7E8E",
			x"0000" when x"7E8F",
			x"0000" when x"7E90",
			x"0000" when x"7E91",
			x"0000" when x"7E92",
			x"0000" when x"7E93",
			x"0000" when x"7E94",
			x"0000" when x"7E95",
			x"0000" when x"7E96",
			x"0000" when x"7E97",
			x"0000" when x"7E98",
			x"0000" when x"7E99",
			x"0000" when x"7E9A",
			x"0000" when x"7E9B",
			x"0000" when x"7E9C",
			x"0000" when x"7E9D",
			x"0000" when x"7E9E",
			x"0000" when x"7E9F",
			x"0000" when x"7EA0",
			x"0000" when x"7EA1",
			x"0000" when x"7EA2",
			x"0000" when x"7EA3",
			x"0000" when x"7EA4",
			x"0000" when x"7EA5",
			x"0000" when x"7EA6",
			x"0000" when x"7EA7",
			x"0000" when x"7EA8",
			x"0000" when x"7EA9",
			x"0000" when x"7EAA",
			x"0000" when x"7EAB",
			x"0000" when x"7EAC",
			x"0000" when x"7EAD",
			x"0000" when x"7EAE",
			x"0000" when x"7EAF",
			x"0000" when x"7EB0",
			x"0000" when x"7EB1",
			x"0000" when x"7EB2",
			x"0000" when x"7EB3",
			x"0000" when x"7EB4",
			x"0000" when x"7EB5",
			x"0000" when x"7EB6",
			x"0000" when x"7EB7",
			x"0000" when x"7EB8",
			x"0000" when x"7EB9",
			x"0000" when x"7EBA",
			x"0000" when x"7EBB",
			x"0000" when x"7EBC",
			x"0000" when x"7EBD",
			x"0000" when x"7EBE",
			x"0000" when x"7EBF",
			x"0000" when x"7EC0",
			x"0000" when x"7EC1",
			x"0000" when x"7EC2",
			x"0000" when x"7EC3",
			x"0000" when x"7EC4",
			x"0000" when x"7EC5",
			x"0000" when x"7EC6",
			x"0000" when x"7EC7",
			x"0000" when x"7EC8",
			x"0000" when x"7EC9",
			x"0000" when x"7ECA",
			x"0000" when x"7ECB",
			x"0000" when x"7ECC",
			x"0000" when x"7ECD",
			x"0000" when x"7ECE",
			x"0000" when x"7ECF",
			x"0000" when x"7ED0",
			x"0000" when x"7ED1",
			x"0000" when x"7ED2",
			x"0000" when x"7ED3",
			x"0000" when x"7ED4",
			x"0000" when x"7ED5",
			x"0000" when x"7ED6",
			x"0000" when x"7ED7",
			x"0000" when x"7ED8",
			x"0000" when x"7ED9",
			x"0000" when x"7EDA",
			x"0000" when x"7EDB",
			x"0000" when x"7EDC",
			x"0000" when x"7EDD",
			x"0000" when x"7EDE",
			x"0000" when x"7EDF",
			x"0000" when x"7EE0",
			x"0000" when x"7EE1",
			x"0000" when x"7EE2",
			x"0000" when x"7EE3",
			x"0000" when x"7EE4",
			x"0000" when x"7EE5",
			x"0000" when x"7EE6",
			x"0000" when x"7EE7",
			x"0000" when x"7EE8",
			x"0000" when x"7EE9",
			x"0000" when x"7EEA",
			x"0000" when x"7EEB",
			x"0000" when x"7EEC",
			x"0000" when x"7EED",
			x"0000" when x"7EEE",
			x"0000" when x"7EEF",
			x"0000" when x"7EF0",
			x"0000" when x"7EF1",
			x"0000" when x"7EF2",
			x"0000" when x"7EF3",
			x"0000" when x"7EF4",
			x"0000" when x"7EF5",
			x"0000" when x"7EF6",
			x"0000" when x"7EF7",
			x"0000" when x"7EF8",
			x"0000" when x"7EF9",
			x"0000" when x"7EFA",
			x"0000" when x"7EFB",
			x"0000" when x"7EFC",
			x"0000" when x"7EFD",
			x"0000" when x"7EFE",
			x"0000" when x"7EFF",
			x"0000" when x"7F00",
			x"0000" when x"7F01",
			x"0000" when x"7F02",
			x"0000" when x"7F03",
			x"0000" when x"7F04",
			x"0000" when x"7F05",
			x"0000" when x"7F06",
			x"0000" when x"7F07",
			x"0000" when x"7F08",
			x"0000" when x"7F09",
			x"0000" when x"7F0A",
			x"0000" when x"7F0B",
			x"0000" when x"7F0C",
			x"0000" when x"7F0D",
			x"0000" when x"7F0E",
			x"0000" when x"7F0F",
			x"0000" when x"7F10",
			x"0000" when x"7F11",
			x"0000" when x"7F12",
			x"0000" when x"7F13",
			x"0000" when x"7F14",
			x"0000" when x"7F15",
			x"0000" when x"7F16",
			x"0000" when x"7F17",
			x"0000" when x"7F18",
			x"0000" when x"7F19",
			x"0000" when x"7F1A",
			x"0000" when x"7F1B",
			x"0000" when x"7F1C",
			x"0000" when x"7F1D",
			x"0000" when x"7F1E",
			x"0000" when x"7F1F",
			x"0000" when x"7F20",
			x"0000" when x"7F21",
			x"0000" when x"7F22",
			x"0000" when x"7F23",
			x"0000" when x"7F24",
			x"0000" when x"7F25",
			x"0000" when x"7F26",
			x"0000" when x"7F27",
			x"0000" when x"7F28",
			x"0000" when x"7F29",
			x"0000" when x"7F2A",
			x"0000" when x"7F2B",
			x"0000" when x"7F2C",
			x"0000" when x"7F2D",
			x"0000" when x"7F2E",
			x"0000" when x"7F2F",
			x"0000" when x"7F30",
			x"0000" when x"7F31",
			x"0000" when x"7F32",
			x"0000" when x"7F33",
			x"0000" when x"7F34",
			x"0000" when x"7F35",
			x"0000" when x"7F36",
			x"0000" when x"7F37",
			x"0000" when x"7F38",
			x"0000" when x"7F39",
			x"0000" when x"7F3A",
			x"0000" when x"7F3B",
			x"0000" when x"7F3C",
			x"0000" when x"7F3D",
			x"0000" when x"7F3E",
			x"0000" when x"7F3F",
			x"0000" when x"7F40",
			x"0000" when x"7F41",
			x"0000" when x"7F42",
			x"0000" when x"7F43",
			x"0000" when x"7F44",
			x"0000" when x"7F45",
			x"0000" when x"7F46",
			x"0000" when x"7F47",
			x"0000" when x"7F48",
			x"0000" when x"7F49",
			x"0000" when x"7F4A",
			x"0000" when x"7F4B",
			x"0000" when x"7F4C",
			x"0000" when x"7F4D",
			x"0000" when x"7F4E",
			x"0000" when x"7F4F",
			x"0000" when x"7F50",
			x"0000" when x"7F51",
			x"0000" when x"7F52",
			x"0000" when x"7F53",
			x"0000" when x"7F54",
			x"0000" when x"7F55",
			x"0000" when x"7F56",
			x"0000" when x"7F57",
			x"0000" when x"7F58",
			x"0000" when x"7F59",
			x"0000" when x"7F5A",
			x"0000" when x"7F5B",
			x"0000" when x"7F5C",
			x"0000" when x"7F5D",
			x"0000" when x"7F5E",
			x"0000" when x"7F5F",
			x"0000" when x"7F60",
			x"0000" when x"7F61",
			x"0000" when x"7F62",
			x"0000" when x"7F63",
			x"0000" when x"7F64",
			x"0000" when x"7F65",
			x"0000" when x"7F66",
			x"0000" when x"7F67",
			x"0000" when x"7F68",
			x"0000" when x"7F69",
			x"0000" when x"7F6A",
			x"0000" when x"7F6B",
			x"0000" when x"7F6C",
			x"0000" when x"7F6D",
			x"0000" when x"7F6E",
			x"0000" when x"7F6F",
			x"0000" when x"7F70",
			x"0000" when x"7F71",
			x"0000" when x"7F72",
			x"0000" when x"7F73",
			x"0000" when x"7F74",
			x"0000" when x"7F75",
			x"0000" when x"7F76",
			x"0000" when x"7F77",
			x"0000" when x"7F78",
			x"0000" when x"7F79",
			x"0000" when x"7F7A",
			x"0000" when x"7F7B",
			x"0000" when x"7F7C",
			x"0000" when x"7F7D",
			x"0000" when x"7F7E",
			x"0000" when x"7F7F",
			x"0000" when x"7F80",
			x"0000" when x"7F81",
			x"0000" when x"7F82",
			x"0000" when x"7F83",
			x"0000" when x"7F84",
			x"0000" when x"7F85",
			x"0000" when x"7F86",
			x"0000" when x"7F87",
			x"0000" when x"7F88",
			x"0000" when x"7F89",
			x"0000" when x"7F8A",
			x"0000" when x"7F8B",
			x"0000" when x"7F8C",
			x"0000" when x"7F8D",
			x"0000" when x"7F8E",
			x"0000" when x"7F8F",
			x"0000" when x"7F90",
			x"0000" when x"7F91",
			x"0000" when x"7F92",
			x"0000" when x"7F93",
			x"0000" when x"7F94",
			x"0000" when x"7F95",
			x"0000" when x"7F96",
			x"0000" when x"7F97",
			x"0000" when x"7F98",
			x"0000" when x"7F99",
			x"0000" when x"7F9A",
			x"0000" when x"7F9B",
			x"0000" when x"7F9C",
			x"0000" when x"7F9D",
			x"0000" when x"7F9E",
			x"0000" when x"7F9F",
			x"0000" when x"7FA0",
			x"0000" when x"7FA1",
			x"0000" when x"7FA2",
			x"0000" when x"7FA3",
			x"0000" when x"7FA4",
			x"0000" when x"7FA5",
			x"0000" when x"7FA6",
			x"0000" when x"7FA7",
			x"0000" when x"7FA8",
			x"0000" when x"7FA9",
			x"0000" when x"7FAA",
			x"0000" when x"7FAB",
			x"0000" when x"7FAC",
			x"0000" when x"7FAD",
			x"0000" when x"7FAE",
			x"0000" when x"7FAF",
			x"0000" when x"7FB0",
			x"0000" when x"7FB1",
			x"0000" when x"7FB2",
			x"0000" when x"7FB3",
			x"0000" when x"7FB4",
			x"0000" when x"7FB5",
			x"0000" when x"7FB6",
			x"0000" when x"7FB7",
			x"0000" when x"7FB8",
			x"0000" when x"7FB9",
			x"0000" when x"7FBA",
			x"0000" when x"7FBB",
			x"0000" when x"7FBC",
			x"0000" when x"7FBD",
			x"0000" when x"7FBE",
			x"0000" when x"7FBF",
			x"0000" when x"7FC0",
			x"0000" when x"7FC1",
			x"0000" when x"7FC2",
			x"0000" when x"7FC3",
			x"0000" when x"7FC4",
			x"0000" when x"7FC5",
			x"0000" when x"7FC6",
			x"0000" when x"7FC7",
			x"0000" when x"7FC8",
			x"0000" when x"7FC9",
			x"0000" when x"7FCA",
			x"0000" when x"7FCB",
			x"0000" when x"7FCC",
			x"0000" when x"7FCD",
			x"0000" when x"7FCE",
			x"0000" when x"7FCF",
			x"0000" when x"7FD0",
			x"0000" when x"7FD1",
			x"0000" when x"7FD2",
			x"0000" when x"7FD3",
			x"0000" when x"7FD4",
			x"0000" when x"7FD5",
			x"0000" when x"7FD6",
			x"0000" when x"7FD7",
			x"0000" when x"7FD8",
			x"0000" when x"7FD9",
			x"0000" when x"7FDA",
			x"0000" when x"7FDB",
			x"0000" when x"7FDC",
			x"0000" when x"7FDD",
			x"0000" when x"7FDE",
			x"0000" when x"7FDF",
			x"0000" when x"7FE0",
			x"0000" when x"7FE1",
			x"0000" when x"7FE2",
			x"0000" when x"7FE3",
			x"0000" when x"7FE4",
			x"0000" when x"7FE5",
			x"0000" when x"7FE6",
			x"0000" when x"7FE7",
			x"0000" when x"7FE8",
			x"0000" when x"7FE9",
			x"0000" when x"7FEA",
			x"0000" when x"7FEB",
			x"0000" when x"7FEC",
			x"0000" when x"7FED",
			x"0000" when x"7FEE",
			x"0000" when x"7FEF",
			x"0000" when x"7FF0",
			x"0000" when x"7FF1",
			x"0000" when x"7FF2",
			x"0000" when x"7FF3",
			x"0000" when x"7FF4",
			x"0000" when x"7FF5",
			x"0000" when x"7FF6",
			x"0000" when x"7FF7",
			x"0000" when x"7FF8",
			x"0000" when x"7FF9",
			x"0000" when x"7FFA",
			x"0000" when x"7FFB",
			x"0000" when x"7FFC",
			x"0000" when x"7FFD",
			x"0000" when x"7FFE",
			x"0000" when x"7FFF",
			x"0000" when x"8000",
			x"0000" when x"8001",
			x"0000" when x"8002",
			x"0000" when x"8003",
			x"0000" when x"8004",
			x"0000" when x"8005",
			x"0000" when x"8006",
			x"0000" when x"8007",
			x"0000" when x"8008",
			x"0000" when x"8009",
			x"0000" when x"800A",
			x"0000" when x"800B",
			x"0000" when x"800C",
			x"0000" when x"800D",
			x"0000" when x"800E",
			x"0000" when x"800F",
			x"0000" when x"8010",
			x"0000" when x"8011",
			x"0000" when x"8012",
			x"0000" when x"8013",
			x"0000" when x"8014",
			x"0000" when x"8015",
			x"0000" when x"8016",
			x"0000" when x"8017",
			x"0000" when x"8018",
			x"0000" when x"8019",
			x"0000" when x"801A",
			x"0000" when x"801B",
			x"0000" when x"801C",
			x"0000" when x"801D",
			x"0000" when x"801E",
			x"0000" when x"801F",
			x"0000" when x"8020",
			x"0000" when x"8021",
			x"0000" when x"8022",
			x"0000" when x"8023",
			x"0000" when x"8024",
			x"0000" when x"8025",
			x"0000" when x"8026",
			x"0000" when x"8027",
			x"0000" when x"8028",
			x"0000" when x"8029",
			x"0000" when x"802A",
			x"0000" when x"802B",
			x"0000" when x"802C",
			x"0000" when x"802D",
			x"0000" when x"802E",
			x"0000" when x"802F",
			x"0000" when x"8030",
			x"0000" when x"8031",
			x"0000" when x"8032",
			x"0000" when x"8033",
			x"0000" when x"8034",
			x"0000" when x"8035",
			x"0000" when x"8036",
			x"0000" when x"8037",
			x"0000" when x"8038",
			x"0000" when x"8039",
			x"0000" when x"803A",
			x"0000" when x"803B",
			x"0000" when x"803C",
			x"0000" when x"803D",
			x"0000" when x"803E",
			x"0000" when x"803F",
			x"0000" when x"8040",
			x"0000" when x"8041",
			x"0000" when x"8042",
			x"0000" when x"8043",
			x"0000" when x"8044",
			x"0000" when x"8045",
			x"0000" when x"8046",
			x"0000" when x"8047",
			x"0000" when x"8048",
			x"0000" when x"8049",
			x"0000" when x"804A",
			x"0000" when x"804B",
			x"0000" when x"804C",
			x"0000" when x"804D",
			x"0000" when x"804E",
			x"0000" when x"804F",
			x"0000" when x"8050",
			x"0000" when x"8051",
			x"0000" when x"8052",
			x"0000" when x"8053",
			x"0000" when x"8054",
			x"0000" when x"8055",
			x"0000" when x"8056",
			x"0000" when x"8057",
			x"0000" when x"8058",
			x"0000" when x"8059",
			x"0000" when x"805A",
			x"0000" when x"805B",
			x"0000" when x"805C",
			x"0000" when x"805D",
			x"0000" when x"805E",
			x"0000" when x"805F",
			x"0000" when x"8060",
			x"0000" when x"8061",
			x"0000" when x"8062",
			x"0000" when x"8063",
			x"0000" when x"8064",
			x"0000" when x"8065",
			x"0000" when x"8066",
			x"0000" when x"8067",
			x"0000" when x"8068",
			x"0000" when x"8069",
			x"0000" when x"806A",
			x"0000" when x"806B",
			x"0000" when x"806C",
			x"0000" when x"806D",
			x"0000" when x"806E",
			x"0000" when x"806F",
			x"0000" when x"8070",
			x"0000" when x"8071",
			x"0000" when x"8072",
			x"0000" when x"8073",
			x"0000" when x"8074",
			x"0000" when x"8075",
			x"0000" when x"8076",
			x"0000" when x"8077",
			x"0000" when x"8078",
			x"0000" when x"8079",
			x"0000" when x"807A",
			x"0000" when x"807B",
			x"0000" when x"807C",
			x"0000" when x"807D",
			x"0000" when x"807E",
			x"0000" when x"807F",
			x"0000" when x"8080",
			x"0000" when x"8081",
			x"0000" when x"8082",
			x"0000" when x"8083",
			x"0000" when x"8084",
			x"0000" when x"8085",
			x"0000" when x"8086",
			x"0000" when x"8087",
			x"0000" when x"8088",
			x"0000" when x"8089",
			x"0000" when x"808A",
			x"0000" when x"808B",
			x"0000" when x"808C",
			x"0000" when x"808D",
			x"0000" when x"808E",
			x"0000" when x"808F",
			x"0000" when x"8090",
			x"0000" when x"8091",
			x"0000" when x"8092",
			x"0000" when x"8093",
			x"0000" when x"8094",
			x"0000" when x"8095",
			x"0000" when x"8096",
			x"0000" when x"8097",
			x"0000" when x"8098",
			x"0000" when x"8099",
			x"0000" when x"809A",
			x"0000" when x"809B",
			x"0000" when x"809C",
			x"0000" when x"809D",
			x"0000" when x"809E",
			x"0000" when x"809F",
			x"0000" when x"80A0",
			x"0000" when x"80A1",
			x"0000" when x"80A2",
			x"0000" when x"80A3",
			x"0000" when x"80A4",
			x"0000" when x"80A5",
			x"0000" when x"80A6",
			x"0000" when x"80A7",
			x"0000" when x"80A8",
			x"0000" when x"80A9",
			x"0000" when x"80AA",
			x"0000" when x"80AB",
			x"0000" when x"80AC",
			x"0000" when x"80AD",
			x"0000" when x"80AE",
			x"0000" when x"80AF",
			x"0000" when x"80B0",
			x"0000" when x"80B1",
			x"0000" when x"80B2",
			x"0000" when x"80B3",
			x"0000" when x"80B4",
			x"0000" when x"80B5",
			x"0000" when x"80B6",
			x"0000" when x"80B7",
			x"0000" when x"80B8",
			x"0000" when x"80B9",
			x"0000" when x"80BA",
			x"0000" when x"80BB",
			x"0000" when x"80BC",
			x"0000" when x"80BD",
			x"0000" when x"80BE",
			x"0000" when x"80BF",
			x"0000" when x"80C0",
			x"0000" when x"80C1",
			x"0000" when x"80C2",
			x"0000" when x"80C3",
			x"0000" when x"80C4",
			x"0000" when x"80C5",
			x"0000" when x"80C6",
			x"0000" when x"80C7",
			x"0000" when x"80C8",
			x"0000" when x"80C9",
			x"0000" when x"80CA",
			x"0000" when x"80CB",
			x"0000" when x"80CC",
			x"0000" when x"80CD",
			x"0000" when x"80CE",
			x"0000" when x"80CF",
			x"0000" when x"80D0",
			x"0000" when x"80D1",
			x"0000" when x"80D2",
			x"0000" when x"80D3",
			x"0000" when x"80D4",
			x"0000" when x"80D5",
			x"0000" when x"80D6",
			x"0000" when x"80D7",
			x"0000" when x"80D8",
			x"0000" when x"80D9",
			x"0000" when x"80DA",
			x"0000" when x"80DB",
			x"0000" when x"80DC",
			x"0000" when x"80DD",
			x"0000" when x"80DE",
			x"0000" when x"80DF",
			x"0000" when x"80E0",
			x"0000" when x"80E1",
			x"0000" when x"80E2",
			x"0000" when x"80E3",
			x"0000" when x"80E4",
			x"0000" when x"80E5",
			x"0000" when x"80E6",
			x"0000" when x"80E7",
			x"0000" when x"80E8",
			x"0000" when x"80E9",
			x"0000" when x"80EA",
			x"0000" when x"80EB",
			x"0000" when x"80EC",
			x"0000" when x"80ED",
			x"0000" when x"80EE",
			x"0000" when x"80EF",
			x"0000" when x"80F0",
			x"0000" when x"80F1",
			x"0000" when x"80F2",
			x"0000" when x"80F3",
			x"0000" when x"80F4",
			x"0000" when x"80F5",
			x"0000" when x"80F6",
			x"0000" when x"80F7",
			x"0000" when x"80F8",
			x"0000" when x"80F9",
			x"0000" when x"80FA",
			x"0000" when x"80FB",
			x"0000" when x"80FC",
			x"0000" when x"80FD",
			x"0000" when x"80FE",
			x"0000" when x"80FF",
			x"0000" when x"8100",
			x"0000" when x"8101",
			x"0000" when x"8102",
			x"0000" when x"8103",
			x"0000" when x"8104",
			x"0000" when x"8105",
			x"0000" when x"8106",
			x"0000" when x"8107",
			x"0000" when x"8108",
			x"0000" when x"8109",
			x"0000" when x"810A",
			x"0000" when x"810B",
			x"0000" when x"810C",
			x"0000" when x"810D",
			x"0000" when x"810E",
			x"0000" when x"810F",
			x"0000" when x"8110",
			x"0000" when x"8111",
			x"0000" when x"8112",
			x"0000" when x"8113",
			x"0000" when x"8114",
			x"0000" when x"8115",
			x"0000" when x"8116",
			x"0000" when x"8117",
			x"0000" when x"8118",
			x"0000" when x"8119",
			x"0000" when x"811A",
			x"0000" when x"811B",
			x"0000" when x"811C",
			x"0000" when x"811D",
			x"0000" when x"811E",
			x"0000" when x"811F",
			x"0000" when x"8120",
			x"0000" when x"8121",
			x"0000" when x"8122",
			x"0000" when x"8123",
			x"0000" when x"8124",
			x"0000" when x"8125",
			x"0000" when x"8126",
			x"0000" when x"8127",
			x"0000" when x"8128",
			x"0000" when x"8129",
			x"0000" when x"812A",
			x"0000" when x"812B",
			x"0000" when x"812C",
			x"0000" when x"812D",
			x"0000" when x"812E",
			x"0000" when x"812F",
			x"0000" when x"8130",
			x"0000" when x"8131",
			x"0000" when x"8132",
			x"0000" when x"8133",
			x"0000" when x"8134",
			x"0000" when x"8135",
			x"0000" when x"8136",
			x"0000" when x"8137",
			x"0000" when x"8138",
			x"0000" when x"8139",
			x"0000" when x"813A",
			x"0000" when x"813B",
			x"0000" when x"813C",
			x"0000" when x"813D",
			x"0000" when x"813E",
			x"0000" when x"813F",
			x"0000" when x"8140",
			x"0000" when x"8141",
			x"0000" when x"8142",
			x"0000" when x"8143",
			x"0000" when x"8144",
			x"0000" when x"8145",
			x"0000" when x"8146",
			x"0000" when x"8147",
			x"0000" when x"8148",
			x"0000" when x"8149",
			x"0000" when x"814A",
			x"0000" when x"814B",
			x"0000" when x"814C",
			x"0000" when x"814D",
			x"0000" when x"814E",
			x"0000" when x"814F",
			x"0000" when x"8150",
			x"0000" when x"8151",
			x"0000" when x"8152",
			x"0000" when x"8153",
			x"0000" when x"8154",
			x"0000" when x"8155",
			x"0000" when x"8156",
			x"0000" when x"8157",
			x"0000" when x"8158",
			x"0000" when x"8159",
			x"0000" when x"815A",
			x"0000" when x"815B",
			x"0000" when x"815C",
			x"0000" when x"815D",
			x"0000" when x"815E",
			x"0000" when x"815F",
			x"0000" when x"8160",
			x"0000" when x"8161",
			x"0000" when x"8162",
			x"0000" when x"8163",
			x"0000" when x"8164",
			x"0000" when x"8165",
			x"0000" when x"8166",
			x"0000" when x"8167",
			x"0000" when x"8168",
			x"0000" when x"8169",
			x"0000" when x"816A",
			x"0000" when x"816B",
			x"0000" when x"816C",
			x"0000" when x"816D",
			x"0000" when x"816E",
			x"0000" when x"816F",
			x"0000" when x"8170",
			x"0000" when x"8171",
			x"0000" when x"8172",
			x"0000" when x"8173",
			x"0000" when x"8174",
			x"0000" when x"8175",
			x"0000" when x"8176",
			x"0000" when x"8177",
			x"0000" when x"8178",
			x"0000" when x"8179",
			x"0000" when x"817A",
			x"0000" when x"817B",
			x"0000" when x"817C",
			x"0000" when x"817D",
			x"0000" when x"817E",
			x"0000" when x"817F",
			x"0000" when x"8180",
			x"0000" when x"8181",
			x"0000" when x"8182",
			x"0000" when x"8183",
			x"0000" when x"8184",
			x"0000" when x"8185",
			x"0000" when x"8186",
			x"0000" when x"8187",
			x"0000" when x"8188",
			x"0000" when x"8189",
			x"0000" when x"818A",
			x"0000" when x"818B",
			x"0000" when x"818C",
			x"0000" when x"818D",
			x"0000" when x"818E",
			x"0000" when x"818F",
			x"0000" when x"8190",
			x"0000" when x"8191",
			x"0000" when x"8192",
			x"0000" when x"8193",
			x"0000" when x"8194",
			x"0000" when x"8195",
			x"0000" when x"8196",
			x"0000" when x"8197",
			x"0000" when x"8198",
			x"0000" when x"8199",
			x"0000" when x"819A",
			x"0000" when x"819B",
			x"0000" when x"819C",
			x"0000" when x"819D",
			x"0000" when x"819E",
			x"0000" when x"819F",
			x"0000" when x"81A0",
			x"0000" when x"81A1",
			x"0000" when x"81A2",
			x"0000" when x"81A3",
			x"0000" when x"81A4",
			x"0000" when x"81A5",
			x"0000" when x"81A6",
			x"0000" when x"81A7",
			x"0000" when x"81A8",
			x"0000" when x"81A9",
			x"0000" when x"81AA",
			x"0000" when x"81AB",
			x"0000" when x"81AC",
			x"0000" when x"81AD",
			x"0000" when x"81AE",
			x"0000" when x"81AF",
			x"0000" when x"81B0",
			x"0000" when x"81B1",
			x"0000" when x"81B2",
			x"0000" when x"81B3",
			x"0000" when x"81B4",
			x"0000" when x"81B5",
			x"0000" when x"81B6",
			x"0000" when x"81B7",
			x"0000" when x"81B8",
			x"0000" when x"81B9",
			x"0000" when x"81BA",
			x"0000" when x"81BB",
			x"0000" when x"81BC",
			x"0000" when x"81BD",
			x"0000" when x"81BE",
			x"0000" when x"81BF",
			x"0000" when x"81C0",
			x"0000" when x"81C1",
			x"0000" when x"81C2",
			x"0000" when x"81C3",
			x"0000" when x"81C4",
			x"0000" when x"81C5",
			x"0000" when x"81C6",
			x"0000" when x"81C7",
			x"0000" when x"81C8",
			x"0000" when x"81C9",
			x"0000" when x"81CA",
			x"0000" when x"81CB",
			x"0000" when x"81CC",
			x"0000" when x"81CD",
			x"0000" when x"81CE",
			x"0000" when x"81CF",
			x"0000" when x"81D0",
			x"0000" when x"81D1",
			x"0000" when x"81D2",
			x"0000" when x"81D3",
			x"0000" when x"81D4",
			x"0000" when x"81D5",
			x"0000" when x"81D6",
			x"0000" when x"81D7",
			x"0000" when x"81D8",
			x"0000" when x"81D9",
			x"0000" when x"81DA",
			x"0000" when x"81DB",
			x"0000" when x"81DC",
			x"0000" when x"81DD",
			x"0000" when x"81DE",
			x"0000" when x"81DF",
			x"0000" when x"81E0",
			x"0000" when x"81E1",
			x"0000" when x"81E2",
			x"0000" when x"81E3",
			x"0000" when x"81E4",
			x"0000" when x"81E5",
			x"0000" when x"81E6",
			x"0000" when x"81E7",
			x"0000" when x"81E8",
			x"0000" when x"81E9",
			x"0000" when x"81EA",
			x"0000" when x"81EB",
			x"0000" when x"81EC",
			x"0000" when x"81ED",
			x"0000" when x"81EE",
			x"0000" when x"81EF",
			x"0000" when x"81F0",
			x"0000" when x"81F1",
			x"0000" when x"81F2",
			x"0000" when x"81F3",
			x"0000" when x"81F4",
			x"0000" when x"81F5",
			x"0000" when x"81F6",
			x"0000" when x"81F7",
			x"0000" when x"81F8",
			x"0000" when x"81F9",
			x"0000" when x"81FA",
			x"0000" when x"81FB",
			x"0000" when x"81FC",
			x"0000" when x"81FD",
			x"0000" when x"81FE",
			x"0000" when x"81FF",
			x"0000" when x"8200",
			x"0000" when x"8201",
			x"0000" when x"8202",
			x"0000" when x"8203",
			x"0000" when x"8204",
			x"0000" when x"8205",
			x"0000" when x"8206",
			x"0000" when x"8207",
			x"0000" when x"8208",
			x"0000" when x"8209",
			x"0000" when x"820A",
			x"0000" when x"820B",
			x"0000" when x"820C",
			x"0000" when x"820D",
			x"0000" when x"820E",
			x"0000" when x"820F",
			x"0000" when x"8210",
			x"0000" when x"8211",
			x"0000" when x"8212",
			x"0000" when x"8213",
			x"0000" when x"8214",
			x"0000" when x"8215",
			x"0000" when x"8216",
			x"0000" when x"8217",
			x"0000" when x"8218",
			x"0000" when x"8219",
			x"0000" when x"821A",
			x"0000" when x"821B",
			x"0000" when x"821C",
			x"0000" when x"821D",
			x"0000" when x"821E",
			x"0000" when x"821F",
			x"0000" when x"8220",
			x"0000" when x"8221",
			x"0000" when x"8222",
			x"0000" when x"8223",
			x"0000" when x"8224",
			x"0000" when x"8225",
			x"0000" when x"8226",
			x"0000" when x"8227",
			x"0000" when x"8228",
			x"0000" when x"8229",
			x"0000" when x"822A",
			x"0000" when x"822B",
			x"0000" when x"822C",
			x"0000" when x"822D",
			x"0000" when x"822E",
			x"0000" when x"822F",
			x"0000" when x"8230",
			x"0000" when x"8231",
			x"0000" when x"8232",
			x"0000" when x"8233",
			x"0000" when x"8234",
			x"0000" when x"8235",
			x"0000" when x"8236",
			x"0000" when x"8237",
			x"0000" when x"8238",
			x"0000" when x"8239",
			x"0000" when x"823A",
			x"0000" when x"823B",
			x"0000" when x"823C",
			x"0000" when x"823D",
			x"0000" when x"823E",
			x"0000" when x"823F",
			x"0000" when x"8240",
			x"0000" when x"8241",
			x"0000" when x"8242",
			x"0000" when x"8243",
			x"0000" when x"8244",
			x"0000" when x"8245",
			x"0000" when x"8246",
			x"0000" when x"8247",
			x"0000" when x"8248",
			x"0000" when x"8249",
			x"0000" when x"824A",
			x"0000" when x"824B",
			x"0000" when x"824C",
			x"0000" when x"824D",
			x"0000" when x"824E",
			x"0000" when x"824F",
			x"0000" when x"8250",
			x"0000" when x"8251",
			x"0000" when x"8252",
			x"0000" when x"8253",
			x"0000" when x"8254",
			x"0000" when x"8255",
			x"0000" when x"8256",
			x"0000" when x"8257",
			x"0000" when x"8258",
			x"0000" when x"8259",
			x"0000" when x"825A",
			x"0000" when x"825B",
			x"0000" when x"825C",
			x"0000" when x"825D",
			x"0000" when x"825E",
			x"0000" when x"825F",
			x"0000" when x"8260",
			x"0000" when x"8261",
			x"0000" when x"8262",
			x"0000" when x"8263",
			x"0000" when x"8264",
			x"0000" when x"8265",
			x"0000" when x"8266",
			x"0000" when x"8267",
			x"0000" when x"8268",
			x"0000" when x"8269",
			x"0000" when x"826A",
			x"0000" when x"826B",
			x"0000" when x"826C",
			x"0000" when x"826D",
			x"0000" when x"826E",
			x"0000" when x"826F",
			x"0000" when x"8270",
			x"0000" when x"8271",
			x"0000" when x"8272",
			x"0000" when x"8273",
			x"0000" when x"8274",
			x"0000" when x"8275",
			x"0000" when x"8276",
			x"0000" when x"8277",
			x"0000" when x"8278",
			x"0000" when x"8279",
			x"0000" when x"827A",
			x"0000" when x"827B",
			x"0000" when x"827C",
			x"0000" when x"827D",
			x"0000" when x"827E",
			x"0000" when x"827F",
			x"0000" when x"8280",
			x"0000" when x"8281",
			x"0000" when x"8282",
			x"0000" when x"8283",
			x"0000" when x"8284",
			x"0000" when x"8285",
			x"0000" when x"8286",
			x"0000" when x"8287",
			x"0000" when x"8288",
			x"0000" when x"8289",
			x"0000" when x"828A",
			x"0000" when x"828B",
			x"0000" when x"828C",
			x"0000" when x"828D",
			x"0000" when x"828E",
			x"0000" when x"828F",
			x"0000" when x"8290",
			x"0000" when x"8291",
			x"0000" when x"8292",
			x"0000" when x"8293",
			x"0000" when x"8294",
			x"0000" when x"8295",
			x"0000" when x"8296",
			x"0000" when x"8297",
			x"0000" when x"8298",
			x"0000" when x"8299",
			x"0000" when x"829A",
			x"0000" when x"829B",
			x"0000" when x"829C",
			x"0000" when x"829D",
			x"0000" when x"829E",
			x"0000" when x"829F",
			x"0000" when x"82A0",
			x"0000" when x"82A1",
			x"0000" when x"82A2",
			x"0000" when x"82A3",
			x"0000" when x"82A4",
			x"0000" when x"82A5",
			x"0000" when x"82A6",
			x"0000" when x"82A7",
			x"0000" when x"82A8",
			x"0000" when x"82A9",
			x"0000" when x"82AA",
			x"0000" when x"82AB",
			x"0000" when x"82AC",
			x"0000" when x"82AD",
			x"0000" when x"82AE",
			x"0000" when x"82AF",
			x"0000" when x"82B0",
			x"0000" when x"82B1",
			x"0000" when x"82B2",
			x"0000" when x"82B3",
			x"0000" when x"82B4",
			x"0000" when x"82B5",
			x"0000" when x"82B6",
			x"0000" when x"82B7",
			x"0000" when x"82B8",
			x"0000" when x"82B9",
			x"0000" when x"82BA",
			x"0000" when x"82BB",
			x"0000" when x"82BC",
			x"0000" when x"82BD",
			x"0000" when x"82BE",
			x"0000" when x"82BF",
			x"0000" when x"82C0",
			x"0000" when x"82C1",
			x"0000" when x"82C2",
			x"0000" when x"82C3",
			x"0000" when x"82C4",
			x"0000" when x"82C5",
			x"0000" when x"82C6",
			x"0000" when x"82C7",
			x"0000" when x"82C8",
			x"0000" when x"82C9",
			x"0000" when x"82CA",
			x"0000" when x"82CB",
			x"0000" when x"82CC",
			x"0000" when x"82CD",
			x"0000" when x"82CE",
			x"0000" when x"82CF",
			x"0000" when x"82D0",
			x"0000" when x"82D1",
			x"0000" when x"82D2",
			x"0000" when x"82D3",
			x"0000" when x"82D4",
			x"0000" when x"82D5",
			x"0000" when x"82D6",
			x"0000" when x"82D7",
			x"0000" when x"82D8",
			x"0000" when x"82D9",
			x"0000" when x"82DA",
			x"0000" when x"82DB",
			x"0000" when x"82DC",
			x"0000" when x"82DD",
			x"0000" when x"82DE",
			x"0000" when x"82DF",
			x"0000" when x"82E0",
			x"0000" when x"82E1",
			x"0000" when x"82E2",
			x"0000" when x"82E3",
			x"0000" when x"82E4",
			x"0000" when x"82E5",
			x"0000" when x"82E6",
			x"0000" when x"82E7",
			x"0000" when x"82E8",
			x"0000" when x"82E9",
			x"0000" when x"82EA",
			x"0000" when x"82EB",
			x"0000" when x"82EC",
			x"0000" when x"82ED",
			x"0000" when x"82EE",
			x"0000" when x"82EF",
			x"0000" when x"82F0",
			x"0000" when x"82F1",
			x"0000" when x"82F2",
			x"0000" when x"82F3",
			x"0000" when x"82F4",
			x"0000" when x"82F5",
			x"0000" when x"82F6",
			x"0000" when x"82F7",
			x"0000" when x"82F8",
			x"0000" when x"82F9",
			x"0000" when x"82FA",
			x"0000" when x"82FB",
			x"0000" when x"82FC",
			x"0000" when x"82FD",
			x"0000" when x"82FE",
			x"0000" when x"82FF",
			x"0000" when x"8300",
			x"0000" when x"8301",
			x"0000" when x"8302",
			x"0000" when x"8303",
			x"0000" when x"8304",
			x"0000" when x"8305",
			x"0000" when x"8306",
			x"0000" when x"8307",
			x"0000" when x"8308",
			x"0000" when x"8309",
			x"0000" when x"830A",
			x"0000" when x"830B",
			x"0000" when x"830C",
			x"0000" when x"830D",
			x"0000" when x"830E",
			x"0000" when x"830F",
			x"0000" when x"8310",
			x"0000" when x"8311",
			x"0000" when x"8312",
			x"0000" when x"8313",
			x"0000" when x"8314",
			x"0000" when x"8315",
			x"0000" when x"8316",
			x"0000" when x"8317",
			x"0000" when x"8318",
			x"0000" when x"8319",
			x"0000" when x"831A",
			x"0000" when x"831B",
			x"0000" when x"831C",
			x"0000" when x"831D",
			x"0000" when x"831E",
			x"0000" when x"831F",
			x"0000" when x"8320",
			x"0000" when x"8321",
			x"0000" when x"8322",
			x"0000" when x"8323",
			x"0000" when x"8324",
			x"0000" when x"8325",
			x"0000" when x"8326",
			x"0000" when x"8327",
			x"0000" when x"8328",
			x"0000" when x"8329",
			x"0000" when x"832A",
			x"0000" when x"832B",
			x"0000" when x"832C",
			x"0000" when x"832D",
			x"0000" when x"832E",
			x"0000" when x"832F",
			x"0000" when x"8330",
			x"0000" when x"8331",
			x"0000" when x"8332",
			x"0000" when x"8333",
			x"0000" when x"8334",
			x"0000" when x"8335",
			x"0000" when x"8336",
			x"0000" when x"8337",
			x"0000" when x"8338",
			x"0000" when x"8339",
			x"0000" when x"833A",
			x"0000" when x"833B",
			x"0000" when x"833C",
			x"0000" when x"833D",
			x"0000" when x"833E",
			x"0000" when x"833F",
			x"0000" when x"8340",
			x"0000" when x"8341",
			x"0000" when x"8342",
			x"0000" when x"8343",
			x"0000" when x"8344",
			x"0000" when x"8345",
			x"0000" when x"8346",
			x"0000" when x"8347",
			x"0000" when x"8348",
			x"0000" when x"8349",
			x"0000" when x"834A",
			x"0000" when x"834B",
			x"0000" when x"834C",
			x"0000" when x"834D",
			x"0000" when x"834E",
			x"0000" when x"834F",
			x"0000" when x"8350",
			x"0000" when x"8351",
			x"0000" when x"8352",
			x"0000" when x"8353",
			x"0000" when x"8354",
			x"0000" when x"8355",
			x"0000" when x"8356",
			x"0000" when x"8357",
			x"0000" when x"8358",
			x"0000" when x"8359",
			x"0000" when x"835A",
			x"0000" when x"835B",
			x"0000" when x"835C",
			x"0000" when x"835D",
			x"0000" when x"835E",
			x"0000" when x"835F",
			x"0000" when x"8360",
			x"0000" when x"8361",
			x"0000" when x"8362",
			x"0000" when x"8363",
			x"0000" when x"8364",
			x"0000" when x"8365",
			x"0000" when x"8366",
			x"0000" when x"8367",
			x"0000" when x"8368",
			x"0000" when x"8369",
			x"0000" when x"836A",
			x"0000" when x"836B",
			x"0000" when x"836C",
			x"0000" when x"836D",
			x"0000" when x"836E",
			x"0000" when x"836F",
			x"0000" when x"8370",
			x"0000" when x"8371",
			x"0000" when x"8372",
			x"0000" when x"8373",
			x"0000" when x"8374",
			x"0000" when x"8375",
			x"0000" when x"8376",
			x"0000" when x"8377",
			x"0000" when x"8378",
			x"0000" when x"8379",
			x"0000" when x"837A",
			x"0000" when x"837B",
			x"0000" when x"837C",
			x"0000" when x"837D",
			x"0000" when x"837E",
			x"0000" when x"837F",
			x"0000" when x"8380",
			x"0000" when x"8381",
			x"0000" when x"8382",
			x"0000" when x"8383",
			x"0000" when x"8384",
			x"0000" when x"8385",
			x"0000" when x"8386",
			x"0000" when x"8387",
			x"0000" when x"8388",
			x"0000" when x"8389",
			x"0000" when x"838A",
			x"0000" when x"838B",
			x"0000" when x"838C",
			x"0000" when x"838D",
			x"0000" when x"838E",
			x"0000" when x"838F",
			x"0000" when x"8390",
			x"0000" when x"8391",
			x"0000" when x"8392",
			x"0000" when x"8393",
			x"0000" when x"8394",
			x"0000" when x"8395",
			x"0000" when x"8396",
			x"0000" when x"8397",
			x"0000" when x"8398",
			x"0000" when x"8399",
			x"0000" when x"839A",
			x"0000" when x"839B",
			x"0000" when x"839C",
			x"0000" when x"839D",
			x"0000" when x"839E",
			x"0000" when x"839F",
			x"0000" when x"83A0",
			x"0000" when x"83A1",
			x"0000" when x"83A2",
			x"0000" when x"83A3",
			x"0000" when x"83A4",
			x"0000" when x"83A5",
			x"0000" when x"83A6",
			x"0000" when x"83A7",
			x"0000" when x"83A8",
			x"0000" when x"83A9",
			x"0000" when x"83AA",
			x"0000" when x"83AB",
			x"0000" when x"83AC",
			x"0000" when x"83AD",
			x"0000" when x"83AE",
			x"0000" when x"83AF",
			x"0000" when x"83B0",
			x"0000" when x"83B1",
			x"0000" when x"83B2",
			x"0000" when x"83B3",
			x"0000" when x"83B4",
			x"0000" when x"83B5",
			x"0000" when x"83B6",
			x"0000" when x"83B7",
			x"0000" when x"83B8",
			x"0000" when x"83B9",
			x"0000" when x"83BA",
			x"0000" when x"83BB",
			x"0000" when x"83BC",
			x"0000" when x"83BD",
			x"0000" when x"83BE",
			x"0000" when x"83BF",
			x"0000" when x"83C0",
			x"0000" when x"83C1",
			x"0000" when x"83C2",
			x"0000" when x"83C3",
			x"0000" when x"83C4",
			x"0000" when x"83C5",
			x"0000" when x"83C6",
			x"0000" when x"83C7",
			x"0000" when x"83C8",
			x"0000" when x"83C9",
			x"0000" when x"83CA",
			x"0000" when x"83CB",
			x"0000" when x"83CC",
			x"0000" when x"83CD",
			x"0000" when x"83CE",
			x"0000" when x"83CF",
			x"0000" when x"83D0",
			x"0000" when x"83D1",
			x"0000" when x"83D2",
			x"0000" when x"83D3",
			x"0000" when x"83D4",
			x"0000" when x"83D5",
			x"0000" when x"83D6",
			x"0000" when x"83D7",
			x"0000" when x"83D8",
			x"0000" when x"83D9",
			x"0000" when x"83DA",
			x"0000" when x"83DB",
			x"0000" when x"83DC",
			x"0000" when x"83DD",
			x"0000" when x"83DE",
			x"0000" when x"83DF",
			x"0000" when x"83E0",
			x"0000" when x"83E1",
			x"0000" when x"83E2",
			x"0000" when x"83E3",
			x"0000" when x"83E4",
			x"0000" when x"83E5",
			x"0000" when x"83E6",
			x"0000" when x"83E7",
			x"0000" when x"83E8",
			x"0000" when x"83E9",
			x"0000" when x"83EA",
			x"0000" when x"83EB",
			x"0000" when x"83EC",
			x"0000" when x"83ED",
			x"0000" when x"83EE",
			x"0000" when x"83EF",
			x"0000" when x"83F0",
			x"0000" when x"83F1",
			x"0000" when x"83F2",
			x"0000" when x"83F3",
			x"0000" when x"83F4",
			x"0000" when x"83F5",
			x"0000" when x"83F6",
			x"0000" when x"83F7",
			x"0000" when x"83F8",
			x"0000" when x"83F9",
			x"0000" when x"83FA",
			x"0000" when x"83FB",
			x"0000" when x"83FC",
			x"0000" when x"83FD",
			x"0000" when x"83FE",
			x"0000" when x"83FF",
			x"0000" when x"8400",
			x"0000" when x"8401",
			x"0000" when x"8402",
			x"0000" when x"8403",
			x"0000" when x"8404",
			x"0000" when x"8405",
			x"0000" when x"8406",
			x"0000" when x"8407",
			x"0000" when x"8408",
			x"0000" when x"8409",
			x"0000" when x"840A",
			x"0000" when x"840B",
			x"0000" when x"840C",
			x"0000" when x"840D",
			x"0000" when x"840E",
			x"0000" when x"840F",
			x"0000" when x"8410",
			x"0000" when x"8411",
			x"0000" when x"8412",
			x"0000" when x"8413",
			x"0000" when x"8414",
			x"0000" when x"8415",
			x"0000" when x"8416",
			x"0000" when x"8417",
			x"0000" when x"8418",
			x"0000" when x"8419",
			x"0000" when x"841A",
			x"0000" when x"841B",
			x"0000" when x"841C",
			x"0000" when x"841D",
			x"0000" when x"841E",
			x"0000" when x"841F",
			x"0000" when x"8420",
			x"0000" when x"8421",
			x"0000" when x"8422",
			x"0000" when x"8423",
			x"0000" when x"8424",
			x"0000" when x"8425",
			x"0000" when x"8426",
			x"0000" when x"8427",
			x"0000" when x"8428",
			x"0000" when x"8429",
			x"0000" when x"842A",
			x"0000" when x"842B",
			x"0000" when x"842C",
			x"0000" when x"842D",
			x"0000" when x"842E",
			x"0000" when x"842F",
			x"0000" when x"8430",
			x"0000" when x"8431",
			x"0000" when x"8432",
			x"0000" when x"8433",
			x"0000" when x"8434",
			x"0000" when x"8435",
			x"0000" when x"8436",
			x"0000" when x"8437",
			x"0000" when x"8438",
			x"0000" when x"8439",
			x"0000" when x"843A",
			x"0000" when x"843B",
			x"0000" when x"843C",
			x"0000" when x"843D",
			x"0000" when x"843E",
			x"0000" when x"843F",
			x"0000" when x"8440",
			x"0000" when x"8441",
			x"0000" when x"8442",
			x"0000" when x"8443",
			x"0000" when x"8444",
			x"0000" when x"8445",
			x"0000" when x"8446",
			x"0000" when x"8447",
			x"0000" when x"8448",
			x"0000" when x"8449",
			x"0000" when x"844A",
			x"0000" when x"844B",
			x"0000" when x"844C",
			x"0000" when x"844D",
			x"0000" when x"844E",
			x"0000" when x"844F",
			x"0000" when x"8450",
			x"0000" when x"8451",
			x"0000" when x"8452",
			x"0000" when x"8453",
			x"0000" when x"8454",
			x"0000" when x"8455",
			x"0000" when x"8456",
			x"0000" when x"8457",
			x"0000" when x"8458",
			x"0000" when x"8459",
			x"0000" when x"845A",
			x"0000" when x"845B",
			x"0000" when x"845C",
			x"0000" when x"845D",
			x"0000" when x"845E",
			x"0000" when x"845F",
			x"0000" when x"8460",
			x"0000" when x"8461",
			x"0000" when x"8462",
			x"0000" when x"8463",
			x"0000" when x"8464",
			x"0000" when x"8465",
			x"0000" when x"8466",
			x"0000" when x"8467",
			x"0000" when x"8468",
			x"0000" when x"8469",
			x"0000" when x"846A",
			x"0000" when x"846B",
			x"0000" when x"846C",
			x"0000" when x"846D",
			x"0000" when x"846E",
			x"0000" when x"846F",
			x"0000" when x"8470",
			x"0000" when x"8471",
			x"0000" when x"8472",
			x"0000" when x"8473",
			x"0000" when x"8474",
			x"0000" when x"8475",
			x"0000" when x"8476",
			x"0000" when x"8477",
			x"0000" when x"8478",
			x"0000" when x"8479",
			x"0000" when x"847A",
			x"0000" when x"847B",
			x"0000" when x"847C",
			x"0000" when x"847D",
			x"0000" when x"847E",
			x"0000" when x"847F",
			x"0000" when x"8480",
			x"0000" when x"8481",
			x"0000" when x"8482",
			x"0000" when x"8483",
			x"0000" when x"8484",
			x"0000" when x"8485",
			x"0000" when x"8486",
			x"0000" when x"8487",
			x"0000" when x"8488",
			x"0000" when x"8489",
			x"0000" when x"848A",
			x"0000" when x"848B",
			x"0000" when x"848C",
			x"0000" when x"848D",
			x"0000" when x"848E",
			x"0000" when x"848F",
			x"0000" when x"8490",
			x"0000" when x"8491",
			x"0000" when x"8492",
			x"0000" when x"8493",
			x"0000" when x"8494",
			x"0000" when x"8495",
			x"0000" when x"8496",
			x"0000" when x"8497",
			x"0000" when x"8498",
			x"0000" when x"8499",
			x"0000" when x"849A",
			x"0000" when x"849B",
			x"0000" when x"849C",
			x"0000" when x"849D",
			x"0000" when x"849E",
			x"0000" when x"849F",
			x"0000" when x"84A0",
			x"0000" when x"84A1",
			x"0000" when x"84A2",
			x"0000" when x"84A3",
			x"0000" when x"84A4",
			x"0000" when x"84A5",
			x"0000" when x"84A6",
			x"0000" when x"84A7",
			x"0000" when x"84A8",
			x"0000" when x"84A9",
			x"0000" when x"84AA",
			x"0000" when x"84AB",
			x"0000" when x"84AC",
			x"0000" when x"84AD",
			x"0000" when x"84AE",
			x"0000" when x"84AF",
			x"0000" when x"84B0",
			x"0000" when x"84B1",
			x"0000" when x"84B2",
			x"0000" when x"84B3",
			x"0000" when x"84B4",
			x"0000" when x"84B5",
			x"0000" when x"84B6",
			x"0000" when x"84B7",
			x"0000" when x"84B8",
			x"0000" when x"84B9",
			x"0000" when x"84BA",
			x"0000" when x"84BB",
			x"0000" when x"84BC",
			x"0000" when x"84BD",
			x"0000" when x"84BE",
			x"0000" when x"84BF",
			x"0000" when x"84C0",
			x"0000" when x"84C1",
			x"0000" when x"84C2",
			x"0000" when x"84C3",
			x"0000" when x"84C4",
			x"0000" when x"84C5",
			x"0000" when x"84C6",
			x"0000" when x"84C7",
			x"0000" when x"84C8",
			x"0000" when x"84C9",
			x"0000" when x"84CA",
			x"0000" when x"84CB",
			x"0000" when x"84CC",
			x"0000" when x"84CD",
			x"0000" when x"84CE",
			x"0000" when x"84CF",
			x"0000" when x"84D0",
			x"0000" when x"84D1",
			x"0000" when x"84D2",
			x"0000" when x"84D3",
			x"0000" when x"84D4",
			x"0000" when x"84D5",
			x"0000" when x"84D6",
			x"0000" when x"84D7",
			x"0000" when x"84D8",
			x"0000" when x"84D9",
			x"0000" when x"84DA",
			x"0000" when x"84DB",
			x"0000" when x"84DC",
			x"0000" when x"84DD",
			x"0000" when x"84DE",
			x"0000" when x"84DF",
			x"0000" when x"84E0",
			x"0000" when x"84E1",
			x"0000" when x"84E2",
			x"0000" when x"84E3",
			x"0000" when x"84E4",
			x"0000" when x"84E5",
			x"0000" when x"84E6",
			x"0000" when x"84E7",
			x"0000" when x"84E8",
			x"0000" when x"84E9",
			x"0000" when x"84EA",
			x"0000" when x"84EB",
			x"0000" when x"84EC",
			x"0000" when x"84ED",
			x"0000" when x"84EE",
			x"0000" when x"84EF",
			x"0000" when x"84F0",
			x"0000" when x"84F1",
			x"0000" when x"84F2",
			x"0000" when x"84F3",
			x"0000" when x"84F4",
			x"0000" when x"84F5",
			x"0000" when x"84F6",
			x"0000" when x"84F7",
			x"0000" when x"84F8",
			x"0000" when x"84F9",
			x"0000" when x"84FA",
			x"0000" when x"84FB",
			x"0000" when x"84FC",
			x"0000" when x"84FD",
			x"0000" when x"84FE",
			x"0000" when x"84FF",
			x"0000" when x"8500",
			x"0000" when x"8501",
			x"0000" when x"8502",
			x"0000" when x"8503",
			x"0000" when x"8504",
			x"0000" when x"8505",
			x"0000" when x"8506",
			x"0000" when x"8507",
			x"0000" when x"8508",
			x"0000" when x"8509",
			x"0000" when x"850A",
			x"0000" when x"850B",
			x"0000" when x"850C",
			x"0000" when x"850D",
			x"0000" when x"850E",
			x"0000" when x"850F",
			x"0000" when x"8510",
			x"0000" when x"8511",
			x"0000" when x"8512",
			x"0000" when x"8513",
			x"0000" when x"8514",
			x"0000" when x"8515",
			x"0000" when x"8516",
			x"0000" when x"8517",
			x"0000" when x"8518",
			x"0000" when x"8519",
			x"0000" when x"851A",
			x"0000" when x"851B",
			x"0000" when x"851C",
			x"0000" when x"851D",
			x"0000" when x"851E",
			x"0000" when x"851F",
			x"0000" when x"8520",
			x"0000" when x"8521",
			x"0000" when x"8522",
			x"0000" when x"8523",
			x"0000" when x"8524",
			x"0000" when x"8525",
			x"0000" when x"8526",
			x"0000" when x"8527",
			x"0000" when x"8528",
			x"0000" when x"8529",
			x"0000" when x"852A",
			x"0000" when x"852B",
			x"0000" when x"852C",
			x"0000" when x"852D",
			x"0000" when x"852E",
			x"0000" when x"852F",
			x"0000" when x"8530",
			x"0000" when x"8531",
			x"0000" when x"8532",
			x"0000" when x"8533",
			x"0000" when x"8534",
			x"0000" when x"8535",
			x"0000" when x"8536",
			x"0000" when x"8537",
			x"0000" when x"8538",
			x"0000" when x"8539",
			x"0000" when x"853A",
			x"0000" when x"853B",
			x"0000" when x"853C",
			x"0000" when x"853D",
			x"0000" when x"853E",
			x"0000" when x"853F",
			x"0000" when x"8540",
			x"0000" when x"8541",
			x"0000" when x"8542",
			x"0000" when x"8543",
			x"0000" when x"8544",
			x"0000" when x"8545",
			x"0000" when x"8546",
			x"0000" when x"8547",
			x"0000" when x"8548",
			x"0000" when x"8549",
			x"0000" when x"854A",
			x"0000" when x"854B",
			x"0000" when x"854C",
			x"0000" when x"854D",
			x"0000" when x"854E",
			x"0000" when x"854F",
			x"0000" when x"8550",
			x"0000" when x"8551",
			x"0000" when x"8552",
			x"0000" when x"8553",
			x"0000" when x"8554",
			x"0000" when x"8555",
			x"0000" when x"8556",
			x"0000" when x"8557",
			x"0000" when x"8558",
			x"0000" when x"8559",
			x"0000" when x"855A",
			x"0000" when x"855B",
			x"0000" when x"855C",
			x"0000" when x"855D",
			x"0000" when x"855E",
			x"0000" when x"855F",
			x"0000" when x"8560",
			x"0000" when x"8561",
			x"0000" when x"8562",
			x"0000" when x"8563",
			x"0000" when x"8564",
			x"0000" when x"8565",
			x"0000" when x"8566",
			x"0000" when x"8567",
			x"0000" when x"8568",
			x"0000" when x"8569",
			x"0000" when x"856A",
			x"0000" when x"856B",
			x"0000" when x"856C",
			x"0000" when x"856D",
			x"0000" when x"856E",
			x"0000" when x"856F",
			x"0000" when x"8570",
			x"0000" when x"8571",
			x"0000" when x"8572",
			x"0000" when x"8573",
			x"0000" when x"8574",
			x"0000" when x"8575",
			x"0000" when x"8576",
			x"0000" when x"8577",
			x"0000" when x"8578",
			x"0000" when x"8579",
			x"0000" when x"857A",
			x"0000" when x"857B",
			x"0000" when x"857C",
			x"0000" when x"857D",
			x"0000" when x"857E",
			x"0000" when x"857F",
			x"0000" when x"8580",
			x"0000" when x"8581",
			x"0000" when x"8582",
			x"0000" when x"8583",
			x"0000" when x"8584",
			x"0000" when x"8585",
			x"0000" when x"8586",
			x"0000" when x"8587",
			x"0000" when x"8588",
			x"0000" when x"8589",
			x"0000" when x"858A",
			x"0000" when x"858B",
			x"0000" when x"858C",
			x"0000" when x"858D",
			x"0000" when x"858E",
			x"0000" when x"858F",
			x"0000" when x"8590",
			x"0000" when x"8591",
			x"0000" when x"8592",
			x"0000" when x"8593",
			x"0000" when x"8594",
			x"0000" when x"8595",
			x"0000" when x"8596",
			x"0000" when x"8597",
			x"0000" when x"8598",
			x"0000" when x"8599",
			x"0000" when x"859A",
			x"0000" when x"859B",
			x"0000" when x"859C",
			x"0000" when x"859D",
			x"0000" when x"859E",
			x"0000" when x"859F",
			x"0000" when x"85A0",
			x"0000" when x"85A1",
			x"0000" when x"85A2",
			x"0000" when x"85A3",
			x"0000" when x"85A4",
			x"0000" when x"85A5",
			x"0000" when x"85A6",
			x"0000" when x"85A7",
			x"0000" when x"85A8",
			x"0000" when x"85A9",
			x"0000" when x"85AA",
			x"0000" when x"85AB",
			x"0000" when x"85AC",
			x"0000" when x"85AD",
			x"0000" when x"85AE",
			x"0000" when x"85AF",
			x"0000" when x"85B0",
			x"0000" when x"85B1",
			x"0000" when x"85B2",
			x"0000" when x"85B3",
			x"0000" when x"85B4",
			x"0000" when x"85B5",
			x"0000" when x"85B6",
			x"0000" when x"85B7",
			x"0000" when x"85B8",
			x"0000" when x"85B9",
			x"0000" when x"85BA",
			x"0000" when x"85BB",
			x"0000" when x"85BC",
			x"0000" when x"85BD",
			x"0000" when x"85BE",
			x"0000" when x"85BF",
			x"0000" when x"85C0",
			x"0000" when x"85C1",
			x"0000" when x"85C2",
			x"0000" when x"85C3",
			x"0000" when x"85C4",
			x"0000" when x"85C5",
			x"0000" when x"85C6",
			x"0000" when x"85C7",
			x"0000" when x"85C8",
			x"0000" when x"85C9",
			x"0000" when x"85CA",
			x"0000" when x"85CB",
			x"0000" when x"85CC",
			x"0000" when x"85CD",
			x"0000" when x"85CE",
			x"0000" when x"85CF",
			x"0000" when x"85D0",
			x"0000" when x"85D1",
			x"0000" when x"85D2",
			x"0000" when x"85D3",
			x"0000" when x"85D4",
			x"0000" when x"85D5",
			x"0000" when x"85D6",
			x"0000" when x"85D7",
			x"0000" when x"85D8",
			x"0000" when x"85D9",
			x"0000" when x"85DA",
			x"0000" when x"85DB",
			x"0000" when x"85DC",
			x"0000" when x"85DD",
			x"0000" when x"85DE",
			x"0000" when x"85DF",
			x"0000" when x"85E0",
			x"0000" when x"85E1",
			x"0000" when x"85E2",
			x"0000" when x"85E3",
			x"0000" when x"85E4",
			x"0000" when x"85E5",
			x"0000" when x"85E6",
			x"0000" when x"85E7",
			x"0000" when x"85E8",
			x"0000" when x"85E9",
			x"0000" when x"85EA",
			x"0000" when x"85EB",
			x"0000" when x"85EC",
			x"0000" when x"85ED",
			x"0000" when x"85EE",
			x"0000" when x"85EF",
			x"0000" when x"85F0",
			x"0000" when x"85F1",
			x"0000" when x"85F2",
			x"0000" when x"85F3",
			x"0000" when x"85F4",
			x"0000" when x"85F5",
			x"0000" when x"85F6",
			x"0000" when x"85F7",
			x"0000" when x"85F8",
			x"0000" when x"85F9",
			x"0000" when x"85FA",
			x"0000" when x"85FB",
			x"0000" when x"85FC",
			x"0000" when x"85FD",
			x"0000" when x"85FE",
			x"0000" when x"85FF",
			x"0000" when x"8600",
			x"0000" when x"8601",
			x"0000" when x"8602",
			x"0000" when x"8603",
			x"0000" when x"8604",
			x"0000" when x"8605",
			x"0000" when x"8606",
			x"0000" when x"8607",
			x"0000" when x"8608",
			x"0000" when x"8609",
			x"0000" when x"860A",
			x"0000" when x"860B",
			x"0000" when x"860C",
			x"0000" when x"860D",
			x"0000" when x"860E",
			x"0000" when x"860F",
			x"0000" when x"8610",
			x"0000" when x"8611",
			x"0000" when x"8612",
			x"0000" when x"8613",
			x"0000" when x"8614",
			x"0000" when x"8615",
			x"0000" when x"8616",
			x"0000" when x"8617",
			x"0000" when x"8618",
			x"0000" when x"8619",
			x"0000" when x"861A",
			x"0000" when x"861B",
			x"0000" when x"861C",
			x"0000" when x"861D",
			x"0000" when x"861E",
			x"0000" when x"861F",
			x"0000" when x"8620",
			x"0000" when x"8621",
			x"0000" when x"8622",
			x"0000" when x"8623",
			x"0000" when x"8624",
			x"0000" when x"8625",
			x"0000" when x"8626",
			x"0000" when x"8627",
			x"0000" when x"8628",
			x"0000" when x"8629",
			x"0000" when x"862A",
			x"0000" when x"862B",
			x"0000" when x"862C",
			x"0000" when x"862D",
			x"0000" when x"862E",
			x"0000" when x"862F",
			x"0000" when x"8630",
			x"0000" when x"8631",
			x"0000" when x"8632",
			x"0000" when x"8633",
			x"0000" when x"8634",
			x"0000" when x"8635",
			x"0000" when x"8636",
			x"0000" when x"8637",
			x"0000" when x"8638",
			x"0000" when x"8639",
			x"0000" when x"863A",
			x"0000" when x"863B",
			x"0000" when x"863C",
			x"0000" when x"863D",
			x"0000" when x"863E",
			x"0000" when x"863F",
			x"0000" when x"8640",
			x"0000" when x"8641",
			x"0000" when x"8642",
			x"0000" when x"8643",
			x"0000" when x"8644",
			x"0000" when x"8645",
			x"0000" when x"8646",
			x"0000" when x"8647",
			x"0000" when x"8648",
			x"0000" when x"8649",
			x"0000" when x"864A",
			x"0000" when x"864B",
			x"0000" when x"864C",
			x"0000" when x"864D",
			x"0000" when x"864E",
			x"0000" when x"864F",
			x"0000" when x"8650",
			x"0000" when x"8651",
			x"0000" when x"8652",
			x"0000" when x"8653",
			x"0000" when x"8654",
			x"0000" when x"8655",
			x"0000" when x"8656",
			x"0000" when x"8657",
			x"0000" when x"8658",
			x"0000" when x"8659",
			x"0000" when x"865A",
			x"0000" when x"865B",
			x"0000" when x"865C",
			x"0000" when x"865D",
			x"0000" when x"865E",
			x"0000" when x"865F",
			x"0000" when x"8660",
			x"0000" when x"8661",
			x"0000" when x"8662",
			x"0000" when x"8663",
			x"0000" when x"8664",
			x"0000" when x"8665",
			x"0000" when x"8666",
			x"0000" when x"8667",
			x"0000" when x"8668",
			x"0000" when x"8669",
			x"0000" when x"866A",
			x"0000" when x"866B",
			x"0000" when x"866C",
			x"0000" when x"866D",
			x"0000" when x"866E",
			x"0000" when x"866F",
			x"0000" when x"8670",
			x"0000" when x"8671",
			x"0000" when x"8672",
			x"0000" when x"8673",
			x"0000" when x"8674",
			x"0000" when x"8675",
			x"0000" when x"8676",
			x"0000" when x"8677",
			x"0000" when x"8678",
			x"0000" when x"8679",
			x"0000" when x"867A",
			x"0000" when x"867B",
			x"0000" when x"867C",
			x"0000" when x"867D",
			x"0000" when x"867E",
			x"0000" when x"867F",
			x"0000" when x"8680",
			x"0000" when x"8681",
			x"0000" when x"8682",
			x"0000" when x"8683",
			x"0000" when x"8684",
			x"0000" when x"8685",
			x"0000" when x"8686",
			x"0000" when x"8687",
			x"0000" when x"8688",
			x"0000" when x"8689",
			x"0000" when x"868A",
			x"0000" when x"868B",
			x"0000" when x"868C",
			x"0000" when x"868D",
			x"0000" when x"868E",
			x"0000" when x"868F",
			x"0000" when x"8690",
			x"0000" when x"8691",
			x"0000" when x"8692",
			x"0000" when x"8693",
			x"0000" when x"8694",
			x"0000" when x"8695",
			x"0000" when x"8696",
			x"0000" when x"8697",
			x"0000" when x"8698",
			x"0000" when x"8699",
			x"0000" when x"869A",
			x"0000" when x"869B",
			x"0000" when x"869C",
			x"0000" when x"869D",
			x"0000" when x"869E",
			x"0000" when x"869F",
			x"0000" when x"86A0",
			x"0000" when x"86A1",
			x"0000" when x"86A2",
			x"0000" when x"86A3",
			x"0000" when x"86A4",
			x"0000" when x"86A5",
			x"0000" when x"86A6",
			x"0000" when x"86A7",
			x"0000" when x"86A8",
			x"0000" when x"86A9",
			x"0000" when x"86AA",
			x"0000" when x"86AB",
			x"0000" when x"86AC",
			x"0000" when x"86AD",
			x"0000" when x"86AE",
			x"0000" when x"86AF",
			x"0000" when x"86B0",
			x"0000" when x"86B1",
			x"0000" when x"86B2",
			x"0000" when x"86B3",
			x"0000" when x"86B4",
			x"0000" when x"86B5",
			x"0000" when x"86B6",
			x"0000" when x"86B7",
			x"0000" when x"86B8",
			x"0000" when x"86B9",
			x"0000" when x"86BA",
			x"0000" when x"86BB",
			x"0000" when x"86BC",
			x"0000" when x"86BD",
			x"0000" when x"86BE",
			x"0000" when x"86BF",
			x"0000" when x"86C0",
			x"0000" when x"86C1",
			x"0000" when x"86C2",
			x"0000" when x"86C3",
			x"0000" when x"86C4",
			x"0000" when x"86C5",
			x"0000" when x"86C6",
			x"0000" when x"86C7",
			x"0000" when x"86C8",
			x"0000" when x"86C9",
			x"0000" when x"86CA",
			x"0000" when x"86CB",
			x"0000" when x"86CC",
			x"0000" when x"86CD",
			x"0000" when x"86CE",
			x"0000" when x"86CF",
			x"0000" when x"86D0",
			x"0000" when x"86D1",
			x"0000" when x"86D2",
			x"0000" when x"86D3",
			x"0000" when x"86D4",
			x"0000" when x"86D5",
			x"0000" when x"86D6",
			x"0000" when x"86D7",
			x"0000" when x"86D8",
			x"0000" when x"86D9",
			x"0000" when x"86DA",
			x"0000" when x"86DB",
			x"0000" when x"86DC",
			x"0000" when x"86DD",
			x"0000" when x"86DE",
			x"0000" when x"86DF",
			x"0000" when x"86E0",
			x"0000" when x"86E1",
			x"0000" when x"86E2",
			x"0000" when x"86E3",
			x"0000" when x"86E4",
			x"0000" when x"86E5",
			x"0000" when x"86E6",
			x"0000" when x"86E7",
			x"0000" when x"86E8",
			x"0000" when x"86E9",
			x"0000" when x"86EA",
			x"0000" when x"86EB",
			x"0000" when x"86EC",
			x"0000" when x"86ED",
			x"0000" when x"86EE",
			x"0000" when x"86EF",
			x"0000" when x"86F0",
			x"0000" when x"86F1",
			x"0000" when x"86F2",
			x"0000" when x"86F3",
			x"0000" when x"86F4",
			x"0000" when x"86F5",
			x"0000" when x"86F6",
			x"0000" when x"86F7",
			x"0000" when x"86F8",
			x"0000" when x"86F9",
			x"0000" when x"86FA",
			x"0000" when x"86FB",
			x"0000" when x"86FC",
			x"0000" when x"86FD",
			x"0000" when x"86FE",
			x"0000" when x"86FF",
			x"0000" when x"8700",
			x"0000" when x"8701",
			x"0000" when x"8702",
			x"0000" when x"8703",
			x"0000" when x"8704",
			x"0000" when x"8705",
			x"0000" when x"8706",
			x"0000" when x"8707",
			x"0000" when x"8708",
			x"0000" when x"8709",
			x"0000" when x"870A",
			x"0000" when x"870B",
			x"0000" when x"870C",
			x"0000" when x"870D",
			x"0000" when x"870E",
			x"0000" when x"870F",
			x"0000" when x"8710",
			x"0000" when x"8711",
			x"0000" when x"8712",
			x"0000" when x"8713",
			x"0000" when x"8714",
			x"0000" when x"8715",
			x"0000" when x"8716",
			x"0000" when x"8717",
			x"0000" when x"8718",
			x"0000" when x"8719",
			x"0000" when x"871A",
			x"0000" when x"871B",
			x"0000" when x"871C",
			x"0000" when x"871D",
			x"0000" when x"871E",
			x"0000" when x"871F",
			x"0000" when x"8720",
			x"0000" when x"8721",
			x"0000" when x"8722",
			x"0000" when x"8723",
			x"0000" when x"8724",
			x"0000" when x"8725",
			x"0000" when x"8726",
			x"0000" when x"8727",
			x"0000" when x"8728",
			x"0000" when x"8729",
			x"0000" when x"872A",
			x"0000" when x"872B",
			x"0000" when x"872C",
			x"0000" when x"872D",
			x"0000" when x"872E",
			x"0000" when x"872F",
			x"0000" when x"8730",
			x"0000" when x"8731",
			x"0000" when x"8732",
			x"0000" when x"8733",
			x"0000" when x"8734",
			x"0000" when x"8735",
			x"0000" when x"8736",
			x"0000" when x"8737",
			x"0000" when x"8738",
			x"0000" when x"8739",
			x"0000" when x"873A",
			x"0000" when x"873B",
			x"0000" when x"873C",
			x"0000" when x"873D",
			x"0000" when x"873E",
			x"0000" when x"873F",
			x"0000" when x"8740",
			x"0000" when x"8741",
			x"0000" when x"8742",
			x"0000" when x"8743",
			x"0000" when x"8744",
			x"0000" when x"8745",
			x"0000" when x"8746",
			x"0000" when x"8747",
			x"0000" when x"8748",
			x"0000" when x"8749",
			x"0000" when x"874A",
			x"0000" when x"874B",
			x"0000" when x"874C",
			x"0000" when x"874D",
			x"0000" when x"874E",
			x"0000" when x"874F",
			x"0000" when x"8750",
			x"0000" when x"8751",
			x"0000" when x"8752",
			x"0000" when x"8753",
			x"0000" when x"8754",
			x"0000" when x"8755",
			x"0000" when x"8756",
			x"0000" when x"8757",
			x"0000" when x"8758",
			x"0000" when x"8759",
			x"0000" when x"875A",
			x"0000" when x"875B",
			x"0000" when x"875C",
			x"0000" when x"875D",
			x"0000" when x"875E",
			x"0000" when x"875F",
			x"0000" when x"8760",
			x"0000" when x"8761",
			x"0000" when x"8762",
			x"0000" when x"8763",
			x"0000" when x"8764",
			x"0000" when x"8765",
			x"0000" when x"8766",
			x"0000" when x"8767",
			x"0000" when x"8768",
			x"0000" when x"8769",
			x"0000" when x"876A",
			x"0000" when x"876B",
			x"0000" when x"876C",
			x"0000" when x"876D",
			x"0000" when x"876E",
			x"0000" when x"876F",
			x"0000" when x"8770",
			x"0000" when x"8771",
			x"0000" when x"8772",
			x"0000" when x"8773",
			x"0000" when x"8774",
			x"0000" when x"8775",
			x"0000" when x"8776",
			x"0000" when x"8777",
			x"0000" when x"8778",
			x"0000" when x"8779",
			x"0000" when x"877A",
			x"0000" when x"877B",
			x"0000" when x"877C",
			x"0000" when x"877D",
			x"0000" when x"877E",
			x"0000" when x"877F",
			x"0000" when x"8780",
			x"0000" when x"8781",
			x"0000" when x"8782",
			x"0000" when x"8783",
			x"0000" when x"8784",
			x"0000" when x"8785",
			x"0000" when x"8786",
			x"0000" when x"8787",
			x"0000" when x"8788",
			x"0000" when x"8789",
			x"0000" when x"878A",
			x"0000" when x"878B",
			x"0000" when x"878C",
			x"0000" when x"878D",
			x"0000" when x"878E",
			x"0000" when x"878F",
			x"0000" when x"8790",
			x"0000" when x"8791",
			x"0000" when x"8792",
			x"0000" when x"8793",
			x"0000" when x"8794",
			x"0000" when x"8795",
			x"0000" when x"8796",
			x"0000" when x"8797",
			x"0000" when x"8798",
			x"0000" when x"8799",
			x"0000" when x"879A",
			x"0000" when x"879B",
			x"0000" when x"879C",
			x"0000" when x"879D",
			x"0000" when x"879E",
			x"0000" when x"879F",
			x"0000" when x"87A0",
			x"0000" when x"87A1",
			x"0000" when x"87A2",
			x"0000" when x"87A3",
			x"0000" when x"87A4",
			x"0000" when x"87A5",
			x"0000" when x"87A6",
			x"0000" when x"87A7",
			x"0000" when x"87A8",
			x"0000" when x"87A9",
			x"0000" when x"87AA",
			x"0000" when x"87AB",
			x"0000" when x"87AC",
			x"0000" when x"87AD",
			x"0000" when x"87AE",
			x"0000" when x"87AF",
			x"0000" when x"87B0",
			x"0000" when x"87B1",
			x"0000" when x"87B2",
			x"0000" when x"87B3",
			x"0000" when x"87B4",
			x"0000" when x"87B5",
			x"0000" when x"87B6",
			x"0000" when x"87B7",
			x"0000" when x"87B8",
			x"0000" when x"87B9",
			x"0000" when x"87BA",
			x"0000" when x"87BB",
			x"0000" when x"87BC",
			x"0000" when x"87BD",
			x"0000" when x"87BE",
			x"0000" when x"87BF",
			x"0000" when x"87C0",
			x"0000" when x"87C1",
			x"0000" when x"87C2",
			x"0000" when x"87C3",
			x"0000" when x"87C4",
			x"0000" when x"87C5",
			x"0000" when x"87C6",
			x"0000" when x"87C7",
			x"0000" when x"87C8",
			x"0000" when x"87C9",
			x"0000" when x"87CA",
			x"0000" when x"87CB",
			x"0000" when x"87CC",
			x"0000" when x"87CD",
			x"0000" when x"87CE",
			x"0000" when x"87CF",
			x"0000" when x"87D0",
			x"0000" when x"87D1",
			x"0000" when x"87D2",
			x"0000" when x"87D3",
			x"0000" when x"87D4",
			x"0000" when x"87D5",
			x"0000" when x"87D6",
			x"0000" when x"87D7",
			x"0000" when x"87D8",
			x"0000" when x"87D9",
			x"0000" when x"87DA",
			x"0000" when x"87DB",
			x"0000" when x"87DC",
			x"0000" when x"87DD",
			x"0000" when x"87DE",
			x"0000" when x"87DF",
			x"0000" when x"87E0",
			x"0000" when x"87E1",
			x"0000" when x"87E2",
			x"0000" when x"87E3",
			x"0000" when x"87E4",
			x"0000" when x"87E5",
			x"0000" when x"87E6",
			x"0000" when x"87E7",
			x"0000" when x"87E8",
			x"0000" when x"87E9",
			x"0000" when x"87EA",
			x"0000" when x"87EB",
			x"0000" when x"87EC",
			x"0000" when x"87ED",
			x"0000" when x"87EE",
			x"0000" when x"87EF",
			x"0000" when x"87F0",
			x"0000" when x"87F1",
			x"0000" when x"87F2",
			x"0000" when x"87F3",
			x"0000" when x"87F4",
			x"0000" when x"87F5",
			x"0000" when x"87F6",
			x"0000" when x"87F7",
			x"0000" when x"87F8",
			x"0000" when x"87F9",
			x"0000" when x"87FA",
			x"0000" when x"87FB",
			x"0000" when x"87FC",
			x"0000" when x"87FD",
			x"0000" when x"87FE",
			x"0000" when x"87FF",
			x"0000" when x"8800",
			x"0000" when x"8801",
			x"0000" when x"8802",
			x"0000" when x"8803",
			x"0000" when x"8804",
			x"0000" when x"8805",
			x"0000" when x"8806",
			x"0000" when x"8807",
			x"0000" when x"8808",
			x"0000" when x"8809",
			x"0000" when x"880A",
			x"0000" when x"880B",
			x"0000" when x"880C",
			x"0000" when x"880D",
			x"0000" when x"880E",
			x"0000" when x"880F",
			x"0000" when x"8810",
			x"0000" when x"8811",
			x"0000" when x"8812",
			x"0000" when x"8813",
			x"0000" when x"8814",
			x"0000" when x"8815",
			x"0000" when x"8816",
			x"0000" when x"8817",
			x"0000" when x"8818",
			x"0000" when x"8819",
			x"0000" when x"881A",
			x"0000" when x"881B",
			x"0000" when x"881C",
			x"0000" when x"881D",
			x"0000" when x"881E",
			x"0000" when x"881F",
			x"0000" when x"8820",
			x"0000" when x"8821",
			x"0000" when x"8822",
			x"0000" when x"8823",
			x"0000" when x"8824",
			x"0000" when x"8825",
			x"0000" when x"8826",
			x"0000" when x"8827",
			x"0000" when x"8828",
			x"0000" when x"8829",
			x"0000" when x"882A",
			x"0000" when x"882B",
			x"0000" when x"882C",
			x"0000" when x"882D",
			x"0000" when x"882E",
			x"0000" when x"882F",
			x"0000" when x"8830",
			x"0000" when x"8831",
			x"0000" when x"8832",
			x"0000" when x"8833",
			x"0000" when x"8834",
			x"0000" when x"8835",
			x"0000" when x"8836",
			x"0000" when x"8837",
			x"0000" when x"8838",
			x"0000" when x"8839",
			x"0000" when x"883A",
			x"0000" when x"883B",
			x"0000" when x"883C",
			x"0000" when x"883D",
			x"0000" when x"883E",
			x"0000" when x"883F",
			x"0000" when x"8840",
			x"0000" when x"8841",
			x"0000" when x"8842",
			x"0000" when x"8843",
			x"0000" when x"8844",
			x"0000" when x"8845",
			x"0000" when x"8846",
			x"0000" when x"8847",
			x"0000" when x"8848",
			x"0000" when x"8849",
			x"0000" when x"884A",
			x"0000" when x"884B",
			x"0000" when x"884C",
			x"0000" when x"884D",
			x"0000" when x"884E",
			x"0000" when x"884F",
			x"0000" when x"8850",
			x"0000" when x"8851",
			x"0000" when x"8852",
			x"0000" when x"8853",
			x"0000" when x"8854",
			x"0000" when x"8855",
			x"0000" when x"8856",
			x"0000" when x"8857",
			x"0000" when x"8858",
			x"0000" when x"8859",
			x"0000" when x"885A",
			x"0000" when x"885B",
			x"0000" when x"885C",
			x"0000" when x"885D",
			x"0000" when x"885E",
			x"0000" when x"885F",
			x"0000" when x"8860",
			x"0000" when x"8861",
			x"0000" when x"8862",
			x"0000" when x"8863",
			x"0000" when x"8864",
			x"0000" when x"8865",
			x"0000" when x"8866",
			x"0000" when x"8867",
			x"0000" when x"8868",
			x"0000" when x"8869",
			x"0000" when x"886A",
			x"0000" when x"886B",
			x"0000" when x"886C",
			x"0000" when x"886D",
			x"0000" when x"886E",
			x"0000" when x"886F",
			x"0000" when x"8870",
			x"0000" when x"8871",
			x"0000" when x"8872",
			x"0000" when x"8873",
			x"0000" when x"8874",
			x"0000" when x"8875",
			x"0000" when x"8876",
			x"0000" when x"8877",
			x"0000" when x"8878",
			x"0000" when x"8879",
			x"0000" when x"887A",
			x"0000" when x"887B",
			x"0000" when x"887C",
			x"0000" when x"887D",
			x"0000" when x"887E",
			x"0000" when x"887F",
			x"0000" when x"8880",
			x"0000" when x"8881",
			x"0000" when x"8882",
			x"0000" when x"8883",
			x"0000" when x"8884",
			x"0000" when x"8885",
			x"0000" when x"8886",
			x"0000" when x"8887",
			x"0000" when x"8888",
			x"0000" when x"8889",
			x"0000" when x"888A",
			x"0000" when x"888B",
			x"0000" when x"888C",
			x"0000" when x"888D",
			x"0000" when x"888E",
			x"0000" when x"888F",
			x"0000" when x"8890",
			x"0000" when x"8891",
			x"0000" when x"8892",
			x"0000" when x"8893",
			x"0000" when x"8894",
			x"0000" when x"8895",
			x"0000" when x"8896",
			x"0000" when x"8897",
			x"0000" when x"8898",
			x"0000" when x"8899",
			x"0000" when x"889A",
			x"0000" when x"889B",
			x"0000" when x"889C",
			x"0000" when x"889D",
			x"0000" when x"889E",
			x"0000" when x"889F",
			x"0000" when x"88A0",
			x"0000" when x"88A1",
			x"0000" when x"88A2",
			x"0000" when x"88A3",
			x"0000" when x"88A4",
			x"0000" when x"88A5",
			x"0000" when x"88A6",
			x"0000" when x"88A7",
			x"0000" when x"88A8",
			x"0000" when x"88A9",
			x"0000" when x"88AA",
			x"0000" when x"88AB",
			x"0000" when x"88AC",
			x"0000" when x"88AD",
			x"0000" when x"88AE",
			x"0000" when x"88AF",
			x"0000" when x"88B0",
			x"0000" when x"88B1",
			x"0000" when x"88B2",
			x"0000" when x"88B3",
			x"0000" when x"88B4",
			x"0000" when x"88B5",
			x"0000" when x"88B6",
			x"0000" when x"88B7",
			x"0000" when x"88B8",
			x"0000" when x"88B9",
			x"0000" when x"88BA",
			x"0000" when x"88BB",
			x"0000" when x"88BC",
			x"0000" when x"88BD",
			x"0000" when x"88BE",
			x"0000" when x"88BF",
			x"0000" when x"88C0",
			x"0000" when x"88C1",
			x"0000" when x"88C2",
			x"0000" when x"88C3",
			x"0000" when x"88C4",
			x"0000" when x"88C5",
			x"0000" when x"88C6",
			x"0000" when x"88C7",
			x"0000" when x"88C8",
			x"0000" when x"88C9",
			x"0000" when x"88CA",
			x"0000" when x"88CB",
			x"0000" when x"88CC",
			x"0000" when x"88CD",
			x"0000" when x"88CE",
			x"0000" when x"88CF",
			x"0000" when x"88D0",
			x"0000" when x"88D1",
			x"0000" when x"88D2",
			x"0000" when x"88D3",
			x"0000" when x"88D4",
			x"0000" when x"88D5",
			x"0000" when x"88D6",
			x"0000" when x"88D7",
			x"0000" when x"88D8",
			x"0000" when x"88D9",
			x"0000" when x"88DA",
			x"0000" when x"88DB",
			x"0000" when x"88DC",
			x"0000" when x"88DD",
			x"0000" when x"88DE",
			x"0000" when x"88DF",
			x"0000" when x"88E0",
			x"0000" when x"88E1",
			x"0000" when x"88E2",
			x"0000" when x"88E3",
			x"0000" when x"88E4",
			x"0000" when x"88E5",
			x"0000" when x"88E6",
			x"0000" when x"88E7",
			x"0000" when x"88E8",
			x"0000" when x"88E9",
			x"0000" when x"88EA",
			x"0000" when x"88EB",
			x"0000" when x"88EC",
			x"0000" when x"88ED",
			x"0000" when x"88EE",
			x"0000" when x"88EF",
			x"0000" when x"88F0",
			x"0000" when x"88F1",
			x"0000" when x"88F2",
			x"0000" when x"88F3",
			x"0000" when x"88F4",
			x"0000" when x"88F5",
			x"0000" when x"88F6",
			x"0000" when x"88F7",
			x"0000" when x"88F8",
			x"0000" when x"88F9",
			x"0000" when x"88FA",
			x"0000" when x"88FB",
			x"0000" when x"88FC",
			x"0000" when x"88FD",
			x"0000" when x"88FE",
			x"0000" when x"88FF",
			x"0000" when x"8900",
			x"0000" when x"8901",
			x"0000" when x"8902",
			x"0000" when x"8903",
			x"0000" when x"8904",
			x"0000" when x"8905",
			x"0000" when x"8906",
			x"0000" when x"8907",
			x"0000" when x"8908",
			x"0000" when x"8909",
			x"0000" when x"890A",
			x"0000" when x"890B",
			x"0000" when x"890C",
			x"0000" when x"890D",
			x"0000" when x"890E",
			x"0000" when x"890F",
			x"0000" when x"8910",
			x"0000" when x"8911",
			x"0000" when x"8912",
			x"0000" when x"8913",
			x"0000" when x"8914",
			x"0000" when x"8915",
			x"0000" when x"8916",
			x"0000" when x"8917",
			x"0000" when x"8918",
			x"0000" when x"8919",
			x"0000" when x"891A",
			x"0000" when x"891B",
			x"0000" when x"891C",
			x"0000" when x"891D",
			x"0000" when x"891E",
			x"0000" when x"891F",
			x"0000" when x"8920",
			x"0000" when x"8921",
			x"0000" when x"8922",
			x"0000" when x"8923",
			x"0000" when x"8924",
			x"0000" when x"8925",
			x"0000" when x"8926",
			x"0000" when x"8927",
			x"0000" when x"8928",
			x"0000" when x"8929",
			x"0000" when x"892A",
			x"0000" when x"892B",
			x"0000" when x"892C",
			x"0000" when x"892D",
			x"0000" when x"892E",
			x"0000" when x"892F",
			x"0000" when x"8930",
			x"0000" when x"8931",
			x"0000" when x"8932",
			x"0000" when x"8933",
			x"0000" when x"8934",
			x"0000" when x"8935",
			x"0000" when x"8936",
			x"0000" when x"8937",
			x"0000" when x"8938",
			x"0000" when x"8939",
			x"0000" when x"893A",
			x"0000" when x"893B",
			x"0000" when x"893C",
			x"0000" when x"893D",
			x"0000" when x"893E",
			x"0000" when x"893F",
			x"0000" when x"8940",
			x"0000" when x"8941",
			x"0000" when x"8942",
			x"0000" when x"8943",
			x"0000" when x"8944",
			x"0000" when x"8945",
			x"0000" when x"8946",
			x"0000" when x"8947",
			x"0000" when x"8948",
			x"0000" when x"8949",
			x"0000" when x"894A",
			x"0000" when x"894B",
			x"0000" when x"894C",
			x"0000" when x"894D",
			x"0000" when x"894E",
			x"0000" when x"894F",
			x"0000" when x"8950",
			x"0000" when x"8951",
			x"0000" when x"8952",
			x"0000" when x"8953",
			x"0000" when x"8954",
			x"0000" when x"8955",
			x"0000" when x"8956",
			x"0000" when x"8957",
			x"0000" when x"8958",
			x"0000" when x"8959",
			x"0000" when x"895A",
			x"0000" when x"895B",
			x"0000" when x"895C",
			x"0000" when x"895D",
			x"0000" when x"895E",
			x"0000" when x"895F",
			x"0000" when x"8960",
			x"0000" when x"8961",
			x"0000" when x"8962",
			x"0000" when x"8963",
			x"0000" when x"8964",
			x"0000" when x"8965",
			x"0000" when x"8966",
			x"0000" when x"8967",
			x"0000" when x"8968",
			x"0000" when x"8969",
			x"0000" when x"896A",
			x"0000" when x"896B",
			x"0000" when x"896C",
			x"0000" when x"896D",
			x"0000" when x"896E",
			x"0000" when x"896F",
			x"0000" when x"8970",
			x"0000" when x"8971",
			x"0000" when x"8972",
			x"0000" when x"8973",
			x"0000" when x"8974",
			x"0000" when x"8975",
			x"0000" when x"8976",
			x"0000" when x"8977",
			x"0000" when x"8978",
			x"0000" when x"8979",
			x"0000" when x"897A",
			x"0000" when x"897B",
			x"0000" when x"897C",
			x"0000" when x"897D",
			x"0000" when x"897E",
			x"0000" when x"897F",
			x"0000" when x"8980",
			x"0000" when x"8981",
			x"0000" when x"8982",
			x"0000" when x"8983",
			x"0000" when x"8984",
			x"0000" when x"8985",
			x"0000" when x"8986",
			x"0000" when x"8987",
			x"0000" when x"8988",
			x"0000" when x"8989",
			x"0000" when x"898A",
			x"0000" when x"898B",
			x"0000" when x"898C",
			x"0000" when x"898D",
			x"0000" when x"898E",
			x"0000" when x"898F",
			x"0000" when x"8990",
			x"0000" when x"8991",
			x"0000" when x"8992",
			x"0000" when x"8993",
			x"0000" when x"8994",
			x"0000" when x"8995",
			x"0000" when x"8996",
			x"0000" when x"8997",
			x"0000" when x"8998",
			x"0000" when x"8999",
			x"0000" when x"899A",
			x"0000" when x"899B",
			x"0000" when x"899C",
			x"0000" when x"899D",
			x"0000" when x"899E",
			x"0000" when x"899F",
			x"0000" when x"89A0",
			x"0000" when x"89A1",
			x"0000" when x"89A2",
			x"0000" when x"89A3",
			x"0000" when x"89A4",
			x"0000" when x"89A5",
			x"0000" when x"89A6",
			x"0000" when x"89A7",
			x"0000" when x"89A8",
			x"0000" when x"89A9",
			x"0000" when x"89AA",
			x"0000" when x"89AB",
			x"0000" when x"89AC",
			x"0000" when x"89AD",
			x"0000" when x"89AE",
			x"0000" when x"89AF",
			x"0000" when x"89B0",
			x"0000" when x"89B1",
			x"0000" when x"89B2",
			x"0000" when x"89B3",
			x"0000" when x"89B4",
			x"0000" when x"89B5",
			x"0000" when x"89B6",
			x"0000" when x"89B7",
			x"0000" when x"89B8",
			x"0000" when x"89B9",
			x"0000" when x"89BA",
			x"0000" when x"89BB",
			x"0000" when x"89BC",
			x"0000" when x"89BD",
			x"0000" when x"89BE",
			x"0000" when x"89BF",
			x"0000" when x"89C0",
			x"0000" when x"89C1",
			x"0000" when x"89C2",
			x"0000" when x"89C3",
			x"0000" when x"89C4",
			x"0000" when x"89C5",
			x"0000" when x"89C6",
			x"0000" when x"89C7",
			x"0000" when x"89C8",
			x"0000" when x"89C9",
			x"0000" when x"89CA",
			x"0000" when x"89CB",
			x"0000" when x"89CC",
			x"0000" when x"89CD",
			x"0000" when x"89CE",
			x"0000" when x"89CF",
			x"0000" when x"89D0",
			x"0000" when x"89D1",
			x"0000" when x"89D2",
			x"0000" when x"89D3",
			x"0000" when x"89D4",
			x"0000" when x"89D5",
			x"0000" when x"89D6",
			x"0000" when x"89D7",
			x"0000" when x"89D8",
			x"0000" when x"89D9",
			x"0000" when x"89DA",
			x"0000" when x"89DB",
			x"0000" when x"89DC",
			x"0000" when x"89DD",
			x"0000" when x"89DE",
			x"0000" when x"89DF",
			x"0000" when x"89E0",
			x"0000" when x"89E1",
			x"0000" when x"89E2",
			x"0000" when x"89E3",
			x"0000" when x"89E4",
			x"0000" when x"89E5",
			x"0000" when x"89E6",
			x"0000" when x"89E7",
			x"0000" when x"89E8",
			x"0000" when x"89E9",
			x"0000" when x"89EA",
			x"0000" when x"89EB",
			x"0000" when x"89EC",
			x"0000" when x"89ED",
			x"0000" when x"89EE",
			x"0000" when x"89EF",
			x"0000" when x"89F0",
			x"0000" when x"89F1",
			x"0000" when x"89F2",
			x"0000" when x"89F3",
			x"0000" when x"89F4",
			x"0000" when x"89F5",
			x"0000" when x"89F6",
			x"0000" when x"89F7",
			x"0000" when x"89F8",
			x"0000" when x"89F9",
			x"0000" when x"89FA",
			x"0000" when x"89FB",
			x"0000" when x"89FC",
			x"0000" when x"89FD",
			x"0000" when x"89FE",
			x"0000" when x"89FF",
			x"0000" when x"8A00",
			x"0000" when x"8A01",
			x"0000" when x"8A02",
			x"0000" when x"8A03",
			x"0000" when x"8A04",
			x"0000" when x"8A05",
			x"0000" when x"8A06",
			x"0000" when x"8A07",
			x"0000" when x"8A08",
			x"0000" when x"8A09",
			x"0000" when x"8A0A",
			x"0000" when x"8A0B",
			x"0000" when x"8A0C",
			x"0000" when x"8A0D",
			x"0000" when x"8A0E",
			x"0000" when x"8A0F",
			x"0000" when x"8A10",
			x"0000" when x"8A11",
			x"0000" when x"8A12",
			x"0000" when x"8A13",
			x"0000" when x"8A14",
			x"0000" when x"8A15",
			x"0000" when x"8A16",
			x"0000" when x"8A17",
			x"0000" when x"8A18",
			x"0000" when x"8A19",
			x"0000" when x"8A1A",
			x"0000" when x"8A1B",
			x"0000" when x"8A1C",
			x"0000" when x"8A1D",
			x"0000" when x"8A1E",
			x"0000" when x"8A1F",
			x"0000" when x"8A20",
			x"0000" when x"8A21",
			x"0000" when x"8A22",
			x"0000" when x"8A23",
			x"0000" when x"8A24",
			x"0000" when x"8A25",
			x"0000" when x"8A26",
			x"0000" when x"8A27",
			x"0000" when x"8A28",
			x"0000" when x"8A29",
			x"0000" when x"8A2A",
			x"0000" when x"8A2B",
			x"0000" when x"8A2C",
			x"0000" when x"8A2D",
			x"0000" when x"8A2E",
			x"0000" when x"8A2F",
			x"0000" when x"8A30",
			x"0000" when x"8A31",
			x"0000" when x"8A32",
			x"0000" when x"8A33",
			x"0000" when x"8A34",
			x"0000" when x"8A35",
			x"0000" when x"8A36",
			x"0000" when x"8A37",
			x"0000" when x"8A38",
			x"0000" when x"8A39",
			x"0000" when x"8A3A",
			x"0000" when x"8A3B",
			x"0000" when x"8A3C",
			x"0000" when x"8A3D",
			x"0000" when x"8A3E",
			x"0000" when x"8A3F",
			x"0000" when x"8A40",
			x"0000" when x"8A41",
			x"0000" when x"8A42",
			x"0000" when x"8A43",
			x"0000" when x"8A44",
			x"0000" when x"8A45",
			x"0000" when x"8A46",
			x"0000" when x"8A47",
			x"0000" when x"8A48",
			x"0000" when x"8A49",
			x"0000" when x"8A4A",
			x"0000" when x"8A4B",
			x"0000" when x"8A4C",
			x"0000" when x"8A4D",
			x"0000" when x"8A4E",
			x"0000" when x"8A4F",
			x"0000" when x"8A50",
			x"0000" when x"8A51",
			x"0000" when x"8A52",
			x"0000" when x"8A53",
			x"0000" when x"8A54",
			x"0000" when x"8A55",
			x"0000" when x"8A56",
			x"0000" when x"8A57",
			x"0000" when x"8A58",
			x"0000" when x"8A59",
			x"0000" when x"8A5A",
			x"0000" when x"8A5B",
			x"0000" when x"8A5C",
			x"0000" when x"8A5D",
			x"0000" when x"8A5E",
			x"0000" when x"8A5F",
			x"0000" when x"8A60",
			x"0000" when x"8A61",
			x"0000" when x"8A62",
			x"0000" when x"8A63",
			x"0000" when x"8A64",
			x"0000" when x"8A65",
			x"0000" when x"8A66",
			x"0000" when x"8A67",
			x"0000" when x"8A68",
			x"0000" when x"8A69",
			x"0000" when x"8A6A",
			x"0000" when x"8A6B",
			x"0000" when x"8A6C",
			x"0000" when x"8A6D",
			x"0000" when x"8A6E",
			x"0000" when x"8A6F",
			x"0000" when x"8A70",
			x"0000" when x"8A71",
			x"0000" when x"8A72",
			x"0000" when x"8A73",
			x"0000" when x"8A74",
			x"0000" when x"8A75",
			x"0000" when x"8A76",
			x"0000" when x"8A77",
			x"0000" when x"8A78",
			x"0000" when x"8A79",
			x"0000" when x"8A7A",
			x"0000" when x"8A7B",
			x"0000" when x"8A7C",
			x"0000" when x"8A7D",
			x"0000" when x"8A7E",
			x"0000" when x"8A7F",
			x"0000" when x"8A80",
			x"0000" when x"8A81",
			x"0000" when x"8A82",
			x"0000" when x"8A83",
			x"0000" when x"8A84",
			x"0000" when x"8A85",
			x"0000" when x"8A86",
			x"0000" when x"8A87",
			x"0000" when x"8A88",
			x"0000" when x"8A89",
			x"0000" when x"8A8A",
			x"0000" when x"8A8B",
			x"0000" when x"8A8C",
			x"0000" when x"8A8D",
			x"0000" when x"8A8E",
			x"0000" when x"8A8F",
			x"0000" when x"8A90",
			x"0000" when x"8A91",
			x"0000" when x"8A92",
			x"0000" when x"8A93",
			x"0000" when x"8A94",
			x"0000" when x"8A95",
			x"0000" when x"8A96",
			x"0000" when x"8A97",
			x"0000" when x"8A98",
			x"0000" when x"8A99",
			x"0000" when x"8A9A",
			x"0000" when x"8A9B",
			x"0000" when x"8A9C",
			x"0000" when x"8A9D",
			x"0000" when x"8A9E",
			x"0000" when x"8A9F",
			x"0000" when x"8AA0",
			x"0000" when x"8AA1",
			x"0000" when x"8AA2",
			x"0000" when x"8AA3",
			x"0000" when x"8AA4",
			x"0000" when x"8AA5",
			x"0000" when x"8AA6",
			x"0000" when x"8AA7",
			x"0000" when x"8AA8",
			x"0000" when x"8AA9",
			x"0000" when x"8AAA",
			x"0000" when x"8AAB",
			x"0000" when x"8AAC",
			x"0000" when x"8AAD",
			x"0000" when x"8AAE",
			x"0000" when x"8AAF",
			x"0000" when x"8AB0",
			x"0000" when x"8AB1",
			x"0000" when x"8AB2",
			x"0000" when x"8AB3",
			x"0000" when x"8AB4",
			x"0000" when x"8AB5",
			x"0000" when x"8AB6",
			x"0000" when x"8AB7",
			x"0000" when x"8AB8",
			x"0000" when x"8AB9",
			x"0000" when x"8ABA",
			x"0000" when x"8ABB",
			x"0000" when x"8ABC",
			x"0000" when x"8ABD",
			x"0000" when x"8ABE",
			x"0000" when x"8ABF",
			x"0000" when x"8AC0",
			x"0000" when x"8AC1",
			x"0000" when x"8AC2",
			x"0000" when x"8AC3",
			x"0000" when x"8AC4",
			x"0000" when x"8AC5",
			x"0000" when x"8AC6",
			x"0000" when x"8AC7",
			x"0000" when x"8AC8",
			x"0000" when x"8AC9",
			x"0000" when x"8ACA",
			x"0000" when x"8ACB",
			x"0000" when x"8ACC",
			x"0000" when x"8ACD",
			x"0000" when x"8ACE",
			x"0000" when x"8ACF",
			x"0000" when x"8AD0",
			x"0000" when x"8AD1",
			x"0000" when x"8AD2",
			x"0000" when x"8AD3",
			x"0000" when x"8AD4",
			x"0000" when x"8AD5",
			x"0000" when x"8AD6",
			x"0000" when x"8AD7",
			x"0000" when x"8AD8",
			x"0000" when x"8AD9",
			x"0000" when x"8ADA",
			x"0000" when x"8ADB",
			x"0000" when x"8ADC",
			x"0000" when x"8ADD",
			x"0000" when x"8ADE",
			x"0000" when x"8ADF",
			x"0000" when x"8AE0",
			x"0000" when x"8AE1",
			x"0000" when x"8AE2",
			x"0000" when x"8AE3",
			x"0000" when x"8AE4",
			x"0000" when x"8AE5",
			x"0000" when x"8AE6",
			x"0000" when x"8AE7",
			x"0000" when x"8AE8",
			x"0000" when x"8AE9",
			x"0000" when x"8AEA",
			x"0000" when x"8AEB",
			x"0000" when x"8AEC",
			x"0000" when x"8AED",
			x"0000" when x"8AEE",
			x"0000" when x"8AEF",
			x"0000" when x"8AF0",
			x"0000" when x"8AF1",
			x"0000" when x"8AF2",
			x"0000" when x"8AF3",
			x"0000" when x"8AF4",
			x"0000" when x"8AF5",
			x"0000" when x"8AF6",
			x"0000" when x"8AF7",
			x"0000" when x"8AF8",
			x"0000" when x"8AF9",
			x"0000" when x"8AFA",
			x"0000" when x"8AFB",
			x"0000" when x"8AFC",
			x"0000" when x"8AFD",
			x"0000" when x"8AFE",
			x"0000" when x"8AFF",
			x"0000" when x"8B00",
			x"0000" when x"8B01",
			x"0000" when x"8B02",
			x"0000" when x"8B03",
			x"0000" when x"8B04",
			x"0000" when x"8B05",
			x"0000" when x"8B06",
			x"0000" when x"8B07",
			x"0000" when x"8B08",
			x"0000" when x"8B09",
			x"0000" when x"8B0A",
			x"0000" when x"8B0B",
			x"0000" when x"8B0C",
			x"0000" when x"8B0D",
			x"0000" when x"8B0E",
			x"0000" when x"8B0F",
			x"0000" when x"8B10",
			x"0000" when x"8B11",
			x"0000" when x"8B12",
			x"0000" when x"8B13",
			x"0000" when x"8B14",
			x"0000" when x"8B15",
			x"0000" when x"8B16",
			x"0000" when x"8B17",
			x"0000" when x"8B18",
			x"0000" when x"8B19",
			x"0000" when x"8B1A",
			x"0000" when x"8B1B",
			x"0000" when x"8B1C",
			x"0000" when x"8B1D",
			x"0000" when x"8B1E",
			x"0000" when x"8B1F",
			x"0000" when x"8B20",
			x"0000" when x"8B21",
			x"0000" when x"8B22",
			x"0000" when x"8B23",
			x"0000" when x"8B24",
			x"0000" when x"8B25",
			x"0000" when x"8B26",
			x"0000" when x"8B27",
			x"0000" when x"8B28",
			x"0000" when x"8B29",
			x"0000" when x"8B2A",
			x"0000" when x"8B2B",
			x"0000" when x"8B2C",
			x"0000" when x"8B2D",
			x"0000" when x"8B2E",
			x"0000" when x"8B2F",
			x"0000" when x"8B30",
			x"0000" when x"8B31",
			x"0000" when x"8B32",
			x"0000" when x"8B33",
			x"0000" when x"8B34",
			x"0000" when x"8B35",
			x"0000" when x"8B36",
			x"0000" when x"8B37",
			x"0000" when x"8B38",
			x"0000" when x"8B39",
			x"0000" when x"8B3A",
			x"0000" when x"8B3B",
			x"0000" when x"8B3C",
			x"0000" when x"8B3D",
			x"0000" when x"8B3E",
			x"0000" when x"8B3F",
			x"0000" when x"8B40",
			x"0000" when x"8B41",
			x"0000" when x"8B42",
			x"0000" when x"8B43",
			x"0000" when x"8B44",
			x"0000" when x"8B45",
			x"0000" when x"8B46",
			x"0000" when x"8B47",
			x"0000" when x"8B48",
			x"0000" when x"8B49",
			x"0000" when x"8B4A",
			x"0000" when x"8B4B",
			x"0000" when x"8B4C",
			x"0000" when x"8B4D",
			x"0000" when x"8B4E",
			x"0000" when x"8B4F",
			x"0000" when x"8B50",
			x"0000" when x"8B51",
			x"0000" when x"8B52",
			x"0000" when x"8B53",
			x"0000" when x"8B54",
			x"0000" when x"8B55",
			x"0000" when x"8B56",
			x"0000" when x"8B57",
			x"0000" when x"8B58",
			x"0000" when x"8B59",
			x"0000" when x"8B5A",
			x"0000" when x"8B5B",
			x"0000" when x"8B5C",
			x"0000" when x"8B5D",
			x"0000" when x"8B5E",
			x"0000" when x"8B5F",
			x"0000" when x"8B60",
			x"0000" when x"8B61",
			x"0000" when x"8B62",
			x"0000" when x"8B63",
			x"0000" when x"8B64",
			x"0000" when x"8B65",
			x"0000" when x"8B66",
			x"0000" when x"8B67",
			x"0000" when x"8B68",
			x"0000" when x"8B69",
			x"0000" when x"8B6A",
			x"0000" when x"8B6B",
			x"0000" when x"8B6C",
			x"0000" when x"8B6D",
			x"0000" when x"8B6E",
			x"0000" when x"8B6F",
			x"0000" when x"8B70",
			x"0000" when x"8B71",
			x"0000" when x"8B72",
			x"0000" when x"8B73",
			x"0000" when x"8B74",
			x"0000" when x"8B75",
			x"0000" when x"8B76",
			x"0000" when x"8B77",
			x"0000" when x"8B78",
			x"0000" when x"8B79",
			x"0000" when x"8B7A",
			x"0000" when x"8B7B",
			x"0000" when x"8B7C",
			x"0000" when x"8B7D",
			x"0000" when x"8B7E",
			x"0000" when x"8B7F",
			x"0000" when x"8B80",
			x"0000" when x"8B81",
			x"0000" when x"8B82",
			x"0000" when x"8B83",
			x"0000" when x"8B84",
			x"0000" when x"8B85",
			x"0000" when x"8B86",
			x"0000" when x"8B87",
			x"0000" when x"8B88",
			x"0000" when x"8B89",
			x"0000" when x"8B8A",
			x"0000" when x"8B8B",
			x"0000" when x"8B8C",
			x"0000" when x"8B8D",
			x"0000" when x"8B8E",
			x"0000" when x"8B8F",
			x"0000" when x"8B90",
			x"0000" when x"8B91",
			x"0000" when x"8B92",
			x"0000" when x"8B93",
			x"0000" when x"8B94",
			x"0000" when x"8B95",
			x"0000" when x"8B96",
			x"0000" when x"8B97",
			x"0000" when x"8B98",
			x"0000" when x"8B99",
			x"0000" when x"8B9A",
			x"0000" when x"8B9B",
			x"0000" when x"8B9C",
			x"0000" when x"8B9D",
			x"0000" when x"8B9E",
			x"0000" when x"8B9F",
			x"0000" when x"8BA0",
			x"0000" when x"8BA1",
			x"0000" when x"8BA2",
			x"0000" when x"8BA3",
			x"0000" when x"8BA4",
			x"0000" when x"8BA5",
			x"0000" when x"8BA6",
			x"0000" when x"8BA7",
			x"0000" when x"8BA8",
			x"0000" when x"8BA9",
			x"0000" when x"8BAA",
			x"0000" when x"8BAB",
			x"0000" when x"8BAC",
			x"0000" when x"8BAD",
			x"0000" when x"8BAE",
			x"0000" when x"8BAF",
			x"0000" when x"8BB0",
			x"0000" when x"8BB1",
			x"0000" when x"8BB2",
			x"0000" when x"8BB3",
			x"0000" when x"8BB4",
			x"0000" when x"8BB5",
			x"0000" when x"8BB6",
			x"0000" when x"8BB7",
			x"0000" when x"8BB8",
			x"0000" when x"8BB9",
			x"0000" when x"8BBA",
			x"0000" when x"8BBB",
			x"0000" when x"8BBC",
			x"0000" when x"8BBD",
			x"0000" when x"8BBE",
			x"0000" when x"8BBF",
			x"0000" when x"8BC0",
			x"0000" when x"8BC1",
			x"0000" when x"8BC2",
			x"0000" when x"8BC3",
			x"0000" when x"8BC4",
			x"0000" when x"8BC5",
			x"0000" when x"8BC6",
			x"0000" when x"8BC7",
			x"0000" when x"8BC8",
			x"0000" when x"8BC9",
			x"0000" when x"8BCA",
			x"0000" when x"8BCB",
			x"0000" when x"8BCC",
			x"0000" when x"8BCD",
			x"0000" when x"8BCE",
			x"0000" when x"8BCF",
			x"0000" when x"8BD0",
			x"0000" when x"8BD1",
			x"0000" when x"8BD2",
			x"0000" when x"8BD3",
			x"0000" when x"8BD4",
			x"0000" when x"8BD5",
			x"0000" when x"8BD6",
			x"0000" when x"8BD7",
			x"0000" when x"8BD8",
			x"0000" when x"8BD9",
			x"0000" when x"8BDA",
			x"0000" when x"8BDB",
			x"0000" when x"8BDC",
			x"0000" when x"8BDD",
			x"0000" when x"8BDE",
			x"0000" when x"8BDF",
			x"0000" when x"8BE0",
			x"0000" when x"8BE1",
			x"0000" when x"8BE2",
			x"0000" when x"8BE3",
			x"0000" when x"8BE4",
			x"0000" when x"8BE5",
			x"0000" when x"8BE6",
			x"0000" when x"8BE7",
			x"0000" when x"8BE8",
			x"0000" when x"8BE9",
			x"0000" when x"8BEA",
			x"0000" when x"8BEB",
			x"0000" when x"8BEC",
			x"0000" when x"8BED",
			x"0000" when x"8BEE",
			x"0000" when x"8BEF",
			x"0000" when x"8BF0",
			x"0000" when x"8BF1",
			x"0000" when x"8BF2",
			x"0000" when x"8BF3",
			x"0000" when x"8BF4",
			x"0000" when x"8BF5",
			x"0000" when x"8BF6",
			x"0000" when x"8BF7",
			x"0000" when x"8BF8",
			x"0000" when x"8BF9",
			x"0000" when x"8BFA",
			x"0000" when x"8BFB",
			x"0000" when x"8BFC",
			x"0000" when x"8BFD",
			x"0000" when x"8BFE",
			x"0000" when x"8BFF",
			x"0000" when x"8C00",
			x"0000" when x"8C01",
			x"0000" when x"8C02",
			x"0000" when x"8C03",
			x"0000" when x"8C04",
			x"0000" when x"8C05",
			x"0000" when x"8C06",
			x"0000" when x"8C07",
			x"0000" when x"8C08",
			x"0000" when x"8C09",
			x"0000" when x"8C0A",
			x"0000" when x"8C0B",
			x"0000" when x"8C0C",
			x"0000" when x"8C0D",
			x"0000" when x"8C0E",
			x"0000" when x"8C0F",
			x"0000" when x"8C10",
			x"0000" when x"8C11",
			x"0000" when x"8C12",
			x"0000" when x"8C13",
			x"0000" when x"8C14",
			x"0000" when x"8C15",
			x"0000" when x"8C16",
			x"0000" when x"8C17",
			x"0000" when x"8C18",
			x"0000" when x"8C19",
			x"0000" when x"8C1A",
			x"0000" when x"8C1B",
			x"0000" when x"8C1C",
			x"0000" when x"8C1D",
			x"0000" when x"8C1E",
			x"0000" when x"8C1F",
			x"0000" when x"8C20",
			x"0000" when x"8C21",
			x"0000" when x"8C22",
			x"0000" when x"8C23",
			x"0000" when x"8C24",
			x"0000" when x"8C25",
			x"0000" when x"8C26",
			x"0000" when x"8C27",
			x"0000" when x"8C28",
			x"0000" when x"8C29",
			x"0000" when x"8C2A",
			x"0000" when x"8C2B",
			x"0000" when x"8C2C",
			x"0000" when x"8C2D",
			x"0000" when x"8C2E",
			x"0000" when x"8C2F",
			x"0000" when x"8C30",
			x"0000" when x"8C31",
			x"0000" when x"8C32",
			x"0000" when x"8C33",
			x"0000" when x"8C34",
			x"0000" when x"8C35",
			x"0000" when x"8C36",
			x"0000" when x"8C37",
			x"0000" when x"8C38",
			x"0000" when x"8C39",
			x"0000" when x"8C3A",
			x"0000" when x"8C3B",
			x"0000" when x"8C3C",
			x"0000" when x"8C3D",
			x"0000" when x"8C3E",
			x"0000" when x"8C3F",
			x"0000" when x"8C40",
			x"0000" when x"8C41",
			x"0000" when x"8C42",
			x"0000" when x"8C43",
			x"0000" when x"8C44",
			x"0000" when x"8C45",
			x"0000" when x"8C46",
			x"0000" when x"8C47",
			x"0000" when x"8C48",
			x"0000" when x"8C49",
			x"0000" when x"8C4A",
			x"0000" when x"8C4B",
			x"0000" when x"8C4C",
			x"0000" when x"8C4D",
			x"0000" when x"8C4E",
			x"0000" when x"8C4F",
			x"0000" when x"8C50",
			x"0000" when x"8C51",
			x"0000" when x"8C52",
			x"0000" when x"8C53",
			x"0000" when x"8C54",
			x"0000" when x"8C55",
			x"0000" when x"8C56",
			x"0000" when x"8C57",
			x"0000" when x"8C58",
			x"0000" when x"8C59",
			x"0000" when x"8C5A",
			x"0000" when x"8C5B",
			x"0000" when x"8C5C",
			x"0000" when x"8C5D",
			x"0000" when x"8C5E",
			x"0000" when x"8C5F",
			x"0000" when x"8C60",
			x"0000" when x"8C61",
			x"0000" when x"8C62",
			x"0000" when x"8C63",
			x"0000" when x"8C64",
			x"0000" when x"8C65",
			x"0000" when x"8C66",
			x"0000" when x"8C67",
			x"0000" when x"8C68",
			x"0000" when x"8C69",
			x"0000" when x"8C6A",
			x"0000" when x"8C6B",
			x"0000" when x"8C6C",
			x"0000" when x"8C6D",
			x"0000" when x"8C6E",
			x"0000" when x"8C6F",
			x"0000" when x"8C70",
			x"0000" when x"8C71",
			x"0000" when x"8C72",
			x"0000" when x"8C73",
			x"0000" when x"8C74",
			x"0000" when x"8C75",
			x"0000" when x"8C76",
			x"0000" when x"8C77",
			x"0000" when x"8C78",
			x"0000" when x"8C79",
			x"0000" when x"8C7A",
			x"0000" when x"8C7B",
			x"0000" when x"8C7C",
			x"0000" when x"8C7D",
			x"0000" when x"8C7E",
			x"0000" when x"8C7F",
			x"0000" when x"8C80",
			x"0000" when x"8C81",
			x"0000" when x"8C82",
			x"0000" when x"8C83",
			x"0000" when x"8C84",
			x"0000" when x"8C85",
			x"0000" when x"8C86",
			x"0000" when x"8C87",
			x"0000" when x"8C88",
			x"0000" when x"8C89",
			x"0000" when x"8C8A",
			x"0000" when x"8C8B",
			x"0000" when x"8C8C",
			x"0000" when x"8C8D",
			x"0000" when x"8C8E",
			x"0000" when x"8C8F",
			x"0000" when x"8C90",
			x"0000" when x"8C91",
			x"0000" when x"8C92",
			x"0000" when x"8C93",
			x"0000" when x"8C94",
			x"0000" when x"8C95",
			x"0000" when x"8C96",
			x"0000" when x"8C97",
			x"0000" when x"8C98",
			x"0000" when x"8C99",
			x"0000" when x"8C9A",
			x"0000" when x"8C9B",
			x"0000" when x"8C9C",
			x"0000" when x"8C9D",
			x"0000" when x"8C9E",
			x"0000" when x"8C9F",
			x"0000" when x"8CA0",
			x"0000" when x"8CA1",
			x"0000" when x"8CA2",
			x"0000" when x"8CA3",
			x"0000" when x"8CA4",
			x"0000" when x"8CA5",
			x"0000" when x"8CA6",
			x"0000" when x"8CA7",
			x"0000" when x"8CA8",
			x"0000" when x"8CA9",
			x"0000" when x"8CAA",
			x"0000" when x"8CAB",
			x"0000" when x"8CAC",
			x"0000" when x"8CAD",
			x"0000" when x"8CAE",
			x"0000" when x"8CAF",
			x"0000" when x"8CB0",
			x"0000" when x"8CB1",
			x"0000" when x"8CB2",
			x"0000" when x"8CB3",
			x"0000" when x"8CB4",
			x"0000" when x"8CB5",
			x"0000" when x"8CB6",
			x"0000" when x"8CB7",
			x"0000" when x"8CB8",
			x"0000" when x"8CB9",
			x"0000" when x"8CBA",
			x"0000" when x"8CBB",
			x"0000" when x"8CBC",
			x"0000" when x"8CBD",
			x"0000" when x"8CBE",
			x"0000" when x"8CBF",
			x"0000" when x"8CC0",
			x"0000" when x"8CC1",
			x"0000" when x"8CC2",
			x"0000" when x"8CC3",
			x"0000" when x"8CC4",
			x"0000" when x"8CC5",
			x"0000" when x"8CC6",
			x"0000" when x"8CC7",
			x"0000" when x"8CC8",
			x"0000" when x"8CC9",
			x"0000" when x"8CCA",
			x"0000" when x"8CCB",
			x"0000" when x"8CCC",
			x"0000" when x"8CCD",
			x"0000" when x"8CCE",
			x"0000" when x"8CCF",
			x"0000" when x"8CD0",
			x"0000" when x"8CD1",
			x"0000" when x"8CD2",
			x"0000" when x"8CD3",
			x"0000" when x"8CD4",
			x"0000" when x"8CD5",
			x"0000" when x"8CD6",
			x"0000" when x"8CD7",
			x"0000" when x"8CD8",
			x"0000" when x"8CD9",
			x"0000" when x"8CDA",
			x"0000" when x"8CDB",
			x"0000" when x"8CDC",
			x"0000" when x"8CDD",
			x"0000" when x"8CDE",
			x"0000" when x"8CDF",
			x"0000" when x"8CE0",
			x"0000" when x"8CE1",
			x"0000" when x"8CE2",
			x"0000" when x"8CE3",
			x"0000" when x"8CE4",
			x"0000" when x"8CE5",
			x"0000" when x"8CE6",
			x"0000" when x"8CE7",
			x"0000" when x"8CE8",
			x"0000" when x"8CE9",
			x"0000" when x"8CEA",
			x"0000" when x"8CEB",
			x"0000" when x"8CEC",
			x"0000" when x"8CED",
			x"0000" when x"8CEE",
			x"0000" when x"8CEF",
			x"0000" when x"8CF0",
			x"0000" when x"8CF1",
			x"0000" when x"8CF2",
			x"0000" when x"8CF3",
			x"0000" when x"8CF4",
			x"0000" when x"8CF5",
			x"0000" when x"8CF6",
			x"0000" when x"8CF7",
			x"0000" when x"8CF8",
			x"0000" when x"8CF9",
			x"0000" when x"8CFA",
			x"0000" when x"8CFB",
			x"0000" when x"8CFC",
			x"0000" when x"8CFD",
			x"0000" when x"8CFE",
			x"0000" when x"8CFF",
			x"0000" when x"8D00",
			x"0000" when x"8D01",
			x"0000" when x"8D02",
			x"0000" when x"8D03",
			x"0000" when x"8D04",
			x"0000" when x"8D05",
			x"0000" when x"8D06",
			x"0000" when x"8D07",
			x"0000" when x"8D08",
			x"0000" when x"8D09",
			x"0000" when x"8D0A",
			x"0000" when x"8D0B",
			x"0000" when x"8D0C",
			x"0000" when x"8D0D",
			x"0000" when x"8D0E",
			x"0000" when x"8D0F",
			x"0000" when x"8D10",
			x"0000" when x"8D11",
			x"0000" when x"8D12",
			x"0000" when x"8D13",
			x"0000" when x"8D14",
			x"0000" when x"8D15",
			x"0000" when x"8D16",
			x"0000" when x"8D17",
			x"0000" when x"8D18",
			x"0000" when x"8D19",
			x"0000" when x"8D1A",
			x"0000" when x"8D1B",
			x"0000" when x"8D1C",
			x"0000" when x"8D1D",
			x"0000" when x"8D1E",
			x"0000" when x"8D1F",
			x"0000" when x"8D20",
			x"0000" when x"8D21",
			x"0000" when x"8D22",
			x"0000" when x"8D23",
			x"0000" when x"8D24",
			x"0000" when x"8D25",
			x"0000" when x"8D26",
			x"0000" when x"8D27",
			x"0000" when x"8D28",
			x"0000" when x"8D29",
			x"0000" when x"8D2A",
			x"0000" when x"8D2B",
			x"0000" when x"8D2C",
			x"0000" when x"8D2D",
			x"0000" when x"8D2E",
			x"0000" when x"8D2F",
			x"0000" when x"8D30",
			x"0000" when x"8D31",
			x"0000" when x"8D32",
			x"0000" when x"8D33",
			x"0000" when x"8D34",
			x"0000" when x"8D35",
			x"0000" when x"8D36",
			x"0000" when x"8D37",
			x"0000" when x"8D38",
			x"0000" when x"8D39",
			x"0000" when x"8D3A",
			x"0000" when x"8D3B",
			x"0000" when x"8D3C",
			x"0000" when x"8D3D",
			x"0000" when x"8D3E",
			x"0000" when x"8D3F",
			x"0000" when x"8D40",
			x"0000" when x"8D41",
			x"0000" when x"8D42",
			x"0000" when x"8D43",
			x"0000" when x"8D44",
			x"0000" when x"8D45",
			x"0000" when x"8D46",
			x"0000" when x"8D47",
			x"0000" when x"8D48",
			x"0000" when x"8D49",
			x"0000" when x"8D4A",
			x"0000" when x"8D4B",
			x"0000" when x"8D4C",
			x"0000" when x"8D4D",
			x"0000" when x"8D4E",
			x"0000" when x"8D4F",
			x"0000" when x"8D50",
			x"0000" when x"8D51",
			x"0000" when x"8D52",
			x"0000" when x"8D53",
			x"0000" when x"8D54",
			x"0000" when x"8D55",
			x"0000" when x"8D56",
			x"0000" when x"8D57",
			x"0000" when x"8D58",
			x"0000" when x"8D59",
			x"0000" when x"8D5A",
			x"0000" when x"8D5B",
			x"0000" when x"8D5C",
			x"0000" when x"8D5D",
			x"0000" when x"8D5E",
			x"0000" when x"8D5F",
			x"0000" when x"8D60",
			x"0000" when x"8D61",
			x"0000" when x"8D62",
			x"0000" when x"8D63",
			x"0000" when x"8D64",
			x"0000" when x"8D65",
			x"0000" when x"8D66",
			x"0000" when x"8D67",
			x"0000" when x"8D68",
			x"0000" when x"8D69",
			x"0000" when x"8D6A",
			x"0000" when x"8D6B",
			x"0000" when x"8D6C",
			x"0000" when x"8D6D",
			x"0000" when x"8D6E",
			x"0000" when x"8D6F",
			x"0000" when x"8D70",
			x"0000" when x"8D71",
			x"0000" when x"8D72",
			x"0000" when x"8D73",
			x"0000" when x"8D74",
			x"0000" when x"8D75",
			x"0000" when x"8D76",
			x"0000" when x"8D77",
			x"0000" when x"8D78",
			x"0000" when x"8D79",
			x"0000" when x"8D7A",
			x"0000" when x"8D7B",
			x"0000" when x"8D7C",
			x"0000" when x"8D7D",
			x"0000" when x"8D7E",
			x"0000" when x"8D7F",
			x"0000" when x"8D80",
			x"0000" when x"8D81",
			x"0000" when x"8D82",
			x"0000" when x"8D83",
			x"0000" when x"8D84",
			x"0000" when x"8D85",
			x"0000" when x"8D86",
			x"0000" when x"8D87",
			x"0000" when x"8D88",
			x"0000" when x"8D89",
			x"0000" when x"8D8A",
			x"0000" when x"8D8B",
			x"0000" when x"8D8C",
			x"0000" when x"8D8D",
			x"0000" when x"8D8E",
			x"0000" when x"8D8F",
			x"0000" when x"8D90",
			x"0000" when x"8D91",
			x"0000" when x"8D92",
			x"0000" when x"8D93",
			x"0000" when x"8D94",
			x"0000" when x"8D95",
			x"0000" when x"8D96",
			x"0000" when x"8D97",
			x"0000" when x"8D98",
			x"0000" when x"8D99",
			x"0000" when x"8D9A",
			x"0000" when x"8D9B",
			x"0000" when x"8D9C",
			x"0000" when x"8D9D",
			x"0000" when x"8D9E",
			x"0000" when x"8D9F",
			x"0000" when x"8DA0",
			x"0000" when x"8DA1",
			x"0000" when x"8DA2",
			x"0000" when x"8DA3",
			x"0000" when x"8DA4",
			x"0000" when x"8DA5",
			x"0000" when x"8DA6",
			x"0000" when x"8DA7",
			x"0000" when x"8DA8",
			x"0000" when x"8DA9",
			x"0000" when x"8DAA",
			x"0000" when x"8DAB",
			x"0000" when x"8DAC",
			x"0000" when x"8DAD",
			x"0000" when x"8DAE",
			x"0000" when x"8DAF",
			x"0000" when x"8DB0",
			x"0000" when x"8DB1",
			x"0000" when x"8DB2",
			x"0000" when x"8DB3",
			x"0000" when x"8DB4",
			x"0000" when x"8DB5",
			x"0000" when x"8DB6",
			x"0000" when x"8DB7",
			x"0000" when x"8DB8",
			x"0000" when x"8DB9",
			x"0000" when x"8DBA",
			x"0000" when x"8DBB",
			x"0000" when x"8DBC",
			x"0000" when x"8DBD",
			x"0000" when x"8DBE",
			x"0000" when x"8DBF",
			x"0000" when x"8DC0",
			x"0000" when x"8DC1",
			x"0000" when x"8DC2",
			x"0000" when x"8DC3",
			x"0000" when x"8DC4",
			x"0000" when x"8DC5",
			x"0000" when x"8DC6",
			x"0000" when x"8DC7",
			x"0000" when x"8DC8",
			x"0000" when x"8DC9",
			x"0000" when x"8DCA",
			x"0000" when x"8DCB",
			x"0000" when x"8DCC",
			x"0000" when x"8DCD",
			x"0000" when x"8DCE",
			x"0000" when x"8DCF",
			x"0000" when x"8DD0",
			x"0000" when x"8DD1",
			x"0000" when x"8DD2",
			x"0000" when x"8DD3",
			x"0000" when x"8DD4",
			x"0000" when x"8DD5",
			x"0000" when x"8DD6",
			x"0000" when x"8DD7",
			x"0000" when x"8DD8",
			x"0000" when x"8DD9",
			x"0000" when x"8DDA",
			x"0000" when x"8DDB",
			x"0000" when x"8DDC",
			x"0000" when x"8DDD",
			x"0000" when x"8DDE",
			x"0000" when x"8DDF",
			x"0000" when x"8DE0",
			x"0000" when x"8DE1",
			x"0000" when x"8DE2",
			x"0000" when x"8DE3",
			x"0000" when x"8DE4",
			x"0000" when x"8DE5",
			x"0000" when x"8DE6",
			x"0000" when x"8DE7",
			x"0000" when x"8DE8",
			x"0000" when x"8DE9",
			x"0000" when x"8DEA",
			x"0000" when x"8DEB",
			x"0000" when x"8DEC",
			x"0000" when x"8DED",
			x"0000" when x"8DEE",
			x"0000" when x"8DEF",
			x"0000" when x"8DF0",
			x"0000" when x"8DF1",
			x"0000" when x"8DF2",
			x"0000" when x"8DF3",
			x"0000" when x"8DF4",
			x"0000" when x"8DF5",
			x"0000" when x"8DF6",
			x"0000" when x"8DF7",
			x"0000" when x"8DF8",
			x"0000" when x"8DF9",
			x"0000" when x"8DFA",
			x"0000" when x"8DFB",
			x"0000" when x"8DFC",
			x"0000" when x"8DFD",
			x"0000" when x"8DFE",
			x"0000" when x"8DFF",
			x"0000" when x"8E00",
			x"0000" when x"8E01",
			x"0000" when x"8E02",
			x"0000" when x"8E03",
			x"0000" when x"8E04",
			x"0000" when x"8E05",
			x"0000" when x"8E06",
			x"0000" when x"8E07",
			x"0000" when x"8E08",
			x"0000" when x"8E09",
			x"0000" when x"8E0A",
			x"0000" when x"8E0B",
			x"0000" when x"8E0C",
			x"0000" when x"8E0D",
			x"0000" when x"8E0E",
			x"0000" when x"8E0F",
			x"0000" when x"8E10",
			x"0000" when x"8E11",
			x"0000" when x"8E12",
			x"0000" when x"8E13",
			x"0000" when x"8E14",
			x"0000" when x"8E15",
			x"0000" when x"8E16",
			x"0000" when x"8E17",
			x"0000" when x"8E18",
			x"0000" when x"8E19",
			x"0000" when x"8E1A",
			x"0000" when x"8E1B",
			x"0000" when x"8E1C",
			x"0000" when x"8E1D",
			x"0000" when x"8E1E",
			x"0000" when x"8E1F",
			x"0000" when x"8E20",
			x"0000" when x"8E21",
			x"0000" when x"8E22",
			x"0000" when x"8E23",
			x"0000" when x"8E24",
			x"0000" when x"8E25",
			x"0000" when x"8E26",
			x"0000" when x"8E27",
			x"0000" when x"8E28",
			x"0000" when x"8E29",
			x"0000" when x"8E2A",
			x"0000" when x"8E2B",
			x"0000" when x"8E2C",
			x"0000" when x"8E2D",
			x"0000" when x"8E2E",
			x"0000" when x"8E2F",
			x"0000" when x"8E30",
			x"0000" when x"8E31",
			x"0000" when x"8E32",
			x"0000" when x"8E33",
			x"0000" when x"8E34",
			x"0000" when x"8E35",
			x"0000" when x"8E36",
			x"0000" when x"8E37",
			x"0000" when x"8E38",
			x"0000" when x"8E39",
			x"0000" when x"8E3A",
			x"0000" when x"8E3B",
			x"0000" when x"8E3C",
			x"0000" when x"8E3D",
			x"0000" when x"8E3E",
			x"0000" when x"8E3F",
			x"0000" when x"8E40",
			x"0000" when x"8E41",
			x"0000" when x"8E42",
			x"0000" when x"8E43",
			x"0000" when x"8E44",
			x"0000" when x"8E45",
			x"0000" when x"8E46",
			x"0000" when x"8E47",
			x"0000" when x"8E48",
			x"0000" when x"8E49",
			x"0000" when x"8E4A",
			x"0000" when x"8E4B",
			x"0000" when x"8E4C",
			x"0000" when x"8E4D",
			x"0000" when x"8E4E",
			x"0000" when x"8E4F",
			x"0000" when x"8E50",
			x"0000" when x"8E51",
			x"0000" when x"8E52",
			x"0000" when x"8E53",
			x"0000" when x"8E54",
			x"0000" when x"8E55",
			x"0000" when x"8E56",
			x"0000" when x"8E57",
			x"0000" when x"8E58",
			x"0000" when x"8E59",
			x"0000" when x"8E5A",
			x"0000" when x"8E5B",
			x"0000" when x"8E5C",
			x"0000" when x"8E5D",
			x"0000" when x"8E5E",
			x"0000" when x"8E5F",
			x"0000" when x"8E60",
			x"0000" when x"8E61",
			x"0000" when x"8E62",
			x"0000" when x"8E63",
			x"0000" when x"8E64",
			x"0000" when x"8E65",
			x"0000" when x"8E66",
			x"0000" when x"8E67",
			x"0000" when x"8E68",
			x"0000" when x"8E69",
			x"0000" when x"8E6A",
			x"0000" when x"8E6B",
			x"0000" when x"8E6C",
			x"0000" when x"8E6D",
			x"0000" when x"8E6E",
			x"0000" when x"8E6F",
			x"0000" when x"8E70",
			x"0000" when x"8E71",
			x"0000" when x"8E72",
			x"0000" when x"8E73",
			x"0000" when x"8E74",
			x"0000" when x"8E75",
			x"0000" when x"8E76",
			x"0000" when x"8E77",
			x"0000" when x"8E78",
			x"0000" when x"8E79",
			x"0000" when x"8E7A",
			x"0000" when x"8E7B",
			x"0000" when x"8E7C",
			x"0000" when x"8E7D",
			x"0000" when x"8E7E",
			x"0000" when x"8E7F",
			x"0000" when x"8E80",
			x"0000" when x"8E81",
			x"0000" when x"8E82",
			x"0000" when x"8E83",
			x"0000" when x"8E84",
			x"0000" when x"8E85",
			x"0000" when x"8E86",
			x"0000" when x"8E87",
			x"0000" when x"8E88",
			x"0000" when x"8E89",
			x"0000" when x"8E8A",
			x"0000" when x"8E8B",
			x"0000" when x"8E8C",
			x"0000" when x"8E8D",
			x"0000" when x"8E8E",
			x"0000" when x"8E8F",
			x"0000" when x"8E90",
			x"0000" when x"8E91",
			x"0000" when x"8E92",
			x"0000" when x"8E93",
			x"0000" when x"8E94",
			x"0000" when x"8E95",
			x"0000" when x"8E96",
			x"0000" when x"8E97",
			x"0000" when x"8E98",
			x"0000" when x"8E99",
			x"0000" when x"8E9A",
			x"0000" when x"8E9B",
			x"0000" when x"8E9C",
			x"0000" when x"8E9D",
			x"0000" when x"8E9E",
			x"0000" when x"8E9F",
			x"0000" when x"8EA0",
			x"0000" when x"8EA1",
			x"0000" when x"8EA2",
			x"0000" when x"8EA3",
			x"0000" when x"8EA4",
			x"0000" when x"8EA5",
			x"0000" when x"8EA6",
			x"0000" when x"8EA7",
			x"0000" when x"8EA8",
			x"0000" when x"8EA9",
			x"0000" when x"8EAA",
			x"0000" when x"8EAB",
			x"0000" when x"8EAC",
			x"0000" when x"8EAD",
			x"0000" when x"8EAE",
			x"0000" when x"8EAF",
			x"0000" when x"8EB0",
			x"0000" when x"8EB1",
			x"0000" when x"8EB2",
			x"0000" when x"8EB3",
			x"0000" when x"8EB4",
			x"0000" when x"8EB5",
			x"0000" when x"8EB6",
			x"0000" when x"8EB7",
			x"0000" when x"8EB8",
			x"0000" when x"8EB9",
			x"0000" when x"8EBA",
			x"0000" when x"8EBB",
			x"0000" when x"8EBC",
			x"0000" when x"8EBD",
			x"0000" when x"8EBE",
			x"0000" when x"8EBF",
			x"0000" when x"8EC0",
			x"0000" when x"8EC1",
			x"0000" when x"8EC2",
			x"0000" when x"8EC3",
			x"0000" when x"8EC4",
			x"0000" when x"8EC5",
			x"0000" when x"8EC6",
			x"0000" when x"8EC7",
			x"0000" when x"8EC8",
			x"0000" when x"8EC9",
			x"0000" when x"8ECA",
			x"0000" when x"8ECB",
			x"0000" when x"8ECC",
			x"0000" when x"8ECD",
			x"0000" when x"8ECE",
			x"0000" when x"8ECF",
			x"0000" when x"8ED0",
			x"0000" when x"8ED1",
			x"0000" when x"8ED2",
			x"0000" when x"8ED3",
			x"0000" when x"8ED4",
			x"0000" when x"8ED5",
			x"0000" when x"8ED6",
			x"0000" when x"8ED7",
			x"0000" when x"8ED8",
			x"0000" when x"8ED9",
			x"0000" when x"8EDA",
			x"0000" when x"8EDB",
			x"0000" when x"8EDC",
			x"0000" when x"8EDD",
			x"0000" when x"8EDE",
			x"0000" when x"8EDF",
			x"0000" when x"8EE0",
			x"0000" when x"8EE1",
			x"0000" when x"8EE2",
			x"0000" when x"8EE3",
			x"0000" when x"8EE4",
			x"0000" when x"8EE5",
			x"0000" when x"8EE6",
			x"0000" when x"8EE7",
			x"0000" when x"8EE8",
			x"0000" when x"8EE9",
			x"0000" when x"8EEA",
			x"0000" when x"8EEB",
			x"0000" when x"8EEC",
			x"0000" when x"8EED",
			x"0000" when x"8EEE",
			x"0000" when x"8EEF",
			x"0000" when x"8EF0",
			x"0000" when x"8EF1",
			x"0000" when x"8EF2",
			x"0000" when x"8EF3",
			x"0000" when x"8EF4",
			x"0000" when x"8EF5",
			x"0000" when x"8EF6",
			x"0000" when x"8EF7",
			x"0000" when x"8EF8",
			x"0000" when x"8EF9",
			x"0000" when x"8EFA",
			x"0000" when x"8EFB",
			x"0000" when x"8EFC",
			x"0000" when x"8EFD",
			x"0000" when x"8EFE",
			x"0000" when x"8EFF",
			x"0000" when x"8F00",
			x"0000" when x"8F01",
			x"0000" when x"8F02",
			x"0000" when x"8F03",
			x"0000" when x"8F04",
			x"0000" when x"8F05",
			x"0000" when x"8F06",
			x"0000" when x"8F07",
			x"0000" when x"8F08",
			x"0000" when x"8F09",
			x"0000" when x"8F0A",
			x"0000" when x"8F0B",
			x"0000" when x"8F0C",
			x"0000" when x"8F0D",
			x"0000" when x"8F0E",
			x"0000" when x"8F0F",
			x"0000" when x"8F10",
			x"0000" when x"8F11",
			x"0000" when x"8F12",
			x"0000" when x"8F13",
			x"0000" when x"8F14",
			x"0000" when x"8F15",
			x"0000" when x"8F16",
			x"0000" when x"8F17",
			x"0000" when x"8F18",
			x"0000" when x"8F19",
			x"0000" when x"8F1A",
			x"0000" when x"8F1B",
			x"0000" when x"8F1C",
			x"0000" when x"8F1D",
			x"0000" when x"8F1E",
			x"0000" when x"8F1F",
			x"0000" when x"8F20",
			x"0000" when x"8F21",
			x"0000" when x"8F22",
			x"0000" when x"8F23",
			x"0000" when x"8F24",
			x"0000" when x"8F25",
			x"0000" when x"8F26",
			x"0000" when x"8F27",
			x"0000" when x"8F28",
			x"0000" when x"8F29",
			x"0000" when x"8F2A",
			x"0000" when x"8F2B",
			x"0000" when x"8F2C",
			x"0000" when x"8F2D",
			x"0000" when x"8F2E",
			x"0000" when x"8F2F",
			x"0000" when x"8F30",
			x"0000" when x"8F31",
			x"0000" when x"8F32",
			x"0000" when x"8F33",
			x"0000" when x"8F34",
			x"0000" when x"8F35",
			x"0000" when x"8F36",
			x"0000" when x"8F37",
			x"0000" when x"8F38",
			x"0000" when x"8F39",
			x"0000" when x"8F3A",
			x"0000" when x"8F3B",
			x"0000" when x"8F3C",
			x"0000" when x"8F3D",
			x"0000" when x"8F3E",
			x"0000" when x"8F3F",
			x"0000" when x"8F40",
			x"0000" when x"8F41",
			x"0000" when x"8F42",
			x"0000" when x"8F43",
			x"0000" when x"8F44",
			x"0000" when x"8F45",
			x"0000" when x"8F46",
			x"0000" when x"8F47",
			x"0000" when x"8F48",
			x"0000" when x"8F49",
			x"0000" when x"8F4A",
			x"0000" when x"8F4B",
			x"0000" when x"8F4C",
			x"0000" when x"8F4D",
			x"0000" when x"8F4E",
			x"0000" when x"8F4F",
			x"0000" when x"8F50",
			x"0000" when x"8F51",
			x"0000" when x"8F52",
			x"0000" when x"8F53",
			x"0000" when x"8F54",
			x"0000" when x"8F55",
			x"0000" when x"8F56",
			x"0000" when x"8F57",
			x"0000" when x"8F58",
			x"0000" when x"8F59",
			x"0000" when x"8F5A",
			x"0000" when x"8F5B",
			x"0000" when x"8F5C",
			x"0000" when x"8F5D",
			x"0000" when x"8F5E",
			x"0000" when x"8F5F",
			x"0000" when x"8F60",
			x"0000" when x"8F61",
			x"0000" when x"8F62",
			x"0000" when x"8F63",
			x"0000" when x"8F64",
			x"0000" when x"8F65",
			x"0000" when x"8F66",
			x"0000" when x"8F67",
			x"0000" when x"8F68",
			x"0000" when x"8F69",
			x"0000" when x"8F6A",
			x"0000" when x"8F6B",
			x"0000" when x"8F6C",
			x"0000" when x"8F6D",
			x"0000" when x"8F6E",
			x"0000" when x"8F6F",
			x"0000" when x"8F70",
			x"0000" when x"8F71",
			x"0000" when x"8F72",
			x"0000" when x"8F73",
			x"0000" when x"8F74",
			x"0000" when x"8F75",
			x"0000" when x"8F76",
			x"0000" when x"8F77",
			x"0000" when x"8F78",
			x"0000" when x"8F79",
			x"0000" when x"8F7A",
			x"0000" when x"8F7B",
			x"0000" when x"8F7C",
			x"0000" when x"8F7D",
			x"0000" when x"8F7E",
			x"0000" when x"8F7F",
			x"0000" when x"8F80",
			x"0000" when x"8F81",
			x"0000" when x"8F82",
			x"0000" when x"8F83",
			x"0000" when x"8F84",
			x"0000" when x"8F85",
			x"0000" when x"8F86",
			x"0000" when x"8F87",
			x"0000" when x"8F88",
			x"0000" when x"8F89",
			x"0000" when x"8F8A",
			x"0000" when x"8F8B",
			x"0000" when x"8F8C",
			x"0000" when x"8F8D",
			x"0000" when x"8F8E",
			x"0000" when x"8F8F",
			x"0000" when x"8F90",
			x"0000" when x"8F91",
			x"0000" when x"8F92",
			x"0000" when x"8F93",
			x"0000" when x"8F94",
			x"0000" when x"8F95",
			x"0000" when x"8F96",
			x"0000" when x"8F97",
			x"0000" when x"8F98",
			x"0000" when x"8F99",
			x"0000" when x"8F9A",
			x"0000" when x"8F9B",
			x"0000" when x"8F9C",
			x"0000" when x"8F9D",
			x"0000" when x"8F9E",
			x"0000" when x"8F9F",
			x"0000" when x"8FA0",
			x"0000" when x"8FA1",
			x"0000" when x"8FA2",
			x"0000" when x"8FA3",
			x"0000" when x"8FA4",
			x"0000" when x"8FA5",
			x"0000" when x"8FA6",
			x"0000" when x"8FA7",
			x"0000" when x"8FA8",
			x"0000" when x"8FA9",
			x"0000" when x"8FAA",
			x"0000" when x"8FAB",
			x"0000" when x"8FAC",
			x"0000" when x"8FAD",
			x"0000" when x"8FAE",
			x"0000" when x"8FAF",
			x"0000" when x"8FB0",
			x"0000" when x"8FB1",
			x"0000" when x"8FB2",
			x"0000" when x"8FB3",
			x"0000" when x"8FB4",
			x"0000" when x"8FB5",
			x"0000" when x"8FB6",
			x"0000" when x"8FB7",
			x"0000" when x"8FB8",
			x"0000" when x"8FB9",
			x"0000" when x"8FBA",
			x"0000" when x"8FBB",
			x"0000" when x"8FBC",
			x"0000" when x"8FBD",
			x"0000" when x"8FBE",
			x"0000" when x"8FBF",
			x"0000" when x"8FC0",
			x"0000" when x"8FC1",
			x"0000" when x"8FC2",
			x"0000" when x"8FC3",
			x"0000" when x"8FC4",
			x"0000" when x"8FC5",
			x"0000" when x"8FC6",
			x"0000" when x"8FC7",
			x"0000" when x"8FC8",
			x"0000" when x"8FC9",
			x"0000" when x"8FCA",
			x"0000" when x"8FCB",
			x"0000" when x"8FCC",
			x"0000" when x"8FCD",
			x"0000" when x"8FCE",
			x"0000" when x"8FCF",
			x"0000" when x"8FD0",
			x"0000" when x"8FD1",
			x"0000" when x"8FD2",
			x"0000" when x"8FD3",
			x"0000" when x"8FD4",
			x"0000" when x"8FD5",
			x"0000" when x"8FD6",
			x"0000" when x"8FD7",
			x"0000" when x"8FD8",
			x"0000" when x"8FD9",
			x"0000" when x"8FDA",
			x"0000" when x"8FDB",
			x"0000" when x"8FDC",
			x"0000" when x"8FDD",
			x"0000" when x"8FDE",
			x"0000" when x"8FDF",
			x"0000" when x"8FE0",
			x"0000" when x"8FE1",
			x"0000" when x"8FE2",
			x"0000" when x"8FE3",
			x"0000" when x"8FE4",
			x"0000" when x"8FE5",
			x"0000" when x"8FE6",
			x"0000" when x"8FE7",
			x"0000" when x"8FE8",
			x"0000" when x"8FE9",
			x"0000" when x"8FEA",
			x"0000" when x"8FEB",
			x"0000" when x"8FEC",
			x"0000" when x"8FED",
			x"0000" when x"8FEE",
			x"0000" when x"8FEF",
			x"0000" when x"8FF0",
			x"0000" when x"8FF1",
			x"0000" when x"8FF2",
			x"0000" when x"8FF3",
			x"0000" when x"8FF4",
			x"0000" when x"8FF5",
			x"0000" when x"8FF6",
			x"0000" when x"8FF7",
			x"0000" when x"8FF8",
			x"0000" when x"8FF9",
			x"0000" when x"8FFA",
			x"0000" when x"8FFB",
			x"0000" when x"8FFC",
			x"0000" when x"8FFD",
			x"0000" when x"8FFE",
			x"0000" when x"8FFF",
			x"0000" when x"9000",
			x"0000" when x"9001",
			x"0000" when x"9002",
			x"0000" when x"9003",
			x"0000" when x"9004",
			x"0000" when x"9005",
			x"0000" when x"9006",
			x"0000" when x"9007",
			x"0000" when x"9008",
			x"0000" when x"9009",
			x"0000" when x"900A",
			x"0000" when x"900B",
			x"0000" when x"900C",
			x"0000" when x"900D",
			x"0000" when x"900E",
			x"0000" when x"900F",
			x"0000" when x"9010",
			x"0000" when x"9011",
			x"0000" when x"9012",
			x"0000" when x"9013",
			x"0000" when x"9014",
			x"0000" when x"9015",
			x"0000" when x"9016",
			x"0000" when x"9017",
			x"0000" when x"9018",
			x"0000" when x"9019",
			x"0000" when x"901A",
			x"0000" when x"901B",
			x"0000" when x"901C",
			x"0000" when x"901D",
			x"0000" when x"901E",
			x"0000" when x"901F",
			x"0000" when x"9020",
			x"0000" when x"9021",
			x"0000" when x"9022",
			x"0000" when x"9023",
			x"0000" when x"9024",
			x"0000" when x"9025",
			x"0000" when x"9026",
			x"0000" when x"9027",
			x"0000" when x"9028",
			x"0000" when x"9029",
			x"0000" when x"902A",
			x"0000" when x"902B",
			x"0000" when x"902C",
			x"0000" when x"902D",
			x"0000" when x"902E",
			x"0000" when x"902F",
			x"0000" when x"9030",
			x"0000" when x"9031",
			x"0000" when x"9032",
			x"0000" when x"9033",
			x"0000" when x"9034",
			x"0000" when x"9035",
			x"0000" when x"9036",
			x"0000" when x"9037",
			x"0000" when x"9038",
			x"0000" when x"9039",
			x"0000" when x"903A",
			x"0000" when x"903B",
			x"0000" when x"903C",
			x"0000" when x"903D",
			x"0000" when x"903E",
			x"0000" when x"903F",
			x"0000" when x"9040",
			x"0000" when x"9041",
			x"0000" when x"9042",
			x"0000" when x"9043",
			x"0000" when x"9044",
			x"0000" when x"9045",
			x"0000" when x"9046",
			x"0000" when x"9047",
			x"0000" when x"9048",
			x"0000" when x"9049",
			x"0000" when x"904A",
			x"0000" when x"904B",
			x"0000" when x"904C",
			x"0000" when x"904D",
			x"0000" when x"904E",
			x"0000" when x"904F",
			x"0000" when x"9050",
			x"0000" when x"9051",
			x"0000" when x"9052",
			x"0000" when x"9053",
			x"0000" when x"9054",
			x"0000" when x"9055",
			x"0000" when x"9056",
			x"0000" when x"9057",
			x"0000" when x"9058",
			x"0000" when x"9059",
			x"0000" when x"905A",
			x"0000" when x"905B",
			x"0000" when x"905C",
			x"0000" when x"905D",
			x"0000" when x"905E",
			x"0000" when x"905F",
			x"0000" when x"9060",
			x"0000" when x"9061",
			x"0000" when x"9062",
			x"0000" when x"9063",
			x"0000" when x"9064",
			x"0000" when x"9065",
			x"0000" when x"9066",
			x"0000" when x"9067",
			x"0000" when x"9068",
			x"0000" when x"9069",
			x"0000" when x"906A",
			x"0000" when x"906B",
			x"0000" when x"906C",
			x"0000" when x"906D",
			x"0000" when x"906E",
			x"0000" when x"906F",
			x"0000" when x"9070",
			x"0000" when x"9071",
			x"0000" when x"9072",
			x"0000" when x"9073",
			x"0000" when x"9074",
			x"0000" when x"9075",
			x"0000" when x"9076",
			x"0000" when x"9077",
			x"0000" when x"9078",
			x"0000" when x"9079",
			x"0000" when x"907A",
			x"0000" when x"907B",
			x"0000" when x"907C",
			x"0000" when x"907D",
			x"0000" when x"907E",
			x"0000" when x"907F",
			x"0000" when x"9080",
			x"0000" when x"9081",
			x"0000" when x"9082",
			x"0000" when x"9083",
			x"0000" when x"9084",
			x"0000" when x"9085",
			x"0000" when x"9086",
			x"0000" when x"9087",
			x"0000" when x"9088",
			x"0000" when x"9089",
			x"0000" when x"908A",
			x"0000" when x"908B",
			x"0000" when x"908C",
			x"0000" when x"908D",
			x"0000" when x"908E",
			x"0000" when x"908F",
			x"0000" when x"9090",
			x"0000" when x"9091",
			x"0000" when x"9092",
			x"0000" when x"9093",
			x"0000" when x"9094",
			x"0000" when x"9095",
			x"0000" when x"9096",
			x"0000" when x"9097",
			x"0000" when x"9098",
			x"0000" when x"9099",
			x"0000" when x"909A",
			x"0000" when x"909B",
			x"0000" when x"909C",
			x"0000" when x"909D",
			x"0000" when x"909E",
			x"0000" when x"909F",
			x"0000" when x"90A0",
			x"0000" when x"90A1",
			x"0000" when x"90A2",
			x"0000" when x"90A3",
			x"0000" when x"90A4",
			x"0000" when x"90A5",
			x"0000" when x"90A6",
			x"0000" when x"90A7",
			x"0000" when x"90A8",
			x"0000" when x"90A9",
			x"0000" when x"90AA",
			x"0000" when x"90AB",
			x"0000" when x"90AC",
			x"0000" when x"90AD",
			x"0000" when x"90AE",
			x"0000" when x"90AF",
			x"0000" when x"90B0",
			x"0000" when x"90B1",
			x"0000" when x"90B2",
			x"0000" when x"90B3",
			x"0000" when x"90B4",
			x"0000" when x"90B5",
			x"0000" when x"90B6",
			x"0000" when x"90B7",
			x"0000" when x"90B8",
			x"0000" when x"90B9",
			x"0000" when x"90BA",
			x"0000" when x"90BB",
			x"0000" when x"90BC",
			x"0000" when x"90BD",
			x"0000" when x"90BE",
			x"0000" when x"90BF",
			x"0000" when x"90C0",
			x"0000" when x"90C1",
			x"0000" when x"90C2",
			x"0000" when x"90C3",
			x"0000" when x"90C4",
			x"0000" when x"90C5",
			x"0000" when x"90C6",
			x"0000" when x"90C7",
			x"0000" when x"90C8",
			x"0000" when x"90C9",
			x"0000" when x"90CA",
			x"0000" when x"90CB",
			x"0000" when x"90CC",
			x"0000" when x"90CD",
			x"0000" when x"90CE",
			x"0000" when x"90CF",
			x"0000" when x"90D0",
			x"0000" when x"90D1",
			x"0000" when x"90D2",
			x"0000" when x"90D3",
			x"0000" when x"90D4",
			x"0000" when x"90D5",
			x"0000" when x"90D6",
			x"0000" when x"90D7",
			x"0000" when x"90D8",
			x"0000" when x"90D9",
			x"0000" when x"90DA",
			x"0000" when x"90DB",
			x"0000" when x"90DC",
			x"0000" when x"90DD",
			x"0000" when x"90DE",
			x"0000" when x"90DF",
			x"0000" when x"90E0",
			x"0000" when x"90E1",
			x"0000" when x"90E2",
			x"0000" when x"90E3",
			x"0000" when x"90E4",
			x"0000" when x"90E5",
			x"0000" when x"90E6",
			x"0000" when x"90E7",
			x"0000" when x"90E8",
			x"0000" when x"90E9",
			x"0000" when x"90EA",
			x"0000" when x"90EB",
			x"0000" when x"90EC",
			x"0000" when x"90ED",
			x"0000" when x"90EE",
			x"0000" when x"90EF",
			x"0000" when x"90F0",
			x"0000" when x"90F1",
			x"0000" when x"90F2",
			x"0000" when x"90F3",
			x"0000" when x"90F4",
			x"0000" when x"90F5",
			x"0000" when x"90F6",
			x"0000" when x"90F7",
			x"0000" when x"90F8",
			x"0000" when x"90F9",
			x"0000" when x"90FA",
			x"0000" when x"90FB",
			x"0000" when x"90FC",
			x"0000" when x"90FD",
			x"0000" when x"90FE",
			x"0000" when x"90FF",
			x"0000" when x"9100",
			x"0000" when x"9101",
			x"0000" when x"9102",
			x"0000" when x"9103",
			x"0000" when x"9104",
			x"0000" when x"9105",
			x"0000" when x"9106",
			x"0000" when x"9107",
			x"0000" when x"9108",
			x"0000" when x"9109",
			x"0000" when x"910A",
			x"0000" when x"910B",
			x"0000" when x"910C",
			x"0000" when x"910D",
			x"0000" when x"910E",
			x"0000" when x"910F",
			x"0000" when x"9110",
			x"0000" when x"9111",
			x"0000" when x"9112",
			x"0000" when x"9113",
			x"0000" when x"9114",
			x"0000" when x"9115",
			x"0000" when x"9116",
			x"0000" when x"9117",
			x"0000" when x"9118",
			x"0000" when x"9119",
			x"0000" when x"911A",
			x"0000" when x"911B",
			x"0000" when x"911C",
			x"0000" when x"911D",
			x"0000" when x"911E",
			x"0000" when x"911F",
			x"0000" when x"9120",
			x"0000" when x"9121",
			x"0000" when x"9122",
			x"0000" when x"9123",
			x"0000" when x"9124",
			x"0000" when x"9125",
			x"0000" when x"9126",
			x"0000" when x"9127",
			x"0000" when x"9128",
			x"0000" when x"9129",
			x"0000" when x"912A",
			x"0000" when x"912B",
			x"0000" when x"912C",
			x"0000" when x"912D",
			x"0000" when x"912E",
			x"0000" when x"912F",
			x"0000" when x"9130",
			x"0000" when x"9131",
			x"0000" when x"9132",
			x"0000" when x"9133",
			x"0000" when x"9134",
			x"0000" when x"9135",
			x"0000" when x"9136",
			x"0000" when x"9137",
			x"0000" when x"9138",
			x"0000" when x"9139",
			x"0000" when x"913A",
			x"0000" when x"913B",
			x"0000" when x"913C",
			x"0000" when x"913D",
			x"0000" when x"913E",
			x"0000" when x"913F",
			x"0000" when x"9140",
			x"0000" when x"9141",
			x"0000" when x"9142",
			x"0000" when x"9143",
			x"0000" when x"9144",
			x"0000" when x"9145",
			x"0000" when x"9146",
			x"0000" when x"9147",
			x"0000" when x"9148",
			x"0000" when x"9149",
			x"0000" when x"914A",
			x"0000" when x"914B",
			x"0000" when x"914C",
			x"0000" when x"914D",
			x"0000" when x"914E",
			x"0000" when x"914F",
			x"0000" when x"9150",
			x"0000" when x"9151",
			x"0000" when x"9152",
			x"0000" when x"9153",
			x"0000" when x"9154",
			x"0000" when x"9155",
			x"0000" when x"9156",
			x"0000" when x"9157",
			x"0000" when x"9158",
			x"0000" when x"9159",
			x"0000" when x"915A",
			x"0000" when x"915B",
			x"0000" when x"915C",
			x"0000" when x"915D",
			x"0000" when x"915E",
			x"0000" when x"915F",
			x"0000" when x"9160",
			x"0000" when x"9161",
			x"0000" when x"9162",
			x"0000" when x"9163",
			x"0000" when x"9164",
			x"0000" when x"9165",
			x"0000" when x"9166",
			x"0000" when x"9167",
			x"0000" when x"9168",
			x"0000" when x"9169",
			x"0000" when x"916A",
			x"0000" when x"916B",
			x"0000" when x"916C",
			x"0000" when x"916D",
			x"0000" when x"916E",
			x"0000" when x"916F",
			x"0000" when x"9170",
			x"0000" when x"9171",
			x"0000" when x"9172",
			x"0000" when x"9173",
			x"0000" when x"9174",
			x"0000" when x"9175",
			x"0000" when x"9176",
			x"0000" when x"9177",
			x"0000" when x"9178",
			x"0000" when x"9179",
			x"0000" when x"917A",
			x"0000" when x"917B",
			x"0000" when x"917C",
			x"0000" when x"917D",
			x"0000" when x"917E",
			x"0000" when x"917F",
			x"0000" when x"9180",
			x"0000" when x"9181",
			x"0000" when x"9182",
			x"0000" when x"9183",
			x"0000" when x"9184",
			x"0000" when x"9185",
			x"0000" when x"9186",
			x"0000" when x"9187",
			x"0000" when x"9188",
			x"0000" when x"9189",
			x"0000" when x"918A",
			x"0000" when x"918B",
			x"0000" when x"918C",
			x"0000" when x"918D",
			x"0000" when x"918E",
			x"0000" when x"918F",
			x"0000" when x"9190",
			x"0000" when x"9191",
			x"0000" when x"9192",
			x"0000" when x"9193",
			x"0000" when x"9194",
			x"0000" when x"9195",
			x"0000" when x"9196",
			x"0000" when x"9197",
			x"0000" when x"9198",
			x"0000" when x"9199",
			x"0000" when x"919A",
			x"0000" when x"919B",
			x"0000" when x"919C",
			x"0000" when x"919D",
			x"0000" when x"919E",
			x"0000" when x"919F",
			x"0000" when x"91A0",
			x"0000" when x"91A1",
			x"0000" when x"91A2",
			x"0000" when x"91A3",
			x"0000" when x"91A4",
			x"0000" when x"91A5",
			x"0000" when x"91A6",
			x"0000" when x"91A7",
			x"0000" when x"91A8",
			x"0000" when x"91A9",
			x"0000" when x"91AA",
			x"0000" when x"91AB",
			x"0000" when x"91AC",
			x"0000" when x"91AD",
			x"0000" when x"91AE",
			x"0000" when x"91AF",
			x"0000" when x"91B0",
			x"0000" when x"91B1",
			x"0000" when x"91B2",
			x"0000" when x"91B3",
			x"0000" when x"91B4",
			x"0000" when x"91B5",
			x"0000" when x"91B6",
			x"0000" when x"91B7",
			x"0000" when x"91B8",
			x"0000" when x"91B9",
			x"0000" when x"91BA",
			x"0000" when x"91BB",
			x"0000" when x"91BC",
			x"0000" when x"91BD",
			x"0000" when x"91BE",
			x"0000" when x"91BF",
			x"0000" when x"91C0",
			x"0000" when x"91C1",
			x"0000" when x"91C2",
			x"0000" when x"91C3",
			x"0000" when x"91C4",
			x"0000" when x"91C5",
			x"0000" when x"91C6",
			x"0000" when x"91C7",
			x"0000" when x"91C8",
			x"0000" when x"91C9",
			x"0000" when x"91CA",
			x"0000" when x"91CB",
			x"0000" when x"91CC",
			x"0000" when x"91CD",
			x"0000" when x"91CE",
			x"0000" when x"91CF",
			x"0000" when x"91D0",
			x"0000" when x"91D1",
			x"0000" when x"91D2",
			x"0000" when x"91D3",
			x"0000" when x"91D4",
			x"0000" when x"91D5",
			x"0000" when x"91D6",
			x"0000" when x"91D7",
			x"0000" when x"91D8",
			x"0000" when x"91D9",
			x"0000" when x"91DA",
			x"0000" when x"91DB",
			x"0000" when x"91DC",
			x"0000" when x"91DD",
			x"0000" when x"91DE",
			x"0000" when x"91DF",
			x"0000" when x"91E0",
			x"0000" when x"91E1",
			x"0000" when x"91E2",
			x"0000" when x"91E3",
			x"0000" when x"91E4",
			x"0000" when x"91E5",
			x"0000" when x"91E6",
			x"0000" when x"91E7",
			x"0000" when x"91E8",
			x"0000" when x"91E9",
			x"0000" when x"91EA",
			x"0000" when x"91EB",
			x"0000" when x"91EC",
			x"0000" when x"91ED",
			x"0000" when x"91EE",
			x"0000" when x"91EF",
			x"0000" when x"91F0",
			x"0000" when x"91F1",
			x"0000" when x"91F2",
			x"0000" when x"91F3",
			x"0000" when x"91F4",
			x"0000" when x"91F5",
			x"0000" when x"91F6",
			x"0000" when x"91F7",
			x"0000" when x"91F8",
			x"0000" when x"91F9",
			x"0000" when x"91FA",
			x"0000" when x"91FB",
			x"0000" when x"91FC",
			x"0000" when x"91FD",
			x"0000" when x"91FE",
			x"0000" when x"91FF",
			x"0000" when x"9200",
			x"0000" when x"9201",
			x"0000" when x"9202",
			x"0000" when x"9203",
			x"0000" when x"9204",
			x"0000" when x"9205",
			x"0000" when x"9206",
			x"0000" when x"9207",
			x"0000" when x"9208",
			x"0000" when x"9209",
			x"0000" when x"920A",
			x"0000" when x"920B",
			x"0000" when x"920C",
			x"0000" when x"920D",
			x"0000" when x"920E",
			x"0000" when x"920F",
			x"0000" when x"9210",
			x"0000" when x"9211",
			x"0000" when x"9212",
			x"0000" when x"9213",
			x"0000" when x"9214",
			x"0000" when x"9215",
			x"0000" when x"9216",
			x"0000" when x"9217",
			x"0000" when x"9218",
			x"0000" when x"9219",
			x"0000" when x"921A",
			x"0000" when x"921B",
			x"0000" when x"921C",
			x"0000" when x"921D",
			x"0000" when x"921E",
			x"0000" when x"921F",
			x"0000" when x"9220",
			x"0000" when x"9221",
			x"0000" when x"9222",
			x"0000" when x"9223",
			x"0000" when x"9224",
			x"0000" when x"9225",
			x"0000" when x"9226",
			x"0000" when x"9227",
			x"0000" when x"9228",
			x"0000" when x"9229",
			x"0000" when x"922A",
			x"0000" when x"922B",
			x"0000" when x"922C",
			x"0000" when x"922D",
			x"0000" when x"922E",
			x"0000" when x"922F",
			x"0000" when x"9230",
			x"0000" when x"9231",
			x"0000" when x"9232",
			x"0000" when x"9233",
			x"0000" when x"9234",
			x"0000" when x"9235",
			x"0000" when x"9236",
			x"0000" when x"9237",
			x"0000" when x"9238",
			x"0000" when x"9239",
			x"0000" when x"923A",
			x"0000" when x"923B",
			x"0000" when x"923C",
			x"0000" when x"923D",
			x"0000" when x"923E",
			x"0000" when x"923F",
			x"0000" when x"9240",
			x"0000" when x"9241",
			x"0000" when x"9242",
			x"0000" when x"9243",
			x"0000" when x"9244",
			x"0000" when x"9245",
			x"0000" when x"9246",
			x"0000" when x"9247",
			x"0000" when x"9248",
			x"0000" when x"9249",
			x"0000" when x"924A",
			x"0000" when x"924B",
			x"0000" when x"924C",
			x"0000" when x"924D",
			x"0000" when x"924E",
			x"0000" when x"924F",
			x"0000" when x"9250",
			x"0000" when x"9251",
			x"0000" when x"9252",
			x"0000" when x"9253",
			x"0000" when x"9254",
			x"0000" when x"9255",
			x"0000" when x"9256",
			x"0000" when x"9257",
			x"0000" when x"9258",
			x"0000" when x"9259",
			x"0000" when x"925A",
			x"0000" when x"925B",
			x"0000" when x"925C",
			x"0000" when x"925D",
			x"0000" when x"925E",
			x"0000" when x"925F",
			x"0000" when x"9260",
			x"0000" when x"9261",
			x"0000" when x"9262",
			x"0000" when x"9263",
			x"0000" when x"9264",
			x"0000" when x"9265",
			x"0000" when x"9266",
			x"0000" when x"9267",
			x"0000" when x"9268",
			x"0000" when x"9269",
			x"0000" when x"926A",
			x"0000" when x"926B",
			x"0000" when x"926C",
			x"0000" when x"926D",
			x"0000" when x"926E",
			x"0000" when x"926F",
			x"0000" when x"9270",
			x"0000" when x"9271",
			x"0000" when x"9272",
			x"0000" when x"9273",
			x"0000" when x"9274",
			x"0000" when x"9275",
			x"0000" when x"9276",
			x"0000" when x"9277",
			x"0000" when x"9278",
			x"0000" when x"9279",
			x"0000" when x"927A",
			x"0000" when x"927B",
			x"0000" when x"927C",
			x"0000" when x"927D",
			x"0000" when x"927E",
			x"0000" when x"927F",
			x"0000" when x"9280",
			x"0000" when x"9281",
			x"0000" when x"9282",
			x"0000" when x"9283",
			x"0000" when x"9284",
			x"0000" when x"9285",
			x"0000" when x"9286",
			x"0000" when x"9287",
			x"0000" when x"9288",
			x"0000" when x"9289",
			x"0000" when x"928A",
			x"0000" when x"928B",
			x"0000" when x"928C",
			x"0000" when x"928D",
			x"0000" when x"928E",
			x"0000" when x"928F",
			x"0000" when x"9290",
			x"0000" when x"9291",
			x"0000" when x"9292",
			x"0000" when x"9293",
			x"0000" when x"9294",
			x"0000" when x"9295",
			x"0000" when x"9296",
			x"0000" when x"9297",
			x"0000" when x"9298",
			x"0000" when x"9299",
			x"0000" when x"929A",
			x"0000" when x"929B",
			x"0000" when x"929C",
			x"0000" when x"929D",
			x"0000" when x"929E",
			x"0000" when x"929F",
			x"0000" when x"92A0",
			x"0000" when x"92A1",
			x"0000" when x"92A2",
			x"0000" when x"92A3",
			x"0000" when x"92A4",
			x"0000" when x"92A5",
			x"0000" when x"92A6",
			x"0000" when x"92A7",
			x"0000" when x"92A8",
			x"0000" when x"92A9",
			x"0000" when x"92AA",
			x"0000" when x"92AB",
			x"0000" when x"92AC",
			x"0000" when x"92AD",
			x"0000" when x"92AE",
			x"0000" when x"92AF",
			x"0000" when x"92B0",
			x"0000" when x"92B1",
			x"0000" when x"92B2",
			x"0000" when x"92B3",
			x"0000" when x"92B4",
			x"0000" when x"92B5",
			x"0000" when x"92B6",
			x"0000" when x"92B7",
			x"0000" when x"92B8",
			x"0000" when x"92B9",
			x"0000" when x"92BA",
			x"0000" when x"92BB",
			x"0000" when x"92BC",
			x"0000" when x"92BD",
			x"0000" when x"92BE",
			x"0000" when x"92BF",
			x"0000" when x"92C0",
			x"0000" when x"92C1",
			x"0000" when x"92C2",
			x"0000" when x"92C3",
			x"0000" when x"92C4",
			x"0000" when x"92C5",
			x"0000" when x"92C6",
			x"0000" when x"92C7",
			x"0000" when x"92C8",
			x"0000" when x"92C9",
			x"0000" when x"92CA",
			x"0000" when x"92CB",
			x"0000" when x"92CC",
			x"0000" when x"92CD",
			x"0000" when x"92CE",
			x"0000" when x"92CF",
			x"0000" when x"92D0",
			x"0000" when x"92D1",
			x"0000" when x"92D2",
			x"0000" when x"92D3",
			x"0000" when x"92D4",
			x"0000" when x"92D5",
			x"0000" when x"92D6",
			x"0000" when x"92D7",
			x"0000" when x"92D8",
			x"0000" when x"92D9",
			x"0000" when x"92DA",
			x"0000" when x"92DB",
			x"0000" when x"92DC",
			x"0000" when x"92DD",
			x"0000" when x"92DE",
			x"0000" when x"92DF",
			x"0000" when x"92E0",
			x"0000" when x"92E1",
			x"0000" when x"92E2",
			x"0000" when x"92E3",
			x"0000" when x"92E4",
			x"0000" when x"92E5",
			x"0000" when x"92E6",
			x"0000" when x"92E7",
			x"0000" when x"92E8",
			x"0000" when x"92E9",
			x"0000" when x"92EA",
			x"0000" when x"92EB",
			x"0000" when x"92EC",
			x"0000" when x"92ED",
			x"0000" when x"92EE",
			x"0000" when x"92EF",
			x"0000" when x"92F0",
			x"0000" when x"92F1",
			x"0000" when x"92F2",
			x"0000" when x"92F3",
			x"0000" when x"92F4",
			x"0000" when x"92F5",
			x"0000" when x"92F6",
			x"0000" when x"92F7",
			x"0000" when x"92F8",
			x"0000" when x"92F9",
			x"0000" when x"92FA",
			x"0000" when x"92FB",
			x"0000" when x"92FC",
			x"0000" when x"92FD",
			x"0000" when x"92FE",
			x"0000" when x"92FF",
			x"0000" when x"9300",
			x"0000" when x"9301",
			x"0000" when x"9302",
			x"0000" when x"9303",
			x"0000" when x"9304",
			x"0000" when x"9305",
			x"0000" when x"9306",
			x"0000" when x"9307",
			x"0000" when x"9308",
			x"0000" when x"9309",
			x"0000" when x"930A",
			x"0000" when x"930B",
			x"0000" when x"930C",
			x"0000" when x"930D",
			x"0000" when x"930E",
			x"0000" when x"930F",
			x"0000" when x"9310",
			x"0000" when x"9311",
			x"0000" when x"9312",
			x"0000" when x"9313",
			x"0000" when x"9314",
			x"0000" when x"9315",
			x"0000" when x"9316",
			x"0000" when x"9317",
			x"0000" when x"9318",
			x"0000" when x"9319",
			x"0000" when x"931A",
			x"0000" when x"931B",
			x"0000" when x"931C",
			x"0000" when x"931D",
			x"0000" when x"931E",
			x"0000" when x"931F",
			x"0000" when x"9320",
			x"0000" when x"9321",
			x"0000" when x"9322",
			x"0000" when x"9323",
			x"0000" when x"9324",
			x"0000" when x"9325",
			x"0000" when x"9326",
			x"0000" when x"9327",
			x"0000" when x"9328",
			x"0000" when x"9329",
			x"0000" when x"932A",
			x"0000" when x"932B",
			x"0000" when x"932C",
			x"0000" when x"932D",
			x"0000" when x"932E",
			x"0000" when x"932F",
			x"0000" when x"9330",
			x"0000" when x"9331",
			x"0000" when x"9332",
			x"0000" when x"9333",
			x"0000" when x"9334",
			x"0000" when x"9335",
			x"0000" when x"9336",
			x"0000" when x"9337",
			x"0000" when x"9338",
			x"0000" when x"9339",
			x"0000" when x"933A",
			x"0000" when x"933B",
			x"0000" when x"933C",
			x"0000" when x"933D",
			x"0000" when x"933E",
			x"0000" when x"933F",
			x"0000" when x"9340",
			x"0000" when x"9341",
			x"0000" when x"9342",
			x"0000" when x"9343",
			x"0000" when x"9344",
			x"0000" when x"9345",
			x"0000" when x"9346",
			x"0000" when x"9347",
			x"0000" when x"9348",
			x"0000" when x"9349",
			x"0000" when x"934A",
			x"0000" when x"934B",
			x"0000" when x"934C",
			x"0000" when x"934D",
			x"0000" when x"934E",
			x"0000" when x"934F",
			x"0000" when x"9350",
			x"0000" when x"9351",
			x"0000" when x"9352",
			x"0000" when x"9353",
			x"0000" when x"9354",
			x"0000" when x"9355",
			x"0000" when x"9356",
			x"0000" when x"9357",
			x"0000" when x"9358",
			x"0000" when x"9359",
			x"0000" when x"935A",
			x"0000" when x"935B",
			x"0000" when x"935C",
			x"0000" when x"935D",
			x"0000" when x"935E",
			x"0000" when x"935F",
			x"0000" when x"9360",
			x"0000" when x"9361",
			x"0000" when x"9362",
			x"0000" when x"9363",
			x"0000" when x"9364",
			x"0000" when x"9365",
			x"0000" when x"9366",
			x"0000" when x"9367",
			x"0000" when x"9368",
			x"0000" when x"9369",
			x"0000" when x"936A",
			x"0000" when x"936B",
			x"0000" when x"936C",
			x"0000" when x"936D",
			x"0000" when x"936E",
			x"0000" when x"936F",
			x"0000" when x"9370",
			x"0000" when x"9371",
			x"0000" when x"9372",
			x"0000" when x"9373",
			x"0000" when x"9374",
			x"0000" when x"9375",
			x"0000" when x"9376",
			x"0000" when x"9377",
			x"0000" when x"9378",
			x"0000" when x"9379",
			x"0000" when x"937A",
			x"0000" when x"937B",
			x"0000" when x"937C",
			x"0000" when x"937D",
			x"0000" when x"937E",
			x"0000" when x"937F",
			x"0000" when x"9380",
			x"0000" when x"9381",
			x"0000" when x"9382",
			x"0000" when x"9383",
			x"0000" when x"9384",
			x"0000" when x"9385",
			x"0000" when x"9386",
			x"0000" when x"9387",
			x"0000" when x"9388",
			x"0000" when x"9389",
			x"0000" when x"938A",
			x"0000" when x"938B",
			x"0000" when x"938C",
			x"0000" when x"938D",
			x"0000" when x"938E",
			x"0000" when x"938F",
			x"0000" when x"9390",
			x"0000" when x"9391",
			x"0000" when x"9392",
			x"0000" when x"9393",
			x"0000" when x"9394",
			x"0000" when x"9395",
			x"0000" when x"9396",
			x"0000" when x"9397",
			x"0000" when x"9398",
			x"0000" when x"9399",
			x"0000" when x"939A",
			x"0000" when x"939B",
			x"0000" when x"939C",
			x"0000" when x"939D",
			x"0000" when x"939E",
			x"0000" when x"939F",
			x"0000" when x"93A0",
			x"0000" when x"93A1",
			x"0000" when x"93A2",
			x"0000" when x"93A3",
			x"0000" when x"93A4",
			x"0000" when x"93A5",
			x"0000" when x"93A6",
			x"0000" when x"93A7",
			x"0000" when x"93A8",
			x"0000" when x"93A9",
			x"0000" when x"93AA",
			x"0000" when x"93AB",
			x"0000" when x"93AC",
			x"0000" when x"93AD",
			x"0000" when x"93AE",
			x"0000" when x"93AF",
			x"0000" when x"93B0",
			x"0000" when x"93B1",
			x"0000" when x"93B2",
			x"0000" when x"93B3",
			x"0000" when x"93B4",
			x"0000" when x"93B5",
			x"0000" when x"93B6",
			x"0000" when x"93B7",
			x"0000" when x"93B8",
			x"0000" when x"93B9",
			x"0000" when x"93BA",
			x"0000" when x"93BB",
			x"0000" when x"93BC",
			x"0000" when x"93BD",
			x"0000" when x"93BE",
			x"0000" when x"93BF",
			x"0000" when x"93C0",
			x"0000" when x"93C1",
			x"0000" when x"93C2",
			x"0000" when x"93C3",
			x"0000" when x"93C4",
			x"0000" when x"93C5",
			x"0000" when x"93C6",
			x"0000" when x"93C7",
			x"0000" when x"93C8",
			x"0000" when x"93C9",
			x"0000" when x"93CA",
			x"0000" when x"93CB",
			x"0000" when x"93CC",
			x"0000" when x"93CD",
			x"0000" when x"93CE",
			x"0000" when x"93CF",
			x"0000" when x"93D0",
			x"0000" when x"93D1",
			x"0000" when x"93D2",
			x"0000" when x"93D3",
			x"0000" when x"93D4",
			x"0000" when x"93D5",
			x"0000" when x"93D6",
			x"0000" when x"93D7",
			x"0000" when x"93D8",
			x"0000" when x"93D9",
			x"0000" when x"93DA",
			x"0000" when x"93DB",
			x"0000" when x"93DC",
			x"0000" when x"93DD",
			x"0000" when x"93DE",
			x"0000" when x"93DF",
			x"0000" when x"93E0",
			x"0000" when x"93E1",
			x"0000" when x"93E2",
			x"0000" when x"93E3",
			x"0000" when x"93E4",
			x"0000" when x"93E5",
			x"0000" when x"93E6",
			x"0000" when x"93E7",
			x"0000" when x"93E8",
			x"0000" when x"93E9",
			x"0000" when x"93EA",
			x"0000" when x"93EB",
			x"0000" when x"93EC",
			x"0000" when x"93ED",
			x"0000" when x"93EE",
			x"0000" when x"93EF",
			x"0000" when x"93F0",
			x"0000" when x"93F1",
			x"0000" when x"93F2",
			x"0000" when x"93F3",
			x"0000" when x"93F4",
			x"0000" when x"93F5",
			x"0000" when x"93F6",
			x"0000" when x"93F7",
			x"0000" when x"93F8",
			x"0000" when x"93F9",
			x"0000" when x"93FA",
			x"0000" when x"93FB",
			x"0000" when x"93FC",
			x"0000" when x"93FD",
			x"0000" when x"93FE",
			x"0000" when x"93FF",
			x"0000" when x"9400",
			x"0000" when x"9401",
			x"0000" when x"9402",
			x"0000" when x"9403",
			x"0000" when x"9404",
			x"0000" when x"9405",
			x"0000" when x"9406",
			x"0000" when x"9407",
			x"0000" when x"9408",
			x"0000" when x"9409",
			x"0000" when x"940A",
			x"0000" when x"940B",
			x"0000" when x"940C",
			x"0000" when x"940D",
			x"0000" when x"940E",
			x"0000" when x"940F",
			x"0000" when x"9410",
			x"0000" when x"9411",
			x"0000" when x"9412",
			x"0000" when x"9413",
			x"0000" when x"9414",
			x"0000" when x"9415",
			x"0000" when x"9416",
			x"0000" when x"9417",
			x"0000" when x"9418",
			x"0000" when x"9419",
			x"0000" when x"941A",
			x"0000" when x"941B",
			x"0000" when x"941C",
			x"0000" when x"941D",
			x"0000" when x"941E",
			x"0000" when x"941F",
			x"0000" when x"9420",
			x"0000" when x"9421",
			x"0000" when x"9422",
			x"0000" when x"9423",
			x"0000" when x"9424",
			x"0000" when x"9425",
			x"0000" when x"9426",
			x"0000" when x"9427",
			x"0000" when x"9428",
			x"0000" when x"9429",
			x"0000" when x"942A",
			x"0000" when x"942B",
			x"0000" when x"942C",
			x"0000" when x"942D",
			x"0000" when x"942E",
			x"0000" when x"942F",
			x"0000" when x"9430",
			x"0000" when x"9431",
			x"0000" when x"9432",
			x"0000" when x"9433",
			x"0000" when x"9434",
			x"0000" when x"9435",
			x"0000" when x"9436",
			x"0000" when x"9437",
			x"0000" when x"9438",
			x"0000" when x"9439",
			x"0000" when x"943A",
			x"0000" when x"943B",
			x"0000" when x"943C",
			x"0000" when x"943D",
			x"0000" when x"943E",
			x"0000" when x"943F",
			x"0000" when x"9440",
			x"0000" when x"9441",
			x"0000" when x"9442",
			x"0000" when x"9443",
			x"0000" when x"9444",
			x"0000" when x"9445",
			x"0000" when x"9446",
			x"0000" when x"9447",
			x"0000" when x"9448",
			x"0000" when x"9449",
			x"0000" when x"944A",
			x"0000" when x"944B",
			x"0000" when x"944C",
			x"0000" when x"944D",
			x"0000" when x"944E",
			x"0000" when x"944F",
			x"0000" when x"9450",
			x"0000" when x"9451",
			x"0000" when x"9452",
			x"0000" when x"9453",
			x"0000" when x"9454",
			x"0000" when x"9455",
			x"0000" when x"9456",
			x"0000" when x"9457",
			x"0000" when x"9458",
			x"0000" when x"9459",
			x"0000" when x"945A",
			x"0000" when x"945B",
			x"0000" when x"945C",
			x"0000" when x"945D",
			x"0000" when x"945E",
			x"0000" when x"945F",
			x"0000" when x"9460",
			x"0000" when x"9461",
			x"0000" when x"9462",
			x"0000" when x"9463",
			x"0000" when x"9464",
			x"0000" when x"9465",
			x"0000" when x"9466",
			x"0000" when x"9467",
			x"0000" when x"9468",
			x"0000" when x"9469",
			x"0000" when x"946A",
			x"0000" when x"946B",
			x"0000" when x"946C",
			x"0000" when x"946D",
			x"0000" when x"946E",
			x"0000" when x"946F",
			x"0000" when x"9470",
			x"0000" when x"9471",
			x"0000" when x"9472",
			x"0000" when x"9473",
			x"0000" when x"9474",
			x"0000" when x"9475",
			x"0000" when x"9476",
			x"0000" when x"9477",
			x"0000" when x"9478",
			x"0000" when x"9479",
			x"0000" when x"947A",
			x"0000" when x"947B",
			x"0000" when x"947C",
			x"0000" when x"947D",
			x"0000" when x"947E",
			x"0000" when x"947F",
			x"0000" when x"9480",
			x"0000" when x"9481",
			x"0000" when x"9482",
			x"0000" when x"9483",
			x"0000" when x"9484",
			x"0000" when x"9485",
			x"0000" when x"9486",
			x"0000" when x"9487",
			x"0000" when x"9488",
			x"0000" when x"9489",
			x"0000" when x"948A",
			x"0000" when x"948B",
			x"0000" when x"948C",
			x"0000" when x"948D",
			x"0000" when x"948E",
			x"0000" when x"948F",
			x"0000" when x"9490",
			x"0000" when x"9491",
			x"0000" when x"9492",
			x"0000" when x"9493",
			x"0000" when x"9494",
			x"0000" when x"9495",
			x"0000" when x"9496",
			x"0000" when x"9497",
			x"0000" when x"9498",
			x"0000" when x"9499",
			x"0000" when x"949A",
			x"0000" when x"949B",
			x"0000" when x"949C",
			x"0000" when x"949D",
			x"0000" when x"949E",
			x"0000" when x"949F",
			x"0000" when x"94A0",
			x"0000" when x"94A1",
			x"0000" when x"94A2",
			x"0000" when x"94A3",
			x"0000" when x"94A4",
			x"0000" when x"94A5",
			x"0000" when x"94A6",
			x"0000" when x"94A7",
			x"0000" when x"94A8",
			x"0000" when x"94A9",
			x"0000" when x"94AA",
			x"0000" when x"94AB",
			x"0000" when x"94AC",
			x"0000" when x"94AD",
			x"0000" when x"94AE",
			x"0000" when x"94AF",
			x"0000" when x"94B0",
			x"0000" when x"94B1",
			x"0000" when x"94B2",
			x"0000" when x"94B3",
			x"0000" when x"94B4",
			x"0000" when x"94B5",
			x"0000" when x"94B6",
			x"0000" when x"94B7",
			x"0000" when x"94B8",
			x"0000" when x"94B9",
			x"0000" when x"94BA",
			x"0000" when x"94BB",
			x"0000" when x"94BC",
			x"0000" when x"94BD",
			x"0000" when x"94BE",
			x"0000" when x"94BF",
			x"0000" when x"94C0",
			x"0000" when x"94C1",
			x"0000" when x"94C2",
			x"0000" when x"94C3",
			x"0000" when x"94C4",
			x"0000" when x"94C5",
			x"0000" when x"94C6",
			x"0000" when x"94C7",
			x"0000" when x"94C8",
			x"0000" when x"94C9",
			x"0000" when x"94CA",
			x"0000" when x"94CB",
			x"0000" when x"94CC",
			x"0000" when x"94CD",
			x"0000" when x"94CE",
			x"0000" when x"94CF",
			x"0000" when x"94D0",
			x"0000" when x"94D1",
			x"0000" when x"94D2",
			x"0000" when x"94D3",
			x"0000" when x"94D4",
			x"0000" when x"94D5",
			x"0000" when x"94D6",
			x"0000" when x"94D7",
			x"0000" when x"94D8",
			x"0000" when x"94D9",
			x"0000" when x"94DA",
			x"0000" when x"94DB",
			x"0000" when x"94DC",
			x"0000" when x"94DD",
			x"0000" when x"94DE",
			x"0000" when x"94DF",
			x"0000" when x"94E0",
			x"0000" when x"94E1",
			x"0000" when x"94E2",
			x"0000" when x"94E3",
			x"0000" when x"94E4",
			x"0000" when x"94E5",
			x"0000" when x"94E6",
			x"0000" when x"94E7",
			x"0000" when x"94E8",
			x"0000" when x"94E9",
			x"0000" when x"94EA",
			x"0000" when x"94EB",
			x"0000" when x"94EC",
			x"0000" when x"94ED",
			x"0000" when x"94EE",
			x"0000" when x"94EF",
			x"0000" when x"94F0",
			x"0000" when x"94F1",
			x"0000" when x"94F2",
			x"0000" when x"94F3",
			x"0000" when x"94F4",
			x"0000" when x"94F5",
			x"0000" when x"94F6",
			x"0000" when x"94F7",
			x"0000" when x"94F8",
			x"0000" when x"94F9",
			x"0000" when x"94FA",
			x"0000" when x"94FB",
			x"0000" when x"94FC",
			x"0000" when x"94FD",
			x"0000" when x"94FE",
			x"0000" when x"94FF",
			x"0000" when x"9500",
			x"0000" when x"9501",
			x"0000" when x"9502",
			x"0000" when x"9503",
			x"0000" when x"9504",
			x"0000" when x"9505",
			x"0000" when x"9506",
			x"0000" when x"9507",
			x"0000" when x"9508",
			x"0000" when x"9509",
			x"0000" when x"950A",
			x"0000" when x"950B",
			x"0000" when x"950C",
			x"0000" when x"950D",
			x"0000" when x"950E",
			x"0000" when x"950F",
			x"0000" when x"9510",
			x"0000" when x"9511",
			x"0000" when x"9512",
			x"0000" when x"9513",
			x"0000" when x"9514",
			x"0000" when x"9515",
			x"0000" when x"9516",
			x"0000" when x"9517",
			x"0000" when x"9518",
			x"0000" when x"9519",
			x"0000" when x"951A",
			x"0000" when x"951B",
			x"0000" when x"951C",
			x"0000" when x"951D",
			x"0000" when x"951E",
			x"0000" when x"951F",
			x"0000" when x"9520",
			x"0000" when x"9521",
			x"0000" when x"9522",
			x"0000" when x"9523",
			x"0000" when x"9524",
			x"0000" when x"9525",
			x"0000" when x"9526",
			x"0000" when x"9527",
			x"0000" when x"9528",
			x"0000" when x"9529",
			x"0000" when x"952A",
			x"0000" when x"952B",
			x"0000" when x"952C",
			x"0000" when x"952D",
			x"0000" when x"952E",
			x"0000" when x"952F",
			x"0000" when x"9530",
			x"0000" when x"9531",
			x"0000" when x"9532",
			x"0000" when x"9533",
			x"0000" when x"9534",
			x"0000" when x"9535",
			x"0000" when x"9536",
			x"0000" when x"9537",
			x"0000" when x"9538",
			x"0000" when x"9539",
			x"0000" when x"953A",
			x"0000" when x"953B",
			x"0000" when x"953C",
			x"0000" when x"953D",
			x"0000" when x"953E",
			x"0000" when x"953F",
			x"0000" when x"9540",
			x"0000" when x"9541",
			x"0000" when x"9542",
			x"0000" when x"9543",
			x"0000" when x"9544",
			x"0000" when x"9545",
			x"0000" when x"9546",
			x"0000" when x"9547",
			x"0000" when x"9548",
			x"0000" when x"9549",
			x"0000" when x"954A",
			x"0000" when x"954B",
			x"0000" when x"954C",
			x"0000" when x"954D",
			x"0000" when x"954E",
			x"0000" when x"954F",
			x"0000" when x"9550",
			x"0000" when x"9551",
			x"0000" when x"9552",
			x"0000" when x"9553",
			x"0000" when x"9554",
			x"0000" when x"9555",
			x"0000" when x"9556",
			x"0000" when x"9557",
			x"0000" when x"9558",
			x"0000" when x"9559",
			x"0000" when x"955A",
			x"0000" when x"955B",
			x"0000" when x"955C",
			x"0000" when x"955D",
			x"0000" when x"955E",
			x"0000" when x"955F",
			x"0000" when x"9560",
			x"0000" when x"9561",
			x"0000" when x"9562",
			x"0000" when x"9563",
			x"0000" when x"9564",
			x"0000" when x"9565",
			x"0000" when x"9566",
			x"0000" when x"9567",
			x"0000" when x"9568",
			x"0000" when x"9569",
			x"0000" when x"956A",
			x"0000" when x"956B",
			x"0000" when x"956C",
			x"0000" when x"956D",
			x"0000" when x"956E",
			x"0000" when x"956F",
			x"0000" when x"9570",
			x"0000" when x"9571",
			x"0000" when x"9572",
			x"0000" when x"9573",
			x"0000" when x"9574",
			x"0000" when x"9575",
			x"0000" when x"9576",
			x"0000" when x"9577",
			x"0000" when x"9578",
			x"0000" when x"9579",
			x"0000" when x"957A",
			x"0000" when x"957B",
			x"0000" when x"957C",
			x"0000" when x"957D",
			x"0000" when x"957E",
			x"0000" when x"957F",
			x"0000" when x"9580",
			x"0000" when x"9581",
			x"0000" when x"9582",
			x"0000" when x"9583",
			x"0000" when x"9584",
			x"0000" when x"9585",
			x"0000" when x"9586",
			x"0000" when x"9587",
			x"0000" when x"9588",
			x"0000" when x"9589",
			x"0000" when x"958A",
			x"0000" when x"958B",
			x"0000" when x"958C",
			x"0000" when x"958D",
			x"0000" when x"958E",
			x"0000" when x"958F",
			x"0000" when x"9590",
			x"0000" when x"9591",
			x"0000" when x"9592",
			x"0000" when x"9593",
			x"0000" when x"9594",
			x"0000" when x"9595",
			x"0000" when x"9596",
			x"0000" when x"9597",
			x"0000" when x"9598",
			x"0000" when x"9599",
			x"0000" when x"959A",
			x"0000" when x"959B",
			x"0000" when x"959C",
			x"0000" when x"959D",
			x"0000" when x"959E",
			x"0000" when x"959F",
			x"0000" when x"95A0",
			x"0000" when x"95A1",
			x"0000" when x"95A2",
			x"0000" when x"95A3",
			x"0000" when x"95A4",
			x"0000" when x"95A5",
			x"0000" when x"95A6",
			x"0000" when x"95A7",
			x"0000" when x"95A8",
			x"0000" when x"95A9",
			x"0000" when x"95AA",
			x"0000" when x"95AB",
			x"0000" when x"95AC",
			x"0000" when x"95AD",
			x"0000" when x"95AE",
			x"0000" when x"95AF",
			x"0000" when x"95B0",
			x"0000" when x"95B1",
			x"0000" when x"95B2",
			x"0000" when x"95B3",
			x"0000" when x"95B4",
			x"0000" when x"95B5",
			x"0000" when x"95B6",
			x"0000" when x"95B7",
			x"0000" when x"95B8",
			x"0000" when x"95B9",
			x"0000" when x"95BA",
			x"0000" when x"95BB",
			x"0000" when x"95BC",
			x"0000" when x"95BD",
			x"0000" when x"95BE",
			x"0000" when x"95BF",
			x"0000" when x"95C0",
			x"0000" when x"95C1",
			x"0000" when x"95C2",
			x"0000" when x"95C3",
			x"0000" when x"95C4",
			x"0000" when x"95C5",
			x"0000" when x"95C6",
			x"0000" when x"95C7",
			x"0000" when x"95C8",
			x"0000" when x"95C9",
			x"0000" when x"95CA",
			x"0000" when x"95CB",
			x"0000" when x"95CC",
			x"0000" when x"95CD",
			x"0000" when x"95CE",
			x"0000" when x"95CF",
			x"0000" when x"95D0",
			x"0000" when x"95D1",
			x"0000" when x"95D2",
			x"0000" when x"95D3",
			x"0000" when x"95D4",
			x"0000" when x"95D5",
			x"0000" when x"95D6",
			x"0000" when x"95D7",
			x"0000" when x"95D8",
			x"0000" when x"95D9",
			x"0000" when x"95DA",
			x"0000" when x"95DB",
			x"0000" when x"95DC",
			x"0000" when x"95DD",
			x"0000" when x"95DE",
			x"0000" when x"95DF",
			x"0000" when x"95E0",
			x"0000" when x"95E1",
			x"0000" when x"95E2",
			x"0000" when x"95E3",
			x"0000" when x"95E4",
			x"0000" when x"95E5",
			x"0000" when x"95E6",
			x"0000" when x"95E7",
			x"0000" when x"95E8",
			x"0000" when x"95E9",
			x"0000" when x"95EA",
			x"0000" when x"95EB",
			x"0000" when x"95EC",
			x"0000" when x"95ED",
			x"0000" when x"95EE",
			x"0000" when x"95EF",
			x"0000" when x"95F0",
			x"0000" when x"95F1",
			x"0000" when x"95F2",
			x"0000" when x"95F3",
			x"0000" when x"95F4",
			x"0000" when x"95F5",
			x"0000" when x"95F6",
			x"0000" when x"95F7",
			x"0000" when x"95F8",
			x"0000" when x"95F9",
			x"0000" when x"95FA",
			x"0000" when x"95FB",
			x"0000" when x"95FC",
			x"0000" when x"95FD",
			x"0000" when x"95FE",
			x"0000" when x"95FF",
			x"0000" when x"9600",
			x"0000" when x"9601",
			x"0000" when x"9602",
			x"0000" when x"9603",
			x"0000" when x"9604",
			x"0000" when x"9605",
			x"0000" when x"9606",
			x"0000" when x"9607",
			x"0000" when x"9608",
			x"0000" when x"9609",
			x"0000" when x"960A",
			x"0000" when x"960B",
			x"0000" when x"960C",
			x"0000" when x"960D",
			x"0000" when x"960E",
			x"0000" when x"960F",
			x"0000" when x"9610",
			x"0000" when x"9611",
			x"0000" when x"9612",
			x"0000" when x"9613",
			x"0000" when x"9614",
			x"0000" when x"9615",
			x"0000" when x"9616",
			x"0000" when x"9617",
			x"0000" when x"9618",
			x"0000" when x"9619",
			x"0000" when x"961A",
			x"0000" when x"961B",
			x"0000" when x"961C",
			x"0000" when x"961D",
			x"0000" when x"961E",
			x"0000" when x"961F",
			x"0000" when x"9620",
			x"0000" when x"9621",
			x"0000" when x"9622",
			x"0000" when x"9623",
			x"0000" when x"9624",
			x"0000" when x"9625",
			x"0000" when x"9626",
			x"0000" when x"9627",
			x"0000" when x"9628",
			x"0000" when x"9629",
			x"0000" when x"962A",
			x"0000" when x"962B",
			x"0000" when x"962C",
			x"0000" when x"962D",
			x"0000" when x"962E",
			x"0000" when x"962F",
			x"0000" when x"9630",
			x"0000" when x"9631",
			x"0000" when x"9632",
			x"0000" when x"9633",
			x"0000" when x"9634",
			x"0000" when x"9635",
			x"0000" when x"9636",
			x"0000" when x"9637",
			x"0000" when x"9638",
			x"0000" when x"9639",
			x"0000" when x"963A",
			x"0000" when x"963B",
			x"0000" when x"963C",
			x"0000" when x"963D",
			x"0000" when x"963E",
			x"0000" when x"963F",
			x"0000" when x"9640",
			x"0000" when x"9641",
			x"0000" when x"9642",
			x"0000" when x"9643",
			x"0000" when x"9644",
			x"0000" when x"9645",
			x"0000" when x"9646",
			x"0000" when x"9647",
			x"0000" when x"9648",
			x"0000" when x"9649",
			x"0000" when x"964A",
			x"0000" when x"964B",
			x"0000" when x"964C",
			x"0000" when x"964D",
			x"0000" when x"964E",
			x"0000" when x"964F",
			x"0000" when x"9650",
			x"0000" when x"9651",
			x"0000" when x"9652",
			x"0000" when x"9653",
			x"0000" when x"9654",
			x"0000" when x"9655",
			x"0000" when x"9656",
			x"0000" when x"9657",
			x"0000" when x"9658",
			x"0000" when x"9659",
			x"0000" when x"965A",
			x"0000" when x"965B",
			x"0000" when x"965C",
			x"0000" when x"965D",
			x"0000" when x"965E",
			x"0000" when x"965F",
			x"0000" when x"9660",
			x"0000" when x"9661",
			x"0000" when x"9662",
			x"0000" when x"9663",
			x"0000" when x"9664",
			x"0000" when x"9665",
			x"0000" when x"9666",
			x"0000" when x"9667",
			x"0000" when x"9668",
			x"0000" when x"9669",
			x"0000" when x"966A",
			x"0000" when x"966B",
			x"0000" when x"966C",
			x"0000" when x"966D",
			x"0000" when x"966E",
			x"0000" when x"966F",
			x"0000" when x"9670",
			x"0000" when x"9671",
			x"0000" when x"9672",
			x"0000" when x"9673",
			x"0000" when x"9674",
			x"0000" when x"9675",
			x"0000" when x"9676",
			x"0000" when x"9677",
			x"0000" when x"9678",
			x"0000" when x"9679",
			x"0000" when x"967A",
			x"0000" when x"967B",
			x"0000" when x"967C",
			x"0000" when x"967D",
			x"0000" when x"967E",
			x"0000" when x"967F",
			x"0000" when x"9680",
			x"0000" when x"9681",
			x"0000" when x"9682",
			x"0000" when x"9683",
			x"0000" when x"9684",
			x"0000" when x"9685",
			x"0000" when x"9686",
			x"0000" when x"9687",
			x"0000" when x"9688",
			x"0000" when x"9689",
			x"0000" when x"968A",
			x"0000" when x"968B",
			x"0000" when x"968C",
			x"0000" when x"968D",
			x"0000" when x"968E",
			x"0000" when x"968F",
			x"0000" when x"9690",
			x"0000" when x"9691",
			x"0000" when x"9692",
			x"0000" when x"9693",
			x"0000" when x"9694",
			x"0000" when x"9695",
			x"0000" when x"9696",
			x"0000" when x"9697",
			x"0000" when x"9698",
			x"0000" when x"9699",
			x"0000" when x"969A",
			x"0000" when x"969B",
			x"0000" when x"969C",
			x"0000" when x"969D",
			x"0000" when x"969E",
			x"0000" when x"969F",
			x"0000" when x"96A0",
			x"0000" when x"96A1",
			x"0000" when x"96A2",
			x"0000" when x"96A3",
			x"0000" when x"96A4",
			x"0000" when x"96A5",
			x"0000" when x"96A6",
			x"0000" when x"96A7",
			x"0000" when x"96A8",
			x"0000" when x"96A9",
			x"0000" when x"96AA",
			x"0000" when x"96AB",
			x"0000" when x"96AC",
			x"0000" when x"96AD",
			x"0000" when x"96AE",
			x"0000" when x"96AF",
			x"0000" when x"96B0",
			x"0000" when x"96B1",
			x"0000" when x"96B2",
			x"0000" when x"96B3",
			x"0000" when x"96B4",
			x"0000" when x"96B5",
			x"0000" when x"96B6",
			x"0000" when x"96B7",
			x"0000" when x"96B8",
			x"0000" when x"96B9",
			x"0000" when x"96BA",
			x"0000" when x"96BB",
			x"0000" when x"96BC",
			x"0000" when x"96BD",
			x"0000" when x"96BE",
			x"0000" when x"96BF",
			x"0000" when x"96C0",
			x"0000" when x"96C1",
			x"0000" when x"96C2",
			x"0000" when x"96C3",
			x"0000" when x"96C4",
			x"0000" when x"96C5",
			x"0000" when x"96C6",
			x"0000" when x"96C7",
			x"0000" when x"96C8",
			x"0000" when x"96C9",
			x"0000" when x"96CA",
			x"0000" when x"96CB",
			x"0000" when x"96CC",
			x"0000" when x"96CD",
			x"0000" when x"96CE",
			x"0000" when x"96CF",
			x"0000" when x"96D0",
			x"0000" when x"96D1",
			x"0000" when x"96D2",
			x"0000" when x"96D3",
			x"0000" when x"96D4",
			x"0000" when x"96D5",
			x"0000" when x"96D6",
			x"0000" when x"96D7",
			x"0000" when x"96D8",
			x"0000" when x"96D9",
			x"0000" when x"96DA",
			x"0000" when x"96DB",
			x"0000" when x"96DC",
			x"0000" when x"96DD",
			x"0000" when x"96DE",
			x"0000" when x"96DF",
			x"0000" when x"96E0",
			x"0000" when x"96E1",
			x"0000" when x"96E2",
			x"0000" when x"96E3",
			x"0000" when x"96E4",
			x"0000" when x"96E5",
			x"0000" when x"96E6",
			x"0000" when x"96E7",
			x"0000" when x"96E8",
			x"0000" when x"96E9",
			x"0000" when x"96EA",
			x"0000" when x"96EB",
			x"0000" when x"96EC",
			x"0000" when x"96ED",
			x"0000" when x"96EE",
			x"0000" when x"96EF",
			x"0000" when x"96F0",
			x"0000" when x"96F1",
			x"0000" when x"96F2",
			x"0000" when x"96F3",
			x"0000" when x"96F4",
			x"0000" when x"96F5",
			x"0000" when x"96F6",
			x"0000" when x"96F7",
			x"0000" when x"96F8",
			x"0000" when x"96F9",
			x"0000" when x"96FA",
			x"0000" when x"96FB",
			x"0000" when x"96FC",
			x"0000" when x"96FD",
			x"0000" when x"96FE",
			x"0000" when x"96FF",
			x"0000" when x"9700",
			x"0000" when x"9701",
			x"0000" when x"9702",
			x"0000" when x"9703",
			x"0000" when x"9704",
			x"0000" when x"9705",
			x"0000" when x"9706",
			x"0000" when x"9707",
			x"0000" when x"9708",
			x"0000" when x"9709",
			x"0000" when x"970A",
			x"0000" when x"970B",
			x"0000" when x"970C",
			x"0000" when x"970D",
			x"0000" when x"970E",
			x"0000" when x"970F",
			x"0000" when x"9710",
			x"0000" when x"9711",
			x"0000" when x"9712",
			x"0000" when x"9713",
			x"0000" when x"9714",
			x"0000" when x"9715",
			x"0000" when x"9716",
			x"0000" when x"9717",
			x"0000" when x"9718",
			x"0000" when x"9719",
			x"0000" when x"971A",
			x"0000" when x"971B",
			x"0000" when x"971C",
			x"0000" when x"971D",
			x"0000" when x"971E",
			x"0000" when x"971F",
			x"0000" when x"9720",
			x"0000" when x"9721",
			x"0000" when x"9722",
			x"0000" when x"9723",
			x"0000" when x"9724",
			x"0000" when x"9725",
			x"0000" when x"9726",
			x"0000" when x"9727",
			x"0000" when x"9728",
			x"0000" when x"9729",
			x"0000" when x"972A",
			x"0000" when x"972B",
			x"0000" when x"972C",
			x"0000" when x"972D",
			x"0000" when x"972E",
			x"0000" when x"972F",
			x"0000" when x"9730",
			x"0000" when x"9731",
			x"0000" when x"9732",
			x"0000" when x"9733",
			x"0000" when x"9734",
			x"0000" when x"9735",
			x"0000" when x"9736",
			x"0000" when x"9737",
			x"0000" when x"9738",
			x"0000" when x"9739",
			x"0000" when x"973A",
			x"0000" when x"973B",
			x"0000" when x"973C",
			x"0000" when x"973D",
			x"0000" when x"973E",
			x"0000" when x"973F",
			x"0000" when x"9740",
			x"0000" when x"9741",
			x"0000" when x"9742",
			x"0000" when x"9743",
			x"0000" when x"9744",
			x"0000" when x"9745",
			x"0000" when x"9746",
			x"0000" when x"9747",
			x"0000" when x"9748",
			x"0000" when x"9749",
			x"0000" when x"974A",
			x"0000" when x"974B",
			x"0000" when x"974C",
			x"0000" when x"974D",
			x"0000" when x"974E",
			x"0000" when x"974F",
			x"0000" when x"9750",
			x"0000" when x"9751",
			x"0000" when x"9752",
			x"0000" when x"9753",
			x"0000" when x"9754",
			x"0000" when x"9755",
			x"0000" when x"9756",
			x"0000" when x"9757",
			x"0000" when x"9758",
			x"0000" when x"9759",
			x"0000" when x"975A",
			x"0000" when x"975B",
			x"0000" when x"975C",
			x"0000" when x"975D",
			x"0000" when x"975E",
			x"0000" when x"975F",
			x"0000" when x"9760",
			x"0000" when x"9761",
			x"0000" when x"9762",
			x"0000" when x"9763",
			x"0000" when x"9764",
			x"0000" when x"9765",
			x"0000" when x"9766",
			x"0000" when x"9767",
			x"0000" when x"9768",
			x"0000" when x"9769",
			x"0000" when x"976A",
			x"0000" when x"976B",
			x"0000" when x"976C",
			x"0000" when x"976D",
			x"0000" when x"976E",
			x"0000" when x"976F",
			x"0000" when x"9770",
			x"0000" when x"9771",
			x"0000" when x"9772",
			x"0000" when x"9773",
			x"0000" when x"9774",
			x"0000" when x"9775",
			x"0000" when x"9776",
			x"0000" when x"9777",
			x"0000" when x"9778",
			x"0000" when x"9779",
			x"0000" when x"977A",
			x"0000" when x"977B",
			x"0000" when x"977C",
			x"0000" when x"977D",
			x"0000" when x"977E",
			x"0000" when x"977F",
			x"0000" when x"9780",
			x"0000" when x"9781",
			x"0000" when x"9782",
			x"0000" when x"9783",
			x"0000" when x"9784",
			x"0000" when x"9785",
			x"0000" when x"9786",
			x"0000" when x"9787",
			x"0000" when x"9788",
			x"0000" when x"9789",
			x"0000" when x"978A",
			x"0000" when x"978B",
			x"0000" when x"978C",
			x"0000" when x"978D",
			x"0000" when x"978E",
			x"0000" when x"978F",
			x"0000" when x"9790",
			x"0000" when x"9791",
			x"0000" when x"9792",
			x"0000" when x"9793",
			x"0000" when x"9794",
			x"0000" when x"9795",
			x"0000" when x"9796",
			x"0000" when x"9797",
			x"0000" when x"9798",
			x"0000" when x"9799",
			x"0000" when x"979A",
			x"0000" when x"979B",
			x"0000" when x"979C",
			x"0000" when x"979D",
			x"0000" when x"979E",
			x"0000" when x"979F",
			x"0000" when x"97A0",
			x"0000" when x"97A1",
			x"0000" when x"97A2",
			x"0000" when x"97A3",
			x"0000" when x"97A4",
			x"0000" when x"97A5",
			x"0000" when x"97A6",
			x"0000" when x"97A7",
			x"0000" when x"97A8",
			x"0000" when x"97A9",
			x"0000" when x"97AA",
			x"0000" when x"97AB",
			x"0000" when x"97AC",
			x"0000" when x"97AD",
			x"0000" when x"97AE",
			x"0000" when x"97AF",
			x"0000" when x"97B0",
			x"0000" when x"97B1",
			x"0000" when x"97B2",
			x"0000" when x"97B3",
			x"0000" when x"97B4",
			x"0000" when x"97B5",
			x"0000" when x"97B6",
			x"0000" when x"97B7",
			x"0000" when x"97B8",
			x"0000" when x"97B9",
			x"0000" when x"97BA",
			x"0000" when x"97BB",
			x"0000" when x"97BC",
			x"0000" when x"97BD",
			x"0000" when x"97BE",
			x"0000" when x"97BF",
			x"0000" when x"97C0",
			x"0000" when x"97C1",
			x"0000" when x"97C2",
			x"0000" when x"97C3",
			x"0000" when x"97C4",
			x"0000" when x"97C5",
			x"0000" when x"97C6",
			x"0000" when x"97C7",
			x"0000" when x"97C8",
			x"0000" when x"97C9",
			x"0000" when x"97CA",
			x"0000" when x"97CB",
			x"0000" when x"97CC",
			x"0000" when x"97CD",
			x"0000" when x"97CE",
			x"0000" when x"97CF",
			x"0000" when x"97D0",
			x"0000" when x"97D1",
			x"0000" when x"97D2",
			x"0000" when x"97D3",
			x"0000" when x"97D4",
			x"0000" when x"97D5",
			x"0000" when x"97D6",
			x"0000" when x"97D7",
			x"0000" when x"97D8",
			x"0000" when x"97D9",
			x"0000" when x"97DA",
			x"0000" when x"97DB",
			x"0000" when x"97DC",
			x"0000" when x"97DD",
			x"0000" when x"97DE",
			x"0000" when x"97DF",
			x"0000" when x"97E0",
			x"0000" when x"97E1",
			x"0000" when x"97E2",
			x"0000" when x"97E3",
			x"0000" when x"97E4",
			x"0000" when x"97E5",
			x"0000" when x"97E6",
			x"0000" when x"97E7",
			x"0000" when x"97E8",
			x"0000" when x"97E9",
			x"0000" when x"97EA",
			x"0000" when x"97EB",
			x"0000" when x"97EC",
			x"0000" when x"97ED",
			x"0000" when x"97EE",
			x"0000" when x"97EF",
			x"0000" when x"97F0",
			x"0000" when x"97F1",
			x"0000" when x"97F2",
			x"0000" when x"97F3",
			x"0000" when x"97F4",
			x"0000" when x"97F5",
			x"0000" when x"97F6",
			x"0000" when x"97F7",
			x"0000" when x"97F8",
			x"0000" when x"97F9",
			x"0000" when x"97FA",
			x"0000" when x"97FB",
			x"0000" when x"97FC",
			x"0000" when x"97FD",
			x"0000" when x"97FE",
			x"0000" when x"97FF",
			x"0000" when x"9800",
			x"0000" when x"9801",
			x"0000" when x"9802",
			x"0000" when x"9803",
			x"0000" when x"9804",
			x"0000" when x"9805",
			x"0000" when x"9806",
			x"0000" when x"9807",
			x"0000" when x"9808",
			x"0000" when x"9809",
			x"0000" when x"980A",
			x"0000" when x"980B",
			x"0000" when x"980C",
			x"0000" when x"980D",
			x"0000" when x"980E",
			x"0000" when x"980F",
			x"0000" when x"9810",
			x"0000" when x"9811",
			x"0000" when x"9812",
			x"0000" when x"9813",
			x"0000" when x"9814",
			x"0000" when x"9815",
			x"0000" when x"9816",
			x"0000" when x"9817",
			x"0000" when x"9818",
			x"0000" when x"9819",
			x"0000" when x"981A",
			x"0000" when x"981B",
			x"0000" when x"981C",
			x"0000" when x"981D",
			x"0000" when x"981E",
			x"0000" when x"981F",
			x"0000" when x"9820",
			x"0000" when x"9821",
			x"0000" when x"9822",
			x"0000" when x"9823",
			x"0000" when x"9824",
			x"0000" when x"9825",
			x"0000" when x"9826",
			x"0000" when x"9827",
			x"0000" when x"9828",
			x"0000" when x"9829",
			x"0000" when x"982A",
			x"0000" when x"982B",
			x"0000" when x"982C",
			x"0000" when x"982D",
			x"0000" when x"982E",
			x"0000" when x"982F",
			x"0000" when x"9830",
			x"0000" when x"9831",
			x"0000" when x"9832",
			x"0000" when x"9833",
			x"0000" when x"9834",
			x"0000" when x"9835",
			x"0000" when x"9836",
			x"0000" when x"9837",
			x"0000" when x"9838",
			x"0000" when x"9839",
			x"0000" when x"983A",
			x"0000" when x"983B",
			x"0000" when x"983C",
			x"0000" when x"983D",
			x"0000" when x"983E",
			x"0000" when x"983F",
			x"0000" when x"9840",
			x"0000" when x"9841",
			x"0000" when x"9842",
			x"0000" when x"9843",
			x"0000" when x"9844",
			x"0000" when x"9845",
			x"0000" when x"9846",
			x"0000" when x"9847",
			x"0000" when x"9848",
			x"0000" when x"9849",
			x"0000" when x"984A",
			x"0000" when x"984B",
			x"0000" when x"984C",
			x"0000" when x"984D",
			x"0000" when x"984E",
			x"0000" when x"984F",
			x"0000" when x"9850",
			x"0000" when x"9851",
			x"0000" when x"9852",
			x"0000" when x"9853",
			x"0000" when x"9854",
			x"0000" when x"9855",
			x"0000" when x"9856",
			x"0000" when x"9857",
			x"0000" when x"9858",
			x"0000" when x"9859",
			x"0000" when x"985A",
			x"0000" when x"985B",
			x"0000" when x"985C",
			x"0000" when x"985D",
			x"0000" when x"985E",
			x"0000" when x"985F",
			x"0000" when x"9860",
			x"0000" when x"9861",
			x"0000" when x"9862",
			x"0000" when x"9863",
			x"0000" when x"9864",
			x"0000" when x"9865",
			x"0000" when x"9866",
			x"0000" when x"9867",
			x"0000" when x"9868",
			x"0000" when x"9869",
			x"0000" when x"986A",
			x"0000" when x"986B",
			x"0000" when x"986C",
			x"0000" when x"986D",
			x"0000" when x"986E",
			x"0000" when x"986F",
			x"0000" when x"9870",
			x"0000" when x"9871",
			x"0000" when x"9872",
			x"0000" when x"9873",
			x"0000" when x"9874",
			x"0000" when x"9875",
			x"0000" when x"9876",
			x"0000" when x"9877",
			x"0000" when x"9878",
			x"0000" when x"9879",
			x"0000" when x"987A",
			x"0000" when x"987B",
			x"0000" when x"987C",
			x"0000" when x"987D",
			x"0000" when x"987E",
			x"0000" when x"987F",
			x"0000" when x"9880",
			x"0000" when x"9881",
			x"0000" when x"9882",
			x"0000" when x"9883",
			x"0000" when x"9884",
			x"0000" when x"9885",
			x"0000" when x"9886",
			x"0000" when x"9887",
			x"0000" when x"9888",
			x"0000" when x"9889",
			x"0000" when x"988A",
			x"0000" when x"988B",
			x"0000" when x"988C",
			x"0000" when x"988D",
			x"0000" when x"988E",
			x"0000" when x"988F",
			x"0000" when x"9890",
			x"0000" when x"9891",
			x"0000" when x"9892",
			x"0000" when x"9893",
			x"0000" when x"9894",
			x"0000" when x"9895",
			x"0000" when x"9896",
			x"0000" when x"9897",
			x"0000" when x"9898",
			x"0000" when x"9899",
			x"0000" when x"989A",
			x"0000" when x"989B",
			x"0000" when x"989C",
			x"0000" when x"989D",
			x"0000" when x"989E",
			x"0000" when x"989F",
			x"0000" when x"98A0",
			x"0000" when x"98A1",
			x"0000" when x"98A2",
			x"0000" when x"98A3",
			x"0000" when x"98A4",
			x"0000" when x"98A5",
			x"0000" when x"98A6",
			x"0000" when x"98A7",
			x"0000" when x"98A8",
			x"0000" when x"98A9",
			x"0000" when x"98AA",
			x"0000" when x"98AB",
			x"0000" when x"98AC",
			x"0000" when x"98AD",
			x"0000" when x"98AE",
			x"0000" when x"98AF",
			x"0000" when x"98B0",
			x"0000" when x"98B1",
			x"0000" when x"98B2",
			x"0000" when x"98B3",
			x"0000" when x"98B4",
			x"0000" when x"98B5",
			x"0000" when x"98B6",
			x"0000" when x"98B7",
			x"0000" when x"98B8",
			x"0000" when x"98B9",
			x"0000" when x"98BA",
			x"0000" when x"98BB",
			x"0000" when x"98BC",
			x"0000" when x"98BD",
			x"0000" when x"98BE",
			x"0000" when x"98BF",
			x"0000" when x"98C0",
			x"0000" when x"98C1",
			x"0000" when x"98C2",
			x"0000" when x"98C3",
			x"0000" when x"98C4",
			x"0000" when x"98C5",
			x"0000" when x"98C6",
			x"0000" when x"98C7",
			x"0000" when x"98C8",
			x"0000" when x"98C9",
			x"0000" when x"98CA",
			x"0000" when x"98CB",
			x"0000" when x"98CC",
			x"0000" when x"98CD",
			x"0000" when x"98CE",
			x"0000" when x"98CF",
			x"0000" when x"98D0",
			x"0000" when x"98D1",
			x"0000" when x"98D2",
			x"0000" when x"98D3",
			x"0000" when x"98D4",
			x"0000" when x"98D5",
			x"0000" when x"98D6",
			x"0000" when x"98D7",
			x"0000" when x"98D8",
			x"0000" when x"98D9",
			x"0000" when x"98DA",
			x"0000" when x"98DB",
			x"0000" when x"98DC",
			x"0000" when x"98DD",
			x"0000" when x"98DE",
			x"0000" when x"98DF",
			x"0000" when x"98E0",
			x"0000" when x"98E1",
			x"0000" when x"98E2",
			x"0000" when x"98E3",
			x"0000" when x"98E4",
			x"0000" when x"98E5",
			x"0000" when x"98E6",
			x"0000" when x"98E7",
			x"0000" when x"98E8",
			x"0000" when x"98E9",
			x"0000" when x"98EA",
			x"0000" when x"98EB",
			x"0000" when x"98EC",
			x"0000" when x"98ED",
			x"0000" when x"98EE",
			x"0000" when x"98EF",
			x"0000" when x"98F0",
			x"0000" when x"98F1",
			x"0000" when x"98F2",
			x"0000" when x"98F3",
			x"0000" when x"98F4",
			x"0000" when x"98F5",
			x"0000" when x"98F6",
			x"0000" when x"98F7",
			x"0000" when x"98F8",
			x"0000" when x"98F9",
			x"0000" when x"98FA",
			x"0000" when x"98FB",
			x"0000" when x"98FC",
			x"0000" when x"98FD",
			x"0000" when x"98FE",
			x"0000" when x"98FF",
			x"0000" when x"9900",
			x"0000" when x"9901",
			x"0000" when x"9902",
			x"0000" when x"9903",
			x"0000" when x"9904",
			x"0000" when x"9905",
			x"0000" when x"9906",
			x"0000" when x"9907",
			x"0000" when x"9908",
			x"0000" when x"9909",
			x"0000" when x"990A",
			x"0000" when x"990B",
			x"0000" when x"990C",
			x"0000" when x"990D",
			x"0000" when x"990E",
			x"0000" when x"990F",
			x"0000" when x"9910",
			x"0000" when x"9911",
			x"0000" when x"9912",
			x"0000" when x"9913",
			x"0000" when x"9914",
			x"0000" when x"9915",
			x"0000" when x"9916",
			x"0000" when x"9917",
			x"0000" when x"9918",
			x"0000" when x"9919",
			x"0000" when x"991A",
			x"0000" when x"991B",
			x"0000" when x"991C",
			x"0000" when x"991D",
			x"0000" when x"991E",
			x"0000" when x"991F",
			x"0000" when x"9920",
			x"0000" when x"9921",
			x"0000" when x"9922",
			x"0000" when x"9923",
			x"0000" when x"9924",
			x"0000" when x"9925",
			x"0000" when x"9926",
			x"0000" when x"9927",
			x"0000" when x"9928",
			x"0000" when x"9929",
			x"0000" when x"992A",
			x"0000" when x"992B",
			x"0000" when x"992C",
			x"0000" when x"992D",
			x"0000" when x"992E",
			x"0000" when x"992F",
			x"0000" when x"9930",
			x"0000" when x"9931",
			x"0000" when x"9932",
			x"0000" when x"9933",
			x"0000" when x"9934",
			x"0000" when x"9935",
			x"0000" when x"9936",
			x"0000" when x"9937",
			x"0000" when x"9938",
			x"0000" when x"9939",
			x"0000" when x"993A",
			x"0000" when x"993B",
			x"0000" when x"993C",
			x"0000" when x"993D",
			x"0000" when x"993E",
			x"0000" when x"993F",
			x"0000" when x"9940",
			x"0000" when x"9941",
			x"0000" when x"9942",
			x"0000" when x"9943",
			x"0000" when x"9944",
			x"0000" when x"9945",
			x"0000" when x"9946",
			x"0000" when x"9947",
			x"0000" when x"9948",
			x"0000" when x"9949",
			x"0000" when x"994A",
			x"0000" when x"994B",
			x"0000" when x"994C",
			x"0000" when x"994D",
			x"0000" when x"994E",
			x"0000" when x"994F",
			x"0000" when x"9950",
			x"0000" when x"9951",
			x"0000" when x"9952",
			x"0000" when x"9953",
			x"0000" when x"9954",
			x"0000" when x"9955",
			x"0000" when x"9956",
			x"0000" when x"9957",
			x"0000" when x"9958",
			x"0000" when x"9959",
			x"0000" when x"995A",
			x"0000" when x"995B",
			x"0000" when x"995C",
			x"0000" when x"995D",
			x"0000" when x"995E",
			x"0000" when x"995F",
			x"0000" when x"9960",
			x"0000" when x"9961",
			x"0000" when x"9962",
			x"0000" when x"9963",
			x"0000" when x"9964",
			x"0000" when x"9965",
			x"0000" when x"9966",
			x"0000" when x"9967",
			x"0000" when x"9968",
			x"0000" when x"9969",
			x"0000" when x"996A",
			x"0000" when x"996B",
			x"0000" when x"996C",
			x"0000" when x"996D",
			x"0000" when x"996E",
			x"0000" when x"996F",
			x"0000" when x"9970",
			x"0000" when x"9971",
			x"0000" when x"9972",
			x"0000" when x"9973",
			x"0000" when x"9974",
			x"0000" when x"9975",
			x"0000" when x"9976",
			x"0000" when x"9977",
			x"0000" when x"9978",
			x"0000" when x"9979",
			x"0000" when x"997A",
			x"0000" when x"997B",
			x"0000" when x"997C",
			x"0000" when x"997D",
			x"0000" when x"997E",
			x"0000" when x"997F",
			x"0000" when x"9980",
			x"0000" when x"9981",
			x"0000" when x"9982",
			x"0000" when x"9983",
			x"0000" when x"9984",
			x"0000" when x"9985",
			x"0000" when x"9986",
			x"0000" when x"9987",
			x"0000" when x"9988",
			x"0000" when x"9989",
			x"0000" when x"998A",
			x"0000" when x"998B",
			x"0000" when x"998C",
			x"0000" when x"998D",
			x"0000" when x"998E",
			x"0000" when x"998F",
			x"0000" when x"9990",
			x"0000" when x"9991",
			x"0000" when x"9992",
			x"0000" when x"9993",
			x"0000" when x"9994",
			x"0000" when x"9995",
			x"0000" when x"9996",
			x"0000" when x"9997",
			x"0000" when x"9998",
			x"0000" when x"9999",
			x"0000" when x"999A",
			x"0000" when x"999B",
			x"0000" when x"999C",
			x"0000" when x"999D",
			x"0000" when x"999E",
			x"0000" when x"999F",
			x"0000" when x"99A0",
			x"0000" when x"99A1",
			x"0000" when x"99A2",
			x"0000" when x"99A3",
			x"0000" when x"99A4",
			x"0000" when x"99A5",
			x"0000" when x"99A6",
			x"0000" when x"99A7",
			x"0000" when x"99A8",
			x"0000" when x"99A9",
			x"0000" when x"99AA",
			x"0000" when x"99AB",
			x"0000" when x"99AC",
			x"0000" when x"99AD",
			x"0000" when x"99AE",
			x"0000" when x"99AF",
			x"0000" when x"99B0",
			x"0000" when x"99B1",
			x"0000" when x"99B2",
			x"0000" when x"99B3",
			x"0000" when x"99B4",
			x"0000" when x"99B5",
			x"0000" when x"99B6",
			x"0000" when x"99B7",
			x"0000" when x"99B8",
			x"0000" when x"99B9",
			x"0000" when x"99BA",
			x"0000" when x"99BB",
			x"0000" when x"99BC",
			x"0000" when x"99BD",
			x"0000" when x"99BE",
			x"0000" when x"99BF",
			x"0000" when x"99C0",
			x"0000" when x"99C1",
			x"0000" when x"99C2",
			x"0000" when x"99C3",
			x"0000" when x"99C4",
			x"0000" when x"99C5",
			x"0000" when x"99C6",
			x"0000" when x"99C7",
			x"0000" when x"99C8",
			x"0000" when x"99C9",
			x"0000" when x"99CA",
			x"0000" when x"99CB",
			x"0000" when x"99CC",
			x"0000" when x"99CD",
			x"0000" when x"99CE",
			x"0000" when x"99CF",
			x"0000" when x"99D0",
			x"0000" when x"99D1",
			x"0000" when x"99D2",
			x"0000" when x"99D3",
			x"0000" when x"99D4",
			x"0000" when x"99D5",
			x"0000" when x"99D6",
			x"0000" when x"99D7",
			x"0000" when x"99D8",
			x"0000" when x"99D9",
			x"0000" when x"99DA",
			x"0000" when x"99DB",
			x"0000" when x"99DC",
			x"0000" when x"99DD",
			x"0000" when x"99DE",
			x"0000" when x"99DF",
			x"0000" when x"99E0",
			x"0000" when x"99E1",
			x"0000" when x"99E2",
			x"0000" when x"99E3",
			x"0000" when x"99E4",
			x"0000" when x"99E5",
			x"0000" when x"99E6",
			x"0000" when x"99E7",
			x"0000" when x"99E8",
			x"0000" when x"99E9",
			x"0000" when x"99EA",
			x"0000" when x"99EB",
			x"0000" when x"99EC",
			x"0000" when x"99ED",
			x"0000" when x"99EE",
			x"0000" when x"99EF",
			x"0000" when x"99F0",
			x"0000" when x"99F1",
			x"0000" when x"99F2",
			x"0000" when x"99F3",
			x"0000" when x"99F4",
			x"0000" when x"99F5",
			x"0000" when x"99F6",
			x"0000" when x"99F7",
			x"0000" when x"99F8",
			x"0000" when x"99F9",
			x"0000" when x"99FA",
			x"0000" when x"99FB",
			x"0000" when x"99FC",
			x"0000" when x"99FD",
			x"0000" when x"99FE",
			x"0000" when x"99FF",
			x"0000" when x"9A00",
			x"0000" when x"9A01",
			x"0000" when x"9A02",
			x"0000" when x"9A03",
			x"0000" when x"9A04",
			x"0000" when x"9A05",
			x"0000" when x"9A06",
			x"0000" when x"9A07",
			x"0000" when x"9A08",
			x"0000" when x"9A09",
			x"0000" when x"9A0A",
			x"0000" when x"9A0B",
			x"0000" when x"9A0C",
			x"0000" when x"9A0D",
			x"0000" when x"9A0E",
			x"0000" when x"9A0F",
			x"0000" when x"9A10",
			x"0000" when x"9A11",
			x"0000" when x"9A12",
			x"0000" when x"9A13",
			x"0000" when x"9A14",
			x"0000" when x"9A15",
			x"0000" when x"9A16",
			x"0000" when x"9A17",
			x"0000" when x"9A18",
			x"0000" when x"9A19",
			x"0000" when x"9A1A",
			x"0000" when x"9A1B",
			x"0000" when x"9A1C",
			x"0000" when x"9A1D",
			x"0000" when x"9A1E",
			x"0000" when x"9A1F",
			x"0000" when x"9A20",
			x"0000" when x"9A21",
			x"0000" when x"9A22",
			x"0000" when x"9A23",
			x"0000" when x"9A24",
			x"0000" when x"9A25",
			x"0000" when x"9A26",
			x"0000" when x"9A27",
			x"0000" when x"9A28",
			x"0000" when x"9A29",
			x"0000" when x"9A2A",
			x"0000" when x"9A2B",
			x"0000" when x"9A2C",
			x"0000" when x"9A2D",
			x"0000" when x"9A2E",
			x"0000" when x"9A2F",
			x"0000" when x"9A30",
			x"0000" when x"9A31",
			x"0000" when x"9A32",
			x"0000" when x"9A33",
			x"0000" when x"9A34",
			x"0000" when x"9A35",
			x"0000" when x"9A36",
			x"0000" when x"9A37",
			x"0000" when x"9A38",
			x"0000" when x"9A39",
			x"0000" when x"9A3A",
			x"0000" when x"9A3B",
			x"0000" when x"9A3C",
			x"0000" when x"9A3D",
			x"0000" when x"9A3E",
			x"0000" when x"9A3F",
			x"0000" when x"9A40",
			x"0000" when x"9A41",
			x"0000" when x"9A42",
			x"0000" when x"9A43",
			x"0000" when x"9A44",
			x"0000" when x"9A45",
			x"0000" when x"9A46",
			x"0000" when x"9A47",
			x"0000" when x"9A48",
			x"0000" when x"9A49",
			x"0000" when x"9A4A",
			x"0000" when x"9A4B",
			x"0000" when x"9A4C",
			x"0000" when x"9A4D",
			x"0000" when x"9A4E",
			x"0000" when x"9A4F",
			x"0000" when x"9A50",
			x"0000" when x"9A51",
			x"0000" when x"9A52",
			x"0000" when x"9A53",
			x"0000" when x"9A54",
			x"0000" when x"9A55",
			x"0000" when x"9A56",
			x"0000" when x"9A57",
			x"0000" when x"9A58",
			x"0000" when x"9A59",
			x"0000" when x"9A5A",
			x"0000" when x"9A5B",
			x"0000" when x"9A5C",
			x"0000" when x"9A5D",
			x"0000" when x"9A5E",
			x"0000" when x"9A5F",
			x"0000" when x"9A60",
			x"0000" when x"9A61",
			x"0000" when x"9A62",
			x"0000" when x"9A63",
			x"0000" when x"9A64",
			x"0000" when x"9A65",
			x"0000" when x"9A66",
			x"0000" when x"9A67",
			x"0000" when x"9A68",
			x"0000" when x"9A69",
			x"0000" when x"9A6A",
			x"0000" when x"9A6B",
			x"0000" when x"9A6C",
			x"0000" when x"9A6D",
			x"0000" when x"9A6E",
			x"0000" when x"9A6F",
			x"0000" when x"9A70",
			x"0000" when x"9A71",
			x"0000" when x"9A72",
			x"0000" when x"9A73",
			x"0000" when x"9A74",
			x"0000" when x"9A75",
			x"0000" when x"9A76",
			x"0000" when x"9A77",
			x"0000" when x"9A78",
			x"0000" when x"9A79",
			x"0000" when x"9A7A",
			x"0000" when x"9A7B",
			x"0000" when x"9A7C",
			x"0000" when x"9A7D",
			x"0000" when x"9A7E",
			x"0000" when x"9A7F",
			x"0000" when x"9A80",
			x"0000" when x"9A81",
			x"0000" when x"9A82",
			x"0000" when x"9A83",
			x"0000" when x"9A84",
			x"0000" when x"9A85",
			x"0000" when x"9A86",
			x"0000" when x"9A87",
			x"0000" when x"9A88",
			x"0000" when x"9A89",
			x"0000" when x"9A8A",
			x"0000" when x"9A8B",
			x"0000" when x"9A8C",
			x"0000" when x"9A8D",
			x"0000" when x"9A8E",
			x"0000" when x"9A8F",
			x"0000" when x"9A90",
			x"0000" when x"9A91",
			x"0000" when x"9A92",
			x"0000" when x"9A93",
			x"0000" when x"9A94",
			x"0000" when x"9A95",
			x"0000" when x"9A96",
			x"0000" when x"9A97",
			x"0000" when x"9A98",
			x"0000" when x"9A99",
			x"0000" when x"9A9A",
			x"0000" when x"9A9B",
			x"0000" when x"9A9C",
			x"0000" when x"9A9D",
			x"0000" when x"9A9E",
			x"0000" when x"9A9F",
			x"0000" when x"9AA0",
			x"0000" when x"9AA1",
			x"0000" when x"9AA2",
			x"0000" when x"9AA3",
			x"0000" when x"9AA4",
			x"0000" when x"9AA5",
			x"0000" when x"9AA6",
			x"0000" when x"9AA7",
			x"0000" when x"9AA8",
			x"0000" when x"9AA9",
			x"0000" when x"9AAA",
			x"0000" when x"9AAB",
			x"0000" when x"9AAC",
			x"0000" when x"9AAD",
			x"0000" when x"9AAE",
			x"0000" when x"9AAF",
			x"0000" when x"9AB0",
			x"0000" when x"9AB1",
			x"0000" when x"9AB2",
			x"0000" when x"9AB3",
			x"0000" when x"9AB4",
			x"0000" when x"9AB5",
			x"0000" when x"9AB6",
			x"0000" when x"9AB7",
			x"0000" when x"9AB8",
			x"0000" when x"9AB9",
			x"0000" when x"9ABA",
			x"0000" when x"9ABB",
			x"0000" when x"9ABC",
			x"0000" when x"9ABD",
			x"0000" when x"9ABE",
			x"0000" when x"9ABF",
			x"0000" when x"9AC0",
			x"0000" when x"9AC1",
			x"0000" when x"9AC2",
			x"0000" when x"9AC3",
			x"0000" when x"9AC4",
			x"0000" when x"9AC5",
			x"0000" when x"9AC6",
			x"0000" when x"9AC7",
			x"0000" when x"9AC8",
			x"0000" when x"9AC9",
			x"0000" when x"9ACA",
			x"0000" when x"9ACB",
			x"0000" when x"9ACC",
			x"0000" when x"9ACD",
			x"0000" when x"9ACE",
			x"0000" when x"9ACF",
			x"0000" when x"9AD0",
			x"0000" when x"9AD1",
			x"0000" when x"9AD2",
			x"0000" when x"9AD3",
			x"0000" when x"9AD4",
			x"0000" when x"9AD5",
			x"0000" when x"9AD6",
			x"0000" when x"9AD7",
			x"0000" when x"9AD8",
			x"0000" when x"9AD9",
			x"0000" when x"9ADA",
			x"0000" when x"9ADB",
			x"0000" when x"9ADC",
			x"0000" when x"9ADD",
			x"0000" when x"9ADE",
			x"0000" when x"9ADF",
			x"0000" when x"9AE0",
			x"0000" when x"9AE1",
			x"0000" when x"9AE2",
			x"0000" when x"9AE3",
			x"0000" when x"9AE4",
			x"0000" when x"9AE5",
			x"0000" when x"9AE6",
			x"0000" when x"9AE7",
			x"0000" when x"9AE8",
			x"0000" when x"9AE9",
			x"0000" when x"9AEA",
			x"0000" when x"9AEB",
			x"0000" when x"9AEC",
			x"0000" when x"9AED",
			x"0000" when x"9AEE",
			x"0000" when x"9AEF",
			x"0000" when x"9AF0",
			x"0000" when x"9AF1",
			x"0000" when x"9AF2",
			x"0000" when x"9AF3",
			x"0000" when x"9AF4",
			x"0000" when x"9AF5",
			x"0000" when x"9AF6",
			x"0000" when x"9AF7",
			x"0000" when x"9AF8",
			x"0000" when x"9AF9",
			x"0000" when x"9AFA",
			x"0000" when x"9AFB",
			x"0000" when x"9AFC",
			x"0000" when x"9AFD",
			x"0000" when x"9AFE",
			x"0000" when x"9AFF",
			x"0000" when x"9B00",
			x"0000" when x"9B01",
			x"0000" when x"9B02",
			x"0000" when x"9B03",
			x"0000" when x"9B04",
			x"0000" when x"9B05",
			x"0000" when x"9B06",
			x"0000" when x"9B07",
			x"0000" when x"9B08",
			x"0000" when x"9B09",
			x"0000" when x"9B0A",
			x"0000" when x"9B0B",
			x"0000" when x"9B0C",
			x"0000" when x"9B0D",
			x"0000" when x"9B0E",
			x"0000" when x"9B0F",
			x"0000" when x"9B10",
			x"0000" when x"9B11",
			x"0000" when x"9B12",
			x"0000" when x"9B13",
			x"0000" when x"9B14",
			x"0000" when x"9B15",
			x"0000" when x"9B16",
			x"0000" when x"9B17",
			x"0000" when x"9B18",
			x"0000" when x"9B19",
			x"0000" when x"9B1A",
			x"0000" when x"9B1B",
			x"0000" when x"9B1C",
			x"0000" when x"9B1D",
			x"0000" when x"9B1E",
			x"0000" when x"9B1F",
			x"0000" when x"9B20",
			x"0000" when x"9B21",
			x"0000" when x"9B22",
			x"0000" when x"9B23",
			x"0000" when x"9B24",
			x"0000" when x"9B25",
			x"0000" when x"9B26",
			x"0000" when x"9B27",
			x"0000" when x"9B28",
			x"0000" when x"9B29",
			x"0000" when x"9B2A",
			x"0000" when x"9B2B",
			x"0000" when x"9B2C",
			x"0000" when x"9B2D",
			x"0000" when x"9B2E",
			x"0000" when x"9B2F",
			x"0000" when x"9B30",
			x"0000" when x"9B31",
			x"0000" when x"9B32",
			x"0000" when x"9B33",
			x"0000" when x"9B34",
			x"0000" when x"9B35",
			x"0000" when x"9B36",
			x"0000" when x"9B37",
			x"0000" when x"9B38",
			x"0000" when x"9B39",
			x"0000" when x"9B3A",
			x"0000" when x"9B3B",
			x"0000" when x"9B3C",
			x"0000" when x"9B3D",
			x"0000" when x"9B3E",
			x"0000" when x"9B3F",
			x"0000" when x"9B40",
			x"0000" when x"9B41",
			x"0000" when x"9B42",
			x"0000" when x"9B43",
			x"0000" when x"9B44",
			x"0000" when x"9B45",
			x"0000" when x"9B46",
			x"0000" when x"9B47",
			x"0000" when x"9B48",
			x"0000" when x"9B49",
			x"0000" when x"9B4A",
			x"0000" when x"9B4B",
			x"0000" when x"9B4C",
			x"0000" when x"9B4D",
			x"0000" when x"9B4E",
			x"0000" when x"9B4F",
			x"0000" when x"9B50",
			x"0000" when x"9B51",
			x"0000" when x"9B52",
			x"0000" when x"9B53",
			x"0000" when x"9B54",
			x"0000" when x"9B55",
			x"0000" when x"9B56",
			x"0000" when x"9B57",
			x"0000" when x"9B58",
			x"0000" when x"9B59",
			x"0000" when x"9B5A",
			x"0000" when x"9B5B",
			x"0000" when x"9B5C",
			x"0000" when x"9B5D",
			x"0000" when x"9B5E",
			x"0000" when x"9B5F",
			x"0000" when x"9B60",
			x"0000" when x"9B61",
			x"0000" when x"9B62",
			x"0000" when x"9B63",
			x"0000" when x"9B64",
			x"0000" when x"9B65",
			x"0000" when x"9B66",
			x"0000" when x"9B67",
			x"0000" when x"9B68",
			x"0000" when x"9B69",
			x"0000" when x"9B6A",
			x"0000" when x"9B6B",
			x"0000" when x"9B6C",
			x"0000" when x"9B6D",
			x"0000" when x"9B6E",
			x"0000" when x"9B6F",
			x"0000" when x"9B70",
			x"0000" when x"9B71",
			x"0000" when x"9B72",
			x"0000" when x"9B73",
			x"0000" when x"9B74",
			x"0000" when x"9B75",
			x"0000" when x"9B76",
			x"0000" when x"9B77",
			x"0000" when x"9B78",
			x"0000" when x"9B79",
			x"0000" when x"9B7A",
			x"0000" when x"9B7B",
			x"0000" when x"9B7C",
			x"0000" when x"9B7D",
			x"0000" when x"9B7E",
			x"0000" when x"9B7F",
			x"0000" when x"9B80",
			x"0000" when x"9B81",
			x"0000" when x"9B82",
			x"0000" when x"9B83",
			x"0000" when x"9B84",
			x"0000" when x"9B85",
			x"0000" when x"9B86",
			x"0000" when x"9B87",
			x"0000" when x"9B88",
			x"0000" when x"9B89",
			x"0000" when x"9B8A",
			x"0000" when x"9B8B",
			x"0000" when x"9B8C",
			x"0000" when x"9B8D",
			x"0000" when x"9B8E",
			x"0000" when x"9B8F",
			x"0000" when x"9B90",
			x"0000" when x"9B91",
			x"0000" when x"9B92",
			x"0000" when x"9B93",
			x"0000" when x"9B94",
			x"0000" when x"9B95",
			x"0000" when x"9B96",
			x"0000" when x"9B97",
			x"0000" when x"9B98",
			x"0000" when x"9B99",
			x"0000" when x"9B9A",
			x"0000" when x"9B9B",
			x"0000" when x"9B9C",
			x"0000" when x"9B9D",
			x"0000" when x"9B9E",
			x"0000" when x"9B9F",
			x"0000" when x"9BA0",
			x"0000" when x"9BA1",
			x"0000" when x"9BA2",
			x"0000" when x"9BA3",
			x"0000" when x"9BA4",
			x"0000" when x"9BA5",
			x"0000" when x"9BA6",
			x"0000" when x"9BA7",
			x"0000" when x"9BA8",
			x"0000" when x"9BA9",
			x"0000" when x"9BAA",
			x"0000" when x"9BAB",
			x"0000" when x"9BAC",
			x"0000" when x"9BAD",
			x"0000" when x"9BAE",
			x"0000" when x"9BAF",
			x"0000" when x"9BB0",
			x"0000" when x"9BB1",
			x"0000" when x"9BB2",
			x"0000" when x"9BB3",
			x"0000" when x"9BB4",
			x"0000" when x"9BB5",
			x"0000" when x"9BB6",
			x"0000" when x"9BB7",
			x"0000" when x"9BB8",
			x"0000" when x"9BB9",
			x"0000" when x"9BBA",
			x"0000" when x"9BBB",
			x"0000" when x"9BBC",
			x"0000" when x"9BBD",
			x"0000" when x"9BBE",
			x"0000" when x"9BBF",
			x"0000" when x"9BC0",
			x"0000" when x"9BC1",
			x"0000" when x"9BC2",
			x"0000" when x"9BC3",
			x"0000" when x"9BC4",
			x"0000" when x"9BC5",
			x"0000" when x"9BC6",
			x"0000" when x"9BC7",
			x"0000" when x"9BC8",
			x"0000" when x"9BC9",
			x"0000" when x"9BCA",
			x"0000" when x"9BCB",
			x"0000" when x"9BCC",
			x"0000" when x"9BCD",
			x"0000" when x"9BCE",
			x"0000" when x"9BCF",
			x"0000" when x"9BD0",
			x"0000" when x"9BD1",
			x"0000" when x"9BD2",
			x"0000" when x"9BD3",
			x"0000" when x"9BD4",
			x"0000" when x"9BD5",
			x"0000" when x"9BD6",
			x"0000" when x"9BD7",
			x"0000" when x"9BD8",
			x"0000" when x"9BD9",
			x"0000" when x"9BDA",
			x"0000" when x"9BDB",
			x"0000" when x"9BDC",
			x"0000" when x"9BDD",
			x"0000" when x"9BDE",
			x"0000" when x"9BDF",
			x"0000" when x"9BE0",
			x"0000" when x"9BE1",
			x"0000" when x"9BE2",
			x"0000" when x"9BE3",
			x"0000" when x"9BE4",
			x"0000" when x"9BE5",
			x"0000" when x"9BE6",
			x"0000" when x"9BE7",
			x"0000" when x"9BE8",
			x"0000" when x"9BE9",
			x"0000" when x"9BEA",
			x"0000" when x"9BEB",
			x"0000" when x"9BEC",
			x"0000" when x"9BED",
			x"0000" when x"9BEE",
			x"0000" when x"9BEF",
			x"0000" when x"9BF0",
			x"0000" when x"9BF1",
			x"0000" when x"9BF2",
			x"0000" when x"9BF3",
			x"0000" when x"9BF4",
			x"0000" when x"9BF5",
			x"0000" when x"9BF6",
			x"0000" when x"9BF7",
			x"0000" when x"9BF8",
			x"0000" when x"9BF9",
			x"0000" when x"9BFA",
			x"0000" when x"9BFB",
			x"0000" when x"9BFC",
			x"0000" when x"9BFD",
			x"0000" when x"9BFE",
			x"0000" when x"9BFF",
			x"0000" when x"9C00",
			x"0000" when x"9C01",
			x"0000" when x"9C02",
			x"0000" when x"9C03",
			x"0000" when x"9C04",
			x"0000" when x"9C05",
			x"0000" when x"9C06",
			x"0000" when x"9C07",
			x"0000" when x"9C08",
			x"0000" when x"9C09",
			x"0000" when x"9C0A",
			x"0000" when x"9C0B",
			x"0000" when x"9C0C",
			x"0000" when x"9C0D",
			x"0000" when x"9C0E",
			x"0000" when x"9C0F",
			x"0000" when x"9C10",
			x"0000" when x"9C11",
			x"0000" when x"9C12",
			x"0000" when x"9C13",
			x"0000" when x"9C14",
			x"0000" when x"9C15",
			x"0000" when x"9C16",
			x"0000" when x"9C17",
			x"0000" when x"9C18",
			x"0000" when x"9C19",
			x"0000" when x"9C1A",
			x"0000" when x"9C1B",
			x"0000" when x"9C1C",
			x"0000" when x"9C1D",
			x"0000" when x"9C1E",
			x"0000" when x"9C1F",
			x"0000" when x"9C20",
			x"0000" when x"9C21",
			x"0000" when x"9C22",
			x"0000" when x"9C23",
			x"0000" when x"9C24",
			x"0000" when x"9C25",
			x"0000" when x"9C26",
			x"0000" when x"9C27",
			x"0000" when x"9C28",
			x"0000" when x"9C29",
			x"0000" when x"9C2A",
			x"0000" when x"9C2B",
			x"0000" when x"9C2C",
			x"0000" when x"9C2D",
			x"0000" when x"9C2E",
			x"0000" when x"9C2F",
			x"0000" when x"9C30",
			x"0000" when x"9C31",
			x"0000" when x"9C32",
			x"0000" when x"9C33",
			x"0000" when x"9C34",
			x"0000" when x"9C35",
			x"0000" when x"9C36",
			x"0000" when x"9C37",
			x"0000" when x"9C38",
			x"0000" when x"9C39",
			x"0000" when x"9C3A",
			x"0000" when x"9C3B",
			x"0000" when x"9C3C",
			x"0000" when x"9C3D",
			x"0000" when x"9C3E",
			x"0000" when x"9C3F",
			x"0000" when x"9C40",
			x"0000" when x"9C41",
			x"0000" when x"9C42",
			x"0000" when x"9C43",
			x"0000" when x"9C44",
			x"0000" when x"9C45",
			x"0000" when x"9C46",
			x"0000" when x"9C47",
			x"0000" when x"9C48",
			x"0000" when x"9C49",
			x"0000" when x"9C4A",
			x"0000" when x"9C4B",
			x"0000" when x"9C4C",
			x"0000" when x"9C4D",
			x"0000" when x"9C4E",
			x"0000" when x"9C4F",
			x"0000" when x"9C50",
			x"0000" when x"9C51",
			x"0000" when x"9C52",
			x"0000" when x"9C53",
			x"0000" when x"9C54",
			x"0000" when x"9C55",
			x"0000" when x"9C56",
			x"0000" when x"9C57",
			x"0000" when x"9C58",
			x"0000" when x"9C59",
			x"0000" when x"9C5A",
			x"0000" when x"9C5B",
			x"0000" when x"9C5C",
			x"0000" when x"9C5D",
			x"0000" when x"9C5E",
			x"0000" when x"9C5F",
			x"0000" when x"9C60",
			x"0000" when x"9C61",
			x"0000" when x"9C62",
			x"0000" when x"9C63",
			x"0000" when x"9C64",
			x"0000" when x"9C65",
			x"0000" when x"9C66",
			x"0000" when x"9C67",
			x"0000" when x"9C68",
			x"0000" when x"9C69",
			x"0000" when x"9C6A",
			x"0000" when x"9C6B",
			x"0000" when x"9C6C",
			x"0000" when x"9C6D",
			x"0000" when x"9C6E",
			x"0000" when x"9C6F",
			x"0000" when x"9C70",
			x"0000" when x"9C71",
			x"0000" when x"9C72",
			x"0000" when x"9C73",
			x"0000" when x"9C74",
			x"0000" when x"9C75",
			x"0000" when x"9C76",
			x"0000" when x"9C77",
			x"0000" when x"9C78",
			x"0000" when x"9C79",
			x"0000" when x"9C7A",
			x"0000" when x"9C7B",
			x"0000" when x"9C7C",
			x"0000" when x"9C7D",
			x"0000" when x"9C7E",
			x"0000" when x"9C7F",
			x"0000" when x"9C80",
			x"0000" when x"9C81",
			x"0000" when x"9C82",
			x"0000" when x"9C83",
			x"0000" when x"9C84",
			x"0000" when x"9C85",
			x"0000" when x"9C86",
			x"0000" when x"9C87",
			x"0000" when x"9C88",
			x"0000" when x"9C89",
			x"0000" when x"9C8A",
			x"0000" when x"9C8B",
			x"0000" when x"9C8C",
			x"0000" when x"9C8D",
			x"0000" when x"9C8E",
			x"0000" when x"9C8F",
			x"0000" when x"9C90",
			x"0000" when x"9C91",
			x"0000" when x"9C92",
			x"0000" when x"9C93",
			x"0000" when x"9C94",
			x"0000" when x"9C95",
			x"0000" when x"9C96",
			x"0000" when x"9C97",
			x"0000" when x"9C98",
			x"0000" when x"9C99",
			x"0000" when x"9C9A",
			x"0000" when x"9C9B",
			x"0000" when x"9C9C",
			x"0000" when x"9C9D",
			x"0000" when x"9C9E",
			x"0000" when x"9C9F",
			x"0000" when x"9CA0",
			x"0000" when x"9CA1",
			x"0000" when x"9CA2",
			x"0000" when x"9CA3",
			x"0000" when x"9CA4",
			x"0000" when x"9CA5",
			x"0000" when x"9CA6",
			x"0000" when x"9CA7",
			x"0000" when x"9CA8",
			x"0000" when x"9CA9",
			x"0000" when x"9CAA",
			x"0000" when x"9CAB",
			x"0000" when x"9CAC",
			x"0000" when x"9CAD",
			x"0000" when x"9CAE",
			x"0000" when x"9CAF",
			x"0000" when x"9CB0",
			x"0000" when x"9CB1",
			x"0000" when x"9CB2",
			x"0000" when x"9CB3",
			x"0000" when x"9CB4",
			x"0000" when x"9CB5",
			x"0000" when x"9CB6",
			x"0000" when x"9CB7",
			x"0000" when x"9CB8",
			x"0000" when x"9CB9",
			x"0000" when x"9CBA",
			x"0000" when x"9CBB",
			x"0000" when x"9CBC",
			x"0000" when x"9CBD",
			x"0000" when x"9CBE",
			x"0000" when x"9CBF",
			x"0000" when x"9CC0",
			x"0000" when x"9CC1",
			x"0000" when x"9CC2",
			x"0000" when x"9CC3",
			x"0000" when x"9CC4",
			x"0000" when x"9CC5",
			x"0000" when x"9CC6",
			x"0000" when x"9CC7",
			x"0000" when x"9CC8",
			x"0000" when x"9CC9",
			x"0000" when x"9CCA",
			x"0000" when x"9CCB",
			x"0000" when x"9CCC",
			x"0000" when x"9CCD",
			x"0000" when x"9CCE",
			x"0000" when x"9CCF",
			x"0000" when x"9CD0",
			x"0000" when x"9CD1",
			x"0000" when x"9CD2",
			x"0000" when x"9CD3",
			x"0000" when x"9CD4",
			x"0000" when x"9CD5",
			x"0000" when x"9CD6",
			x"0000" when x"9CD7",
			x"0000" when x"9CD8",
			x"0000" when x"9CD9",
			x"0000" when x"9CDA",
			x"0000" when x"9CDB",
			x"0000" when x"9CDC",
			x"0000" when x"9CDD",
			x"0000" when x"9CDE",
			x"0000" when x"9CDF",
			x"0000" when x"9CE0",
			x"0000" when x"9CE1",
			x"0000" when x"9CE2",
			x"0000" when x"9CE3",
			x"0000" when x"9CE4",
			x"0000" when x"9CE5",
			x"0000" when x"9CE6",
			x"0000" when x"9CE7",
			x"0000" when x"9CE8",
			x"0000" when x"9CE9",
			x"0000" when x"9CEA",
			x"0000" when x"9CEB",
			x"0000" when x"9CEC",
			x"0000" when x"9CED",
			x"0000" when x"9CEE",
			x"0000" when x"9CEF",
			x"0000" when x"9CF0",
			x"0000" when x"9CF1",
			x"0000" when x"9CF2",
			x"0000" when x"9CF3",
			x"0000" when x"9CF4",
			x"0000" when x"9CF5",
			x"0000" when x"9CF6",
			x"0000" when x"9CF7",
			x"0000" when x"9CF8",
			x"0000" when x"9CF9",
			x"0000" when x"9CFA",
			x"0000" when x"9CFB",
			x"0000" when x"9CFC",
			x"0000" when x"9CFD",
			x"0000" when x"9CFE",
			x"0000" when x"9CFF",
			x"0000" when x"9D00",
			x"0000" when x"9D01",
			x"0000" when x"9D02",
			x"0000" when x"9D03",
			x"0000" when x"9D04",
			x"0000" when x"9D05",
			x"0000" when x"9D06",
			x"0000" when x"9D07",
			x"0000" when x"9D08",
			x"0000" when x"9D09",
			x"0000" when x"9D0A",
			x"0000" when x"9D0B",
			x"0000" when x"9D0C",
			x"0000" when x"9D0D",
			x"0000" when x"9D0E",
			x"0000" when x"9D0F",
			x"0000" when x"9D10",
			x"0000" when x"9D11",
			x"0000" when x"9D12",
			x"0000" when x"9D13",
			x"0000" when x"9D14",
			x"0000" when x"9D15",
			x"0000" when x"9D16",
			x"0000" when x"9D17",
			x"0000" when x"9D18",
			x"0000" when x"9D19",
			x"0000" when x"9D1A",
			x"0000" when x"9D1B",
			x"0000" when x"9D1C",
			x"0000" when x"9D1D",
			x"0000" when x"9D1E",
			x"0000" when x"9D1F",
			x"0000" when x"9D20",
			x"0000" when x"9D21",
			x"0000" when x"9D22",
			x"0000" when x"9D23",
			x"0000" when x"9D24",
			x"0000" when x"9D25",
			x"0000" when x"9D26",
			x"0000" when x"9D27",
			x"0000" when x"9D28",
			x"0000" when x"9D29",
			x"0000" when x"9D2A",
			x"0000" when x"9D2B",
			x"0000" when x"9D2C",
			x"0000" when x"9D2D",
			x"0000" when x"9D2E",
			x"0000" when x"9D2F",
			x"0000" when x"9D30",
			x"0000" when x"9D31",
			x"0000" when x"9D32",
			x"0000" when x"9D33",
			x"0000" when x"9D34",
			x"0000" when x"9D35",
			x"0000" when x"9D36",
			x"0000" when x"9D37",
			x"0000" when x"9D38",
			x"0000" when x"9D39",
			x"0000" when x"9D3A",
			x"0000" when x"9D3B",
			x"0000" when x"9D3C",
			x"0000" when x"9D3D",
			x"0000" when x"9D3E",
			x"0000" when x"9D3F",
			x"0000" when x"9D40",
			x"0000" when x"9D41",
			x"0000" when x"9D42",
			x"0000" when x"9D43",
			x"0000" when x"9D44",
			x"0000" when x"9D45",
			x"0000" when x"9D46",
			x"0000" when x"9D47",
			x"0000" when x"9D48",
			x"0000" when x"9D49",
			x"0000" when x"9D4A",
			x"0000" when x"9D4B",
			x"0000" when x"9D4C",
			x"0000" when x"9D4D",
			x"0000" when x"9D4E",
			x"0000" when x"9D4F",
			x"0000" when x"9D50",
			x"0000" when x"9D51",
			x"0000" when x"9D52",
			x"0000" when x"9D53",
			x"0000" when x"9D54",
			x"0000" when x"9D55",
			x"0000" when x"9D56",
			x"0000" when x"9D57",
			x"0000" when x"9D58",
			x"0000" when x"9D59",
			x"0000" when x"9D5A",
			x"0000" when x"9D5B",
			x"0000" when x"9D5C",
			x"0000" when x"9D5D",
			x"0000" when x"9D5E",
			x"0000" when x"9D5F",
			x"0000" when x"9D60",
			x"0000" when x"9D61",
			x"0000" when x"9D62",
			x"0000" when x"9D63",
			x"0000" when x"9D64",
			x"0000" when x"9D65",
			x"0000" when x"9D66",
			x"0000" when x"9D67",
			x"0000" when x"9D68",
			x"0000" when x"9D69",
			x"0000" when x"9D6A",
			x"0000" when x"9D6B",
			x"0000" when x"9D6C",
			x"0000" when x"9D6D",
			x"0000" when x"9D6E",
			x"0000" when x"9D6F",
			x"0000" when x"9D70",
			x"0000" when x"9D71",
			x"0000" when x"9D72",
			x"0000" when x"9D73",
			x"0000" when x"9D74",
			x"0000" when x"9D75",
			x"0000" when x"9D76",
			x"0000" when x"9D77",
			x"0000" when x"9D78",
			x"0000" when x"9D79",
			x"0000" when x"9D7A",
			x"0000" when x"9D7B",
			x"0000" when x"9D7C",
			x"0000" when x"9D7D",
			x"0000" when x"9D7E",
			x"0000" when x"9D7F",
			x"0000" when x"9D80",
			x"0000" when x"9D81",
			x"0000" when x"9D82",
			x"0000" when x"9D83",
			x"0000" when x"9D84",
			x"0000" when x"9D85",
			x"0000" when x"9D86",
			x"0000" when x"9D87",
			x"0000" when x"9D88",
			x"0000" when x"9D89",
			x"0000" when x"9D8A",
			x"0000" when x"9D8B",
			x"0000" when x"9D8C",
			x"0000" when x"9D8D",
			x"0000" when x"9D8E",
			x"0000" when x"9D8F",
			x"0000" when x"9D90",
			x"0000" when x"9D91",
			x"0000" when x"9D92",
			x"0000" when x"9D93",
			x"0000" when x"9D94",
			x"0000" when x"9D95",
			x"0000" when x"9D96",
			x"0000" when x"9D97",
			x"0000" when x"9D98",
			x"0000" when x"9D99",
			x"0000" when x"9D9A",
			x"0000" when x"9D9B",
			x"0000" when x"9D9C",
			x"0000" when x"9D9D",
			x"0000" when x"9D9E",
			x"0000" when x"9D9F",
			x"0000" when x"9DA0",
			x"0000" when x"9DA1",
			x"0000" when x"9DA2",
			x"0000" when x"9DA3",
			x"0000" when x"9DA4",
			x"0000" when x"9DA5",
			x"0000" when x"9DA6",
			x"0000" when x"9DA7",
			x"0000" when x"9DA8",
			x"0000" when x"9DA9",
			x"0000" when x"9DAA",
			x"0000" when x"9DAB",
			x"0000" when x"9DAC",
			x"0000" when x"9DAD",
			x"0000" when x"9DAE",
			x"0000" when x"9DAF",
			x"0000" when x"9DB0",
			x"0000" when x"9DB1",
			x"0000" when x"9DB2",
			x"0000" when x"9DB3",
			x"0000" when x"9DB4",
			x"0000" when x"9DB5",
			x"0000" when x"9DB6",
			x"0000" when x"9DB7",
			x"0000" when x"9DB8",
			x"0000" when x"9DB9",
			x"0000" when x"9DBA",
			x"0000" when x"9DBB",
			x"0000" when x"9DBC",
			x"0000" when x"9DBD",
			x"0000" when x"9DBE",
			x"0000" when x"9DBF",
			x"0000" when x"9DC0",
			x"0000" when x"9DC1",
			x"0000" when x"9DC2",
			x"0000" when x"9DC3",
			x"0000" when x"9DC4",
			x"0000" when x"9DC5",
			x"0000" when x"9DC6",
			x"0000" when x"9DC7",
			x"0000" when x"9DC8",
			x"0000" when x"9DC9",
			x"0000" when x"9DCA",
			x"0000" when x"9DCB",
			x"0000" when x"9DCC",
			x"0000" when x"9DCD",
			x"0000" when x"9DCE",
			x"0000" when x"9DCF",
			x"0000" when x"9DD0",
			x"0000" when x"9DD1",
			x"0000" when x"9DD2",
			x"0000" when x"9DD3",
			x"0000" when x"9DD4",
			x"0000" when x"9DD5",
			x"0000" when x"9DD6",
			x"0000" when x"9DD7",
			x"0000" when x"9DD8",
			x"0000" when x"9DD9",
			x"0000" when x"9DDA",
			x"0000" when x"9DDB",
			x"0000" when x"9DDC",
			x"0000" when x"9DDD",
			x"0000" when x"9DDE",
			x"0000" when x"9DDF",
			x"0000" when x"9DE0",
			x"0000" when x"9DE1",
			x"0000" when x"9DE2",
			x"0000" when x"9DE3",
			x"0000" when x"9DE4",
			x"0000" when x"9DE5",
			x"0000" when x"9DE6",
			x"0000" when x"9DE7",
			x"0000" when x"9DE8",
			x"0000" when x"9DE9",
			x"0000" when x"9DEA",
			x"0000" when x"9DEB",
			x"0000" when x"9DEC",
			x"0000" when x"9DED",
			x"0000" when x"9DEE",
			x"0000" when x"9DEF",
			x"0000" when x"9DF0",
			x"0000" when x"9DF1",
			x"0000" when x"9DF2",
			x"0000" when x"9DF3",
			x"0000" when x"9DF4",
			x"0000" when x"9DF5",
			x"0000" when x"9DF6",
			x"0000" when x"9DF7",
			x"0000" when x"9DF8",
			x"0000" when x"9DF9",
			x"0000" when x"9DFA",
			x"0000" when x"9DFB",
			x"0000" when x"9DFC",
			x"0000" when x"9DFD",
			x"0000" when x"9DFE",
			x"0000" when x"9DFF",
			x"0000" when x"9E00",
			x"0000" when x"9E01",
			x"0000" when x"9E02",
			x"0000" when x"9E03",
			x"0000" when x"9E04",
			x"0000" when x"9E05",
			x"0000" when x"9E06",
			x"0000" when x"9E07",
			x"0000" when x"9E08",
			x"0000" when x"9E09",
			x"0000" when x"9E0A",
			x"0000" when x"9E0B",
			x"0000" when x"9E0C",
			x"0000" when x"9E0D",
			x"0000" when x"9E0E",
			x"0000" when x"9E0F",
			x"0000" when x"9E10",
			x"0000" when x"9E11",
			x"0000" when x"9E12",
			x"0000" when x"9E13",
			x"0000" when x"9E14",
			x"0000" when x"9E15",
			x"0000" when x"9E16",
			x"0000" when x"9E17",
			x"0000" when x"9E18",
			x"0000" when x"9E19",
			x"0000" when x"9E1A",
			x"0000" when x"9E1B",
			x"0000" when x"9E1C",
			x"0000" when x"9E1D",
			x"0000" when x"9E1E",
			x"0000" when x"9E1F",
			x"0000" when x"9E20",
			x"0000" when x"9E21",
			x"0000" when x"9E22",
			x"0000" when x"9E23",
			x"0000" when x"9E24",
			x"0000" when x"9E25",
			x"0000" when x"9E26",
			x"0000" when x"9E27",
			x"0000" when x"9E28",
			x"0000" when x"9E29",
			x"0000" when x"9E2A",
			x"0000" when x"9E2B",
			x"0000" when x"9E2C",
			x"0000" when x"9E2D",
			x"0000" when x"9E2E",
			x"0000" when x"9E2F",
			x"0000" when x"9E30",
			x"0000" when x"9E31",
			x"0000" when x"9E32",
			x"0000" when x"9E33",
			x"0000" when x"9E34",
			x"0000" when x"9E35",
			x"0000" when x"9E36",
			x"0000" when x"9E37",
			x"0000" when x"9E38",
			x"0000" when x"9E39",
			x"0000" when x"9E3A",
			x"0000" when x"9E3B",
			x"0000" when x"9E3C",
			x"0000" when x"9E3D",
			x"0000" when x"9E3E",
			x"0000" when x"9E3F",
			x"0000" when x"9E40",
			x"0000" when x"9E41",
			x"0000" when x"9E42",
			x"0000" when x"9E43",
			x"0000" when x"9E44",
			x"0000" when x"9E45",
			x"0000" when x"9E46",
			x"0000" when x"9E47",
			x"0000" when x"9E48",
			x"0000" when x"9E49",
			x"0000" when x"9E4A",
			x"0000" when x"9E4B",
			x"0000" when x"9E4C",
			x"0000" when x"9E4D",
			x"0000" when x"9E4E",
			x"0000" when x"9E4F",
			x"0000" when x"9E50",
			x"0000" when x"9E51",
			x"0000" when x"9E52",
			x"0000" when x"9E53",
			x"0000" when x"9E54",
			x"0000" when x"9E55",
			x"0000" when x"9E56",
			x"0000" when x"9E57",
			x"0000" when x"9E58",
			x"0000" when x"9E59",
			x"0000" when x"9E5A",
			x"0000" when x"9E5B",
			x"0000" when x"9E5C",
			x"0000" when x"9E5D",
			x"0000" when x"9E5E",
			x"0000" when x"9E5F",
			x"0000" when x"9E60",
			x"0000" when x"9E61",
			x"0000" when x"9E62",
			x"0000" when x"9E63",
			x"0000" when x"9E64",
			x"0000" when x"9E65",
			x"0000" when x"9E66",
			x"0000" when x"9E67",
			x"0000" when x"9E68",
			x"0000" when x"9E69",
			x"0000" when x"9E6A",
			x"0000" when x"9E6B",
			x"0000" when x"9E6C",
			x"0000" when x"9E6D",
			x"0000" when x"9E6E",
			x"0000" when x"9E6F",
			x"0000" when x"9E70",
			x"0000" when x"9E71",
			x"0000" when x"9E72",
			x"0000" when x"9E73",
			x"0000" when x"9E74",
			x"0000" when x"9E75",
			x"0000" when x"9E76",
			x"0000" when x"9E77",
			x"0000" when x"9E78",
			x"0000" when x"9E79",
			x"0000" when x"9E7A",
			x"0000" when x"9E7B",
			x"0000" when x"9E7C",
			x"0000" when x"9E7D",
			x"0000" when x"9E7E",
			x"0000" when x"9E7F",
			x"0000" when x"9E80",
			x"0000" when x"9E81",
			x"0000" when x"9E82",
			x"0000" when x"9E83",
			x"0000" when x"9E84",
			x"0000" when x"9E85",
			x"0000" when x"9E86",
			x"0000" when x"9E87",
			x"0000" when x"9E88",
			x"0000" when x"9E89",
			x"0000" when x"9E8A",
			x"0000" when x"9E8B",
			x"0000" when x"9E8C",
			x"0000" when x"9E8D",
			x"0000" when x"9E8E",
			x"0000" when x"9E8F",
			x"0000" when x"9E90",
			x"0000" when x"9E91",
			x"0000" when x"9E92",
			x"0000" when x"9E93",
			x"0000" when x"9E94",
			x"0000" when x"9E95",
			x"0000" when x"9E96",
			x"0000" when x"9E97",
			x"0000" when x"9E98",
			x"0000" when x"9E99",
			x"0000" when x"9E9A",
			x"0000" when x"9E9B",
			x"0000" when x"9E9C",
			x"0000" when x"9E9D",
			x"0000" when x"9E9E",
			x"0000" when x"9E9F",
			x"0000" when x"9EA0",
			x"0000" when x"9EA1",
			x"0000" when x"9EA2",
			x"0000" when x"9EA3",
			x"0000" when x"9EA4",
			x"0000" when x"9EA5",
			x"0000" when x"9EA6",
			x"0000" when x"9EA7",
			x"0000" when x"9EA8",
			x"0000" when x"9EA9",
			x"0000" when x"9EAA",
			x"0000" when x"9EAB",
			x"0000" when x"9EAC",
			x"0000" when x"9EAD",
			x"0000" when x"9EAE",
			x"0000" when x"9EAF",
			x"0000" when x"9EB0",
			x"0000" when x"9EB1",
			x"0000" when x"9EB2",
			x"0000" when x"9EB3",
			x"0000" when x"9EB4",
			x"0000" when x"9EB5",
			x"0000" when x"9EB6",
			x"0000" when x"9EB7",
			x"0000" when x"9EB8",
			x"0000" when x"9EB9",
			x"0000" when x"9EBA",
			x"0000" when x"9EBB",
			x"0000" when x"9EBC",
			x"0000" when x"9EBD",
			x"0000" when x"9EBE",
			x"0000" when x"9EBF",
			x"0000" when x"9EC0",
			x"0000" when x"9EC1",
			x"0000" when x"9EC2",
			x"0000" when x"9EC3",
			x"0000" when x"9EC4",
			x"0000" when x"9EC5",
			x"0000" when x"9EC6",
			x"0000" when x"9EC7",
			x"0000" when x"9EC8",
			x"0000" when x"9EC9",
			x"0000" when x"9ECA",
			x"0000" when x"9ECB",
			x"0000" when x"9ECC",
			x"0000" when x"9ECD",
			x"0000" when x"9ECE",
			x"0000" when x"9ECF",
			x"0000" when x"9ED0",
			x"0000" when x"9ED1",
			x"0000" when x"9ED2",
			x"0000" when x"9ED3",
			x"0000" when x"9ED4",
			x"0000" when x"9ED5",
			x"0000" when x"9ED6",
			x"0000" when x"9ED7",
			x"0000" when x"9ED8",
			x"0000" when x"9ED9",
			x"0000" when x"9EDA",
			x"0000" when x"9EDB",
			x"0000" when x"9EDC",
			x"0000" when x"9EDD",
			x"0000" when x"9EDE",
			x"0000" when x"9EDF",
			x"0000" when x"9EE0",
			x"0000" when x"9EE1",
			x"0000" when x"9EE2",
			x"0000" when x"9EE3",
			x"0000" when x"9EE4",
			x"0000" when x"9EE5",
			x"0000" when x"9EE6",
			x"0000" when x"9EE7",
			x"0000" when x"9EE8",
			x"0000" when x"9EE9",
			x"0000" when x"9EEA",
			x"0000" when x"9EEB",
			x"0000" when x"9EEC",
			x"0000" when x"9EED",
			x"0000" when x"9EEE",
			x"0000" when x"9EEF",
			x"0000" when x"9EF0",
			x"0000" when x"9EF1",
			x"0000" when x"9EF2",
			x"0000" when x"9EF3",
			x"0000" when x"9EF4",
			x"0000" when x"9EF5",
			x"0000" when x"9EF6",
			x"0000" when x"9EF7",
			x"0000" when x"9EF8",
			x"0000" when x"9EF9",
			x"0000" when x"9EFA",
			x"0000" when x"9EFB",
			x"0000" when x"9EFC",
			x"0000" when x"9EFD",
			x"0000" when x"9EFE",
			x"0000" when x"9EFF",
			x"0000" when x"9F00",
			x"0000" when x"9F01",
			x"0000" when x"9F02",
			x"0000" when x"9F03",
			x"0000" when x"9F04",
			x"0000" when x"9F05",
			x"0000" when x"9F06",
			x"0000" when x"9F07",
			x"0000" when x"9F08",
			x"0000" when x"9F09",
			x"0000" when x"9F0A",
			x"0000" when x"9F0B",
			x"0000" when x"9F0C",
			x"0000" when x"9F0D",
			x"0000" when x"9F0E",
			x"0000" when x"9F0F",
			x"0000" when x"9F10",
			x"0000" when x"9F11",
			x"0000" when x"9F12",
			x"0000" when x"9F13",
			x"0000" when x"9F14",
			x"0000" when x"9F15",
			x"0000" when x"9F16",
			x"0000" when x"9F17",
			x"0000" when x"9F18",
			x"0000" when x"9F19",
			x"0000" when x"9F1A",
			x"0000" when x"9F1B",
			x"0000" when x"9F1C",
			x"0000" when x"9F1D",
			x"0000" when x"9F1E",
			x"0000" when x"9F1F",
			x"0000" when x"9F20",
			x"0000" when x"9F21",
			x"0000" when x"9F22",
			x"0000" when x"9F23",
			x"0000" when x"9F24",
			x"0000" when x"9F25",
			x"0000" when x"9F26",
			x"0000" when x"9F27",
			x"0000" when x"9F28",
			x"0000" when x"9F29",
			x"0000" when x"9F2A",
			x"0000" when x"9F2B",
			x"0000" when x"9F2C",
			x"0000" when x"9F2D",
			x"0000" when x"9F2E",
			x"0000" when x"9F2F",
			x"0000" when x"9F30",
			x"0000" when x"9F31",
			x"0000" when x"9F32",
			x"0000" when x"9F33",
			x"0000" when x"9F34",
			x"0000" when x"9F35",
			x"0000" when x"9F36",
			x"0000" when x"9F37",
			x"0000" when x"9F38",
			x"0000" when x"9F39",
			x"0000" when x"9F3A",
			x"0000" when x"9F3B",
			x"0000" when x"9F3C",
			x"0000" when x"9F3D",
			x"0000" when x"9F3E",
			x"0000" when x"9F3F",
			x"0000" when x"9F40",
			x"0000" when x"9F41",
			x"0000" when x"9F42",
			x"0000" when x"9F43",
			x"0000" when x"9F44",
			x"0000" when x"9F45",
			x"0000" when x"9F46",
			x"0000" when x"9F47",
			x"0000" when x"9F48",
			x"0000" when x"9F49",
			x"0000" when x"9F4A",
			x"0000" when x"9F4B",
			x"0000" when x"9F4C",
			x"0000" when x"9F4D",
			x"0000" when x"9F4E",
			x"0000" when x"9F4F",
			x"0000" when x"9F50",
			x"0000" when x"9F51",
			x"0000" when x"9F52",
			x"0000" when x"9F53",
			x"0000" when x"9F54",
			x"0000" when x"9F55",
			x"0000" when x"9F56",
			x"0000" when x"9F57",
			x"0000" when x"9F58",
			x"0000" when x"9F59",
			x"0000" when x"9F5A",
			x"0000" when x"9F5B",
			x"0000" when x"9F5C",
			x"0000" when x"9F5D",
			x"0000" when x"9F5E",
			x"0000" when x"9F5F",
			x"0000" when x"9F60",
			x"0000" when x"9F61",
			x"0000" when x"9F62",
			x"0000" when x"9F63",
			x"0000" when x"9F64",
			x"0000" when x"9F65",
			x"0000" when x"9F66",
			x"0000" when x"9F67",
			x"0000" when x"9F68",
			x"0000" when x"9F69",
			x"0000" when x"9F6A",
			x"0000" when x"9F6B",
			x"0000" when x"9F6C",
			x"0000" when x"9F6D",
			x"0000" when x"9F6E",
			x"0000" when x"9F6F",
			x"0000" when x"9F70",
			x"0000" when x"9F71",
			x"0000" when x"9F72",
			x"0000" when x"9F73",
			x"0000" when x"9F74",
			x"0000" when x"9F75",
			x"0000" when x"9F76",
			x"0000" when x"9F77",
			x"0000" when x"9F78",
			x"0000" when x"9F79",
			x"0000" when x"9F7A",
			x"0000" when x"9F7B",
			x"0000" when x"9F7C",
			x"0000" when x"9F7D",
			x"0000" when x"9F7E",
			x"0000" when x"9F7F",
			x"0000" when x"9F80",
			x"0000" when x"9F81",
			x"0000" when x"9F82",
			x"0000" when x"9F83",
			x"0000" when x"9F84",
			x"0000" when x"9F85",
			x"0000" when x"9F86",
			x"0000" when x"9F87",
			x"0000" when x"9F88",
			x"0000" when x"9F89",
			x"0000" when x"9F8A",
			x"0000" when x"9F8B",
			x"0000" when x"9F8C",
			x"0000" when x"9F8D",
			x"0000" when x"9F8E",
			x"0000" when x"9F8F",
			x"0000" when x"9F90",
			x"0000" when x"9F91",
			x"0000" when x"9F92",
			x"0000" when x"9F93",
			x"0000" when x"9F94",
			x"0000" when x"9F95",
			x"0000" when x"9F96",
			x"0000" when x"9F97",
			x"0000" when x"9F98",
			x"0000" when x"9F99",
			x"0000" when x"9F9A",
			x"0000" when x"9F9B",
			x"0000" when x"9F9C",
			x"0000" when x"9F9D",
			x"0000" when x"9F9E",
			x"0000" when x"9F9F",
			x"0000" when x"9FA0",
			x"0000" when x"9FA1",
			x"0000" when x"9FA2",
			x"0000" when x"9FA3",
			x"0000" when x"9FA4",
			x"0000" when x"9FA5",
			x"0000" when x"9FA6",
			x"0000" when x"9FA7",
			x"0000" when x"9FA8",
			x"0000" when x"9FA9",
			x"0000" when x"9FAA",
			x"0000" when x"9FAB",
			x"0000" when x"9FAC",
			x"0000" when x"9FAD",
			x"0000" when x"9FAE",
			x"0000" when x"9FAF",
			x"0000" when x"9FB0",
			x"0000" when x"9FB1",
			x"0000" when x"9FB2",
			x"0000" when x"9FB3",
			x"0000" when x"9FB4",
			x"0000" when x"9FB5",
			x"0000" when x"9FB6",
			x"0000" when x"9FB7",
			x"0000" when x"9FB8",
			x"0000" when x"9FB9",
			x"0000" when x"9FBA",
			x"0000" when x"9FBB",
			x"0000" when x"9FBC",
			x"0000" when x"9FBD",
			x"0000" when x"9FBE",
			x"0000" when x"9FBF",
			x"0000" when x"9FC0",
			x"0000" when x"9FC1",
			x"0000" when x"9FC2",
			x"0000" when x"9FC3",
			x"0000" when x"9FC4",
			x"0000" when x"9FC5",
			x"0000" when x"9FC6",
			x"0000" when x"9FC7",
			x"0000" when x"9FC8",
			x"0000" when x"9FC9",
			x"0000" when x"9FCA",
			x"0000" when x"9FCB",
			x"0000" when x"9FCC",
			x"0000" when x"9FCD",
			x"0000" when x"9FCE",
			x"0000" when x"9FCF",
			x"0000" when x"9FD0",
			x"0000" when x"9FD1",
			x"0000" when x"9FD2",
			x"0000" when x"9FD3",
			x"0000" when x"9FD4",
			x"0000" when x"9FD5",
			x"0000" when x"9FD6",
			x"0000" when x"9FD7",
			x"0000" when x"9FD8",
			x"0000" when x"9FD9",
			x"0000" when x"9FDA",
			x"0000" when x"9FDB",
			x"0000" when x"9FDC",
			x"0000" when x"9FDD",
			x"0000" when x"9FDE",
			x"0000" when x"9FDF",
			x"0000" when x"9FE0",
			x"0000" when x"9FE1",
			x"0000" when x"9FE2",
			x"0000" when x"9FE3",
			x"0000" when x"9FE4",
			x"0000" when x"9FE5",
			x"0000" when x"9FE6",
			x"0000" when x"9FE7",
			x"0000" when x"9FE8",
			x"0000" when x"9FE9",
			x"0000" when x"9FEA",
			x"0000" when x"9FEB",
			x"0000" when x"9FEC",
			x"0000" when x"9FED",
			x"0000" when x"9FEE",
			x"0000" when x"9FEF",
			x"0000" when x"9FF0",
			x"0000" when x"9FF1",
			x"0000" when x"9FF2",
			x"0000" when x"9FF3",
			x"0000" when x"9FF4",
			x"0000" when x"9FF5",
			x"0000" when x"9FF6",
			x"0000" when x"9FF7",
			x"0000" when x"9FF8",
			x"0000" when x"9FF9",
			x"0000" when x"9FFA",
			x"0000" when x"9FFB",
			x"0000" when x"9FFC",
			x"0000" when x"9FFD",
			x"0000" when x"9FFE",
			x"0000" when x"9FFF",
			x"0000" when x"A000",
			x"0000" when x"A001",
			x"0000" when x"A002",
			x"0000" when x"A003",
			x"0000" when x"A004",
			x"0000" when x"A005",
			x"0000" when x"A006",
			x"0000" when x"A007",
			x"0000" when x"A008",
			x"0000" when x"A009",
			x"0000" when x"A00A",
			x"0000" when x"A00B",
			x"0000" when x"A00C",
			x"0000" when x"A00D",
			x"0000" when x"A00E",
			x"0000" when x"A00F",
			x"0000" when x"A010",
			x"0000" when x"A011",
			x"0000" when x"A012",
			x"0000" when x"A013",
			x"0000" when x"A014",
			x"0000" when x"A015",
			x"0000" when x"A016",
			x"0000" when x"A017",
			x"0000" when x"A018",
			x"0000" when x"A019",
			x"0000" when x"A01A",
			x"0000" when x"A01B",
			x"0000" when x"A01C",
			x"0000" when x"A01D",
			x"0000" when x"A01E",
			x"0000" when x"A01F",
			x"0000" when x"A020",
			x"0000" when x"A021",
			x"0000" when x"A022",
			x"0000" when x"A023",
			x"0000" when x"A024",
			x"0000" when x"A025",
			x"0000" when x"A026",
			x"0000" when x"A027",
			x"0000" when x"A028",
			x"0000" when x"A029",
			x"0000" when x"A02A",
			x"0000" when x"A02B",
			x"0000" when x"A02C",
			x"0000" when x"A02D",
			x"0000" when x"A02E",
			x"0000" when x"A02F",
			x"0000" when x"A030",
			x"0000" when x"A031",
			x"0000" when x"A032",
			x"0000" when x"A033",
			x"0000" when x"A034",
			x"0000" when x"A035",
			x"0000" when x"A036",
			x"0000" when x"A037",
			x"0000" when x"A038",
			x"0000" when x"A039",
			x"0000" when x"A03A",
			x"0000" when x"A03B",
			x"0000" when x"A03C",
			x"0000" when x"A03D",
			x"0000" when x"A03E",
			x"0000" when x"A03F",
			x"0000" when x"A040",
			x"0000" when x"A041",
			x"0000" when x"A042",
			x"0000" when x"A043",
			x"0000" when x"A044",
			x"0000" when x"A045",
			x"0000" when x"A046",
			x"0000" when x"A047",
			x"0000" when x"A048",
			x"0000" when x"A049",
			x"0000" when x"A04A",
			x"0000" when x"A04B",
			x"0000" when x"A04C",
			x"0000" when x"A04D",
			x"0000" when x"A04E",
			x"0000" when x"A04F",
			x"0000" when x"A050",
			x"0000" when x"A051",
			x"0000" when x"A052",
			x"0000" when x"A053",
			x"0000" when x"A054",
			x"0000" when x"A055",
			x"0000" when x"A056",
			x"0000" when x"A057",
			x"0000" when x"A058",
			x"0000" when x"A059",
			x"0000" when x"A05A",
			x"0000" when x"A05B",
			x"0000" when x"A05C",
			x"0000" when x"A05D",
			x"0000" when x"A05E",
			x"0000" when x"A05F",
			x"0000" when x"A060",
			x"0000" when x"A061",
			x"0000" when x"A062",
			x"0000" when x"A063",
			x"0000" when x"A064",
			x"0000" when x"A065",
			x"0000" when x"A066",
			x"0000" when x"A067",
			x"0000" when x"A068",
			x"0000" when x"A069",
			x"0000" when x"A06A",
			x"0000" when x"A06B",
			x"0000" when x"A06C",
			x"0000" when x"A06D",
			x"0000" when x"A06E",
			x"0000" when x"A06F",
			x"0000" when x"A070",
			x"0000" when x"A071",
			x"0000" when x"A072",
			x"0000" when x"A073",
			x"0000" when x"A074",
			x"0000" when x"A075",
			x"0000" when x"A076",
			x"0000" when x"A077",
			x"0000" when x"A078",
			x"0000" when x"A079",
			x"0000" when x"A07A",
			x"0000" when x"A07B",
			x"0000" when x"A07C",
			x"0000" when x"A07D",
			x"0000" when x"A07E",
			x"0000" when x"A07F",
			x"0000" when x"A080",
			x"0000" when x"A081",
			x"0000" when x"A082",
			x"0000" when x"A083",
			x"0000" when x"A084",
			x"0000" when x"A085",
			x"0000" when x"A086",
			x"0000" when x"A087",
			x"0000" when x"A088",
			x"0000" when x"A089",
			x"0000" when x"A08A",
			x"0000" when x"A08B",
			x"0000" when x"A08C",
			x"0000" when x"A08D",
			x"0000" when x"A08E",
			x"0000" when x"A08F",
			x"0000" when x"A090",
			x"0000" when x"A091",
			x"0000" when x"A092",
			x"0000" when x"A093",
			x"0000" when x"A094",
			x"0000" when x"A095",
			x"0000" when x"A096",
			x"0000" when x"A097",
			x"0000" when x"A098",
			x"0000" when x"A099",
			x"0000" when x"A09A",
			x"0000" when x"A09B",
			x"0000" when x"A09C",
			x"0000" when x"A09D",
			x"0000" when x"A09E",
			x"0000" when x"A09F",
			x"0000" when x"A0A0",
			x"0000" when x"A0A1",
			x"0000" when x"A0A2",
			x"0000" when x"A0A3",
			x"0000" when x"A0A4",
			x"0000" when x"A0A5",
			x"0000" when x"A0A6",
			x"0000" when x"A0A7",
			x"0000" when x"A0A8",
			x"0000" when x"A0A9",
			x"0000" when x"A0AA",
			x"0000" when x"A0AB",
			x"0000" when x"A0AC",
			x"0000" when x"A0AD",
			x"0000" when x"A0AE",
			x"0000" when x"A0AF",
			x"0000" when x"A0B0",
			x"0000" when x"A0B1",
			x"0000" when x"A0B2",
			x"0000" when x"A0B3",
			x"0000" when x"A0B4",
			x"0000" when x"A0B5",
			x"0000" when x"A0B6",
			x"0000" when x"A0B7",
			x"0000" when x"A0B8",
			x"0000" when x"A0B9",
			x"0000" when x"A0BA",
			x"0000" when x"A0BB",
			x"0000" when x"A0BC",
			x"0000" when x"A0BD",
			x"0000" when x"A0BE",
			x"0000" when x"A0BF",
			x"0000" when x"A0C0",
			x"0000" when x"A0C1",
			x"0000" when x"A0C2",
			x"0000" when x"A0C3",
			x"0000" when x"A0C4",
			x"0000" when x"A0C5",
			x"0000" when x"A0C6",
			x"0000" when x"A0C7",
			x"0000" when x"A0C8",
			x"0000" when x"A0C9",
			x"0000" when x"A0CA",
			x"0000" when x"A0CB",
			x"0000" when x"A0CC",
			x"0000" when x"A0CD",
			x"0000" when x"A0CE",
			x"0000" when x"A0CF",
			x"0000" when x"A0D0",
			x"0000" when x"A0D1",
			x"0000" when x"A0D2",
			x"0000" when x"A0D3",
			x"0000" when x"A0D4",
			x"0000" when x"A0D5",
			x"0000" when x"A0D6",
			x"0000" when x"A0D7",
			x"0000" when x"A0D8",
			x"0000" when x"A0D9",
			x"0000" when x"A0DA",
			x"0000" when x"A0DB",
			x"0000" when x"A0DC",
			x"0000" when x"A0DD",
			x"0000" when x"A0DE",
			x"0000" when x"A0DF",
			x"0000" when x"A0E0",
			x"0000" when x"A0E1",
			x"0000" when x"A0E2",
			x"0000" when x"A0E3",
			x"0000" when x"A0E4",
			x"0000" when x"A0E5",
			x"0000" when x"A0E6",
			x"0000" when x"A0E7",
			x"0000" when x"A0E8",
			x"0000" when x"A0E9",
			x"0000" when x"A0EA",
			x"0000" when x"A0EB",
			x"0000" when x"A0EC",
			x"0000" when x"A0ED",
			x"0000" when x"A0EE",
			x"0000" when x"A0EF",
			x"0000" when x"A0F0",
			x"0000" when x"A0F1",
			x"0000" when x"A0F2",
			x"0000" when x"A0F3",
			x"0000" when x"A0F4",
			x"0000" when x"A0F5",
			x"0000" when x"A0F6",
			x"0000" when x"A0F7",
			x"0000" when x"A0F8",
			x"0000" when x"A0F9",
			x"0000" when x"A0FA",
			x"0000" when x"A0FB",
			x"0000" when x"A0FC",
			x"0000" when x"A0FD",
			x"0000" when x"A0FE",
			x"0000" when x"A0FF",
			x"0000" when x"A100",
			x"0000" when x"A101",
			x"0000" when x"A102",
			x"0000" when x"A103",
			x"0000" when x"A104",
			x"0000" when x"A105",
			x"0000" when x"A106",
			x"0000" when x"A107",
			x"0000" when x"A108",
			x"0000" when x"A109",
			x"0000" when x"A10A",
			x"0000" when x"A10B",
			x"0000" when x"A10C",
			x"0000" when x"A10D",
			x"0000" when x"A10E",
			x"0000" when x"A10F",
			x"0000" when x"A110",
			x"0000" when x"A111",
			x"0000" when x"A112",
			x"0000" when x"A113",
			x"0000" when x"A114",
			x"0000" when x"A115",
			x"0000" when x"A116",
			x"0000" when x"A117",
			x"0000" when x"A118",
			x"0000" when x"A119",
			x"0000" when x"A11A",
			x"0000" when x"A11B",
			x"0000" when x"A11C",
			x"0000" when x"A11D",
			x"0000" when x"A11E",
			x"0000" when x"A11F",
			x"0000" when x"A120",
			x"0000" when x"A121",
			x"0000" when x"A122",
			x"0000" when x"A123",
			x"0000" when x"A124",
			x"0000" when x"A125",
			x"0000" when x"A126",
			x"0000" when x"A127",
			x"0000" when x"A128",
			x"0000" when x"A129",
			x"0000" when x"A12A",
			x"0000" when x"A12B",
			x"0000" when x"A12C",
			x"0000" when x"A12D",
			x"0000" when x"A12E",
			x"0000" when x"A12F",
			x"0000" when x"A130",
			x"0000" when x"A131",
			x"0000" when x"A132",
			x"0000" when x"A133",
			x"0000" when x"A134",
			x"0000" when x"A135",
			x"0000" when x"A136",
			x"0000" when x"A137",
			x"0000" when x"A138",
			x"0000" when x"A139",
			x"0000" when x"A13A",
			x"0000" when x"A13B",
			x"0000" when x"A13C",
			x"0000" when x"A13D",
			x"0000" when x"A13E",
			x"0000" when x"A13F",
			x"0000" when x"A140",
			x"0000" when x"A141",
			x"0000" when x"A142",
			x"0000" when x"A143",
			x"0000" when x"A144",
			x"0000" when x"A145",
			x"0000" when x"A146",
			x"0000" when x"A147",
			x"0000" when x"A148",
			x"0000" when x"A149",
			x"0000" when x"A14A",
			x"0000" when x"A14B",
			x"0000" when x"A14C",
			x"0000" when x"A14D",
			x"0000" when x"A14E",
			x"0000" when x"A14F",
			x"0000" when x"A150",
			x"0000" when x"A151",
			x"0000" when x"A152",
			x"0000" when x"A153",
			x"0000" when x"A154",
			x"0000" when x"A155",
			x"0000" when x"A156",
			x"0000" when x"A157",
			x"0000" when x"A158",
			x"0000" when x"A159",
			x"0000" when x"A15A",
			x"0000" when x"A15B",
			x"0000" when x"A15C",
			x"0000" when x"A15D",
			x"0000" when x"A15E",
			x"0000" when x"A15F",
			x"0000" when x"A160",
			x"0000" when x"A161",
			x"0000" when x"A162",
			x"0000" when x"A163",
			x"0000" when x"A164",
			x"0000" when x"A165",
			x"0000" when x"A166",
			x"0000" when x"A167",
			x"0000" when x"A168",
			x"0000" when x"A169",
			x"0000" when x"A16A",
			x"0000" when x"A16B",
			x"0000" when x"A16C",
			x"0000" when x"A16D",
			x"0000" when x"A16E",
			x"0000" when x"A16F",
			x"0000" when x"A170",
			x"0000" when x"A171",
			x"0000" when x"A172",
			x"0000" when x"A173",
			x"0000" when x"A174",
			x"0000" when x"A175",
			x"0000" when x"A176",
			x"0000" when x"A177",
			x"0000" when x"A178",
			x"0000" when x"A179",
			x"0000" when x"A17A",
			x"0000" when x"A17B",
			x"0000" when x"A17C",
			x"0000" when x"A17D",
			x"0000" when x"A17E",
			x"0000" when x"A17F",
			x"0000" when x"A180",
			x"0000" when x"A181",
			x"0000" when x"A182",
			x"0000" when x"A183",
			x"0000" when x"A184",
			x"0000" when x"A185",
			x"0000" when x"A186",
			x"0000" when x"A187",
			x"0000" when x"A188",
			x"0000" when x"A189",
			x"0000" when x"A18A",
			x"0000" when x"A18B",
			x"0000" when x"A18C",
			x"0000" when x"A18D",
			x"0000" when x"A18E",
			x"0000" when x"A18F",
			x"0000" when x"A190",
			x"0000" when x"A191",
			x"0000" when x"A192",
			x"0000" when x"A193",
			x"0000" when x"A194",
			x"0000" when x"A195",
			x"0000" when x"A196",
			x"0000" when x"A197",
			x"0000" when x"A198",
			x"0000" when x"A199",
			x"0000" when x"A19A",
			x"0000" when x"A19B",
			x"0000" when x"A19C",
			x"0000" when x"A19D",
			x"0000" when x"A19E",
			x"0000" when x"A19F",
			x"0000" when x"A1A0",
			x"0000" when x"A1A1",
			x"0000" when x"A1A2",
			x"0000" when x"A1A3",
			x"0000" when x"A1A4",
			x"0000" when x"A1A5",
			x"0000" when x"A1A6",
			x"0000" when x"A1A7",
			x"0000" when x"A1A8",
			x"0000" when x"A1A9",
			x"0000" when x"A1AA",
			x"0000" when x"A1AB",
			x"0000" when x"A1AC",
			x"0000" when x"A1AD",
			x"0000" when x"A1AE",
			x"0000" when x"A1AF",
			x"0000" when x"A1B0",
			x"0000" when x"A1B1",
			x"0000" when x"A1B2",
			x"0000" when x"A1B3",
			x"0000" when x"A1B4",
			x"0000" when x"A1B5",
			x"0000" when x"A1B6",
			x"0000" when x"A1B7",
			x"0000" when x"A1B8",
			x"0000" when x"A1B9",
			x"0000" when x"A1BA",
			x"0000" when x"A1BB",
			x"0000" when x"A1BC",
			x"0000" when x"A1BD",
			x"0000" when x"A1BE",
			x"0000" when x"A1BF",
			x"0000" when x"A1C0",
			x"0000" when x"A1C1",
			x"0000" when x"A1C2",
			x"0000" when x"A1C3",
			x"0000" when x"A1C4",
			x"0000" when x"A1C5",
			x"0000" when x"A1C6",
			x"0000" when x"A1C7",
			x"0000" when x"A1C8",
			x"0000" when x"A1C9",
			x"0000" when x"A1CA",
			x"0000" when x"A1CB",
			x"0000" when x"A1CC",
			x"0000" when x"A1CD",
			x"0000" when x"A1CE",
			x"0000" when x"A1CF",
			x"0000" when x"A1D0",
			x"0000" when x"A1D1",
			x"0000" when x"A1D2",
			x"0000" when x"A1D3",
			x"0000" when x"A1D4",
			x"0000" when x"A1D5",
			x"0000" when x"A1D6",
			x"0000" when x"A1D7",
			x"0000" when x"A1D8",
			x"0000" when x"A1D9",
			x"0000" when x"A1DA",
			x"0000" when x"A1DB",
			x"0000" when x"A1DC",
			x"0000" when x"A1DD",
			x"0000" when x"A1DE",
			x"0000" when x"A1DF",
			x"0000" when x"A1E0",
			x"0000" when x"A1E1",
			x"0000" when x"A1E2",
			x"0000" when x"A1E3",
			x"0000" when x"A1E4",
			x"0000" when x"A1E5",
			x"0000" when x"A1E6",
			x"0000" when x"A1E7",
			x"0000" when x"A1E8",
			x"0000" when x"A1E9",
			x"0000" when x"A1EA",
			x"0000" when x"A1EB",
			x"0000" when x"A1EC",
			x"0000" when x"A1ED",
			x"0000" when x"A1EE",
			x"0000" when x"A1EF",
			x"0000" when x"A1F0",
			x"0000" when x"A1F1",
			x"0000" when x"A1F2",
			x"0000" when x"A1F3",
			x"0000" when x"A1F4",
			x"0000" when x"A1F5",
			x"0000" when x"A1F6",
			x"0000" when x"A1F7",
			x"0000" when x"A1F8",
			x"0000" when x"A1F9",
			x"0000" when x"A1FA",
			x"0000" when x"A1FB",
			x"0000" when x"A1FC",
			x"0000" when x"A1FD",
			x"0000" when x"A1FE",
			x"0000" when x"A1FF",
			x"0000" when x"A200",
			x"0000" when x"A201",
			x"0000" when x"A202",
			x"0000" when x"A203",
			x"0000" when x"A204",
			x"0000" when x"A205",
			x"0000" when x"A206",
			x"0000" when x"A207",
			x"0000" when x"A208",
			x"0000" when x"A209",
			x"0000" when x"A20A",
			x"0000" when x"A20B",
			x"0000" when x"A20C",
			x"0000" when x"A20D",
			x"0000" when x"A20E",
			x"0000" when x"A20F",
			x"0000" when x"A210",
			x"0000" when x"A211",
			x"0000" when x"A212",
			x"0000" when x"A213",
			x"0000" when x"A214",
			x"0000" when x"A215",
			x"0000" when x"A216",
			x"0000" when x"A217",
			x"0000" when x"A218",
			x"0000" when x"A219",
			x"0000" when x"A21A",
			x"0000" when x"A21B",
			x"0000" when x"A21C",
			x"0000" when x"A21D",
			x"0000" when x"A21E",
			x"0000" when x"A21F",
			x"0000" when x"A220",
			x"0000" when x"A221",
			x"0000" when x"A222",
			x"0000" when x"A223",
			x"0000" when x"A224",
			x"0000" when x"A225",
			x"0000" when x"A226",
			x"0000" when x"A227",
			x"0000" when x"A228",
			x"0000" when x"A229",
			x"0000" when x"A22A",
			x"0000" when x"A22B",
			x"0000" when x"A22C",
			x"0000" when x"A22D",
			x"0000" when x"A22E",
			x"0000" when x"A22F",
			x"0000" when x"A230",
			x"0000" when x"A231",
			x"0000" when x"A232",
			x"0000" when x"A233",
			x"0000" when x"A234",
			x"0000" when x"A235",
			x"0000" when x"A236",
			x"0000" when x"A237",
			x"0000" when x"A238",
			x"0000" when x"A239",
			x"0000" when x"A23A",
			x"0000" when x"A23B",
			x"0000" when x"A23C",
			x"0000" when x"A23D",
			x"0000" when x"A23E",
			x"0000" when x"A23F",
			x"0000" when x"A240",
			x"0000" when x"A241",
			x"0000" when x"A242",
			x"0000" when x"A243",
			x"0000" when x"A244",
			x"0000" when x"A245",
			x"0000" when x"A246",
			x"0000" when x"A247",
			x"0000" when x"A248",
			x"0000" when x"A249",
			x"0000" when x"A24A",
			x"0000" when x"A24B",
			x"0000" when x"A24C",
			x"0000" when x"A24D",
			x"0000" when x"A24E",
			x"0000" when x"A24F",
			x"0000" when x"A250",
			x"0000" when x"A251",
			x"0000" when x"A252",
			x"0000" when x"A253",
			x"0000" when x"A254",
			x"0000" when x"A255",
			x"0000" when x"A256",
			x"0000" when x"A257",
			x"0000" when x"A258",
			x"0000" when x"A259",
			x"0000" when x"A25A",
			x"0000" when x"A25B",
			x"0000" when x"A25C",
			x"0000" when x"A25D",
			x"0000" when x"A25E",
			x"0000" when x"A25F",
			x"0000" when x"A260",
			x"0000" when x"A261",
			x"0000" when x"A262",
			x"0000" when x"A263",
			x"0000" when x"A264",
			x"0000" when x"A265",
			x"0000" when x"A266",
			x"0000" when x"A267",
			x"0000" when x"A268",
			x"0000" when x"A269",
			x"0000" when x"A26A",
			x"0000" when x"A26B",
			x"0000" when x"A26C",
			x"0000" when x"A26D",
			x"0000" when x"A26E",
			x"0000" when x"A26F",
			x"0000" when x"A270",
			x"0000" when x"A271",
			x"0000" when x"A272",
			x"0000" when x"A273",
			x"0000" when x"A274",
			x"0000" when x"A275",
			x"0000" when x"A276",
			x"0000" when x"A277",
			x"0000" when x"A278",
			x"0000" when x"A279",
			x"0000" when x"A27A",
			x"0000" when x"A27B",
			x"0000" when x"A27C",
			x"0000" when x"A27D",
			x"0000" when x"A27E",
			x"0000" when x"A27F",
			x"0000" when x"A280",
			x"0000" when x"A281",
			x"0000" when x"A282",
			x"0000" when x"A283",
			x"0000" when x"A284",
			x"0000" when x"A285",
			x"0000" when x"A286",
			x"0000" when x"A287",
			x"0000" when x"A288",
			x"0000" when x"A289",
			x"0000" when x"A28A",
			x"0000" when x"A28B",
			x"0000" when x"A28C",
			x"0000" when x"A28D",
			x"0000" when x"A28E",
			x"0000" when x"A28F",
			x"0000" when x"A290",
			x"0000" when x"A291",
			x"0000" when x"A292",
			x"0000" when x"A293",
			x"0000" when x"A294",
			x"0000" when x"A295",
			x"0000" when x"A296",
			x"0000" when x"A297",
			x"0000" when x"A298",
			x"0000" when x"A299",
			x"0000" when x"A29A",
			x"0000" when x"A29B",
			x"0000" when x"A29C",
			x"0000" when x"A29D",
			x"0000" when x"A29E",
			x"0000" when x"A29F",
			x"0000" when x"A2A0",
			x"0000" when x"A2A1",
			x"0000" when x"A2A2",
			x"0000" when x"A2A3",
			x"0000" when x"A2A4",
			x"0000" when x"A2A5",
			x"0000" when x"A2A6",
			x"0000" when x"A2A7",
			x"0000" when x"A2A8",
			x"0000" when x"A2A9",
			x"0000" when x"A2AA",
			x"0000" when x"A2AB",
			x"0000" when x"A2AC",
			x"0000" when x"A2AD",
			x"0000" when x"A2AE",
			x"0000" when x"A2AF",
			x"0000" when x"A2B0",
			x"0000" when x"A2B1",
			x"0000" when x"A2B2",
			x"0000" when x"A2B3",
			x"0000" when x"A2B4",
			x"0000" when x"A2B5",
			x"0000" when x"A2B6",
			x"0000" when x"A2B7",
			x"0000" when x"A2B8",
			x"0000" when x"A2B9",
			x"0000" when x"A2BA",
			x"0000" when x"A2BB",
			x"0000" when x"A2BC",
			x"0000" when x"A2BD",
			x"0000" when x"A2BE",
			x"0000" when x"A2BF",
			x"0000" when x"A2C0",
			x"0000" when x"A2C1",
			x"0000" when x"A2C2",
			x"0000" when x"A2C3",
			x"0000" when x"A2C4",
			x"0000" when x"A2C5",
			x"0000" when x"A2C6",
			x"0000" when x"A2C7",
			x"0000" when x"A2C8",
			x"0000" when x"A2C9",
			x"0000" when x"A2CA",
			x"0000" when x"A2CB",
			x"0000" when x"A2CC",
			x"0000" when x"A2CD",
			x"0000" when x"A2CE",
			x"0000" when x"A2CF",
			x"0000" when x"A2D0",
			x"0000" when x"A2D1",
			x"0000" when x"A2D2",
			x"0000" when x"A2D3",
			x"0000" when x"A2D4",
			x"0000" when x"A2D5",
			x"0000" when x"A2D6",
			x"0000" when x"A2D7",
			x"0000" when x"A2D8",
			x"0000" when x"A2D9",
			x"0000" when x"A2DA",
			x"0000" when x"A2DB",
			x"0000" when x"A2DC",
			x"0000" when x"A2DD",
			x"0000" when x"A2DE",
			x"0000" when x"A2DF",
			x"0000" when x"A2E0",
			x"0000" when x"A2E1",
			x"0000" when x"A2E2",
			x"0000" when x"A2E3",
			x"0000" when x"A2E4",
			x"0000" when x"A2E5",
			x"0000" when x"A2E6",
			x"0000" when x"A2E7",
			x"0000" when x"A2E8",
			x"0000" when x"A2E9",
			x"0000" when x"A2EA",
			x"0000" when x"A2EB",
			x"0000" when x"A2EC",
			x"0000" when x"A2ED",
			x"0000" when x"A2EE",
			x"0000" when x"A2EF",
			x"0000" when x"A2F0",
			x"0000" when x"A2F1",
			x"0000" when x"A2F2",
			x"0000" when x"A2F3",
			x"0000" when x"A2F4",
			x"0000" when x"A2F5",
			x"0000" when x"A2F6",
			x"0000" when x"A2F7",
			x"0000" when x"A2F8",
			x"0000" when x"A2F9",
			x"0000" when x"A2FA",
			x"0000" when x"A2FB",
			x"0000" when x"A2FC",
			x"0000" when x"A2FD",
			x"0000" when x"A2FE",
			x"0000" when x"A2FF",
			x"0000" when x"A300",
			x"0000" when x"A301",
			x"0000" when x"A302",
			x"0000" when x"A303",
			x"0000" when x"A304",
			x"0000" when x"A305",
			x"0000" when x"A306",
			x"0000" when x"A307",
			x"0000" when x"A308",
			x"0000" when x"A309",
			x"0000" when x"A30A",
			x"0000" when x"A30B",
			x"0000" when x"A30C",
			x"0000" when x"A30D",
			x"0000" when x"A30E",
			x"0000" when x"A30F",
			x"0000" when x"A310",
			x"0000" when x"A311",
			x"0000" when x"A312",
			x"0000" when x"A313",
			x"0000" when x"A314",
			x"0000" when x"A315",
			x"0000" when x"A316",
			x"0000" when x"A317",
			x"0000" when x"A318",
			x"0000" when x"A319",
			x"0000" when x"A31A",
			x"0000" when x"A31B",
			x"0000" when x"A31C",
			x"0000" when x"A31D",
			x"0000" when x"A31E",
			x"0000" when x"A31F",
			x"0000" when x"A320",
			x"0000" when x"A321",
			x"0000" when x"A322",
			x"0000" when x"A323",
			x"0000" when x"A324",
			x"0000" when x"A325",
			x"0000" when x"A326",
			x"0000" when x"A327",
			x"0000" when x"A328",
			x"0000" when x"A329",
			x"0000" when x"A32A",
			x"0000" when x"A32B",
			x"0000" when x"A32C",
			x"0000" when x"A32D",
			x"0000" when x"A32E",
			x"0000" when x"A32F",
			x"0000" when x"A330",
			x"0000" when x"A331",
			x"0000" when x"A332",
			x"0000" when x"A333",
			x"0000" when x"A334",
			x"0000" when x"A335",
			x"0000" when x"A336",
			x"0000" when x"A337",
			x"0000" when x"A338",
			x"0000" when x"A339",
			x"0000" when x"A33A",
			x"0000" when x"A33B",
			x"0000" when x"A33C",
			x"0000" when x"A33D",
			x"0000" when x"A33E",
			x"0000" when x"A33F",
			x"0000" when x"A340",
			x"0000" when x"A341",
			x"0000" when x"A342",
			x"0000" when x"A343",
			x"0000" when x"A344",
			x"0000" when x"A345",
			x"0000" when x"A346",
			x"0000" when x"A347",
			x"0000" when x"A348",
			x"0000" when x"A349",
			x"0000" when x"A34A",
			x"0000" when x"A34B",
			x"0000" when x"A34C",
			x"0000" when x"A34D",
			x"0000" when x"A34E",
			x"0000" when x"A34F",
			x"0000" when x"A350",
			x"0000" when x"A351",
			x"0000" when x"A352",
			x"0000" when x"A353",
			x"0000" when x"A354",
			x"0000" when x"A355",
			x"0000" when x"A356",
			x"0000" when x"A357",
			x"0000" when x"A358",
			x"0000" when x"A359",
			x"0000" when x"A35A",
			x"0000" when x"A35B",
			x"0000" when x"A35C",
			x"0000" when x"A35D",
			x"0000" when x"A35E",
			x"0000" when x"A35F",
			x"0000" when x"A360",
			x"0000" when x"A361",
			x"0000" when x"A362",
			x"0000" when x"A363",
			x"0000" when x"A364",
			x"0000" when x"A365",
			x"0000" when x"A366",
			x"0000" when x"A367",
			x"0000" when x"A368",
			x"0000" when x"A369",
			x"0000" when x"A36A",
			x"0000" when x"A36B",
			x"0000" when x"A36C",
			x"0000" when x"A36D",
			x"0000" when x"A36E",
			x"0000" when x"A36F",
			x"0000" when x"A370",
			x"0000" when x"A371",
			x"0000" when x"A372",
			x"0000" when x"A373",
			x"0000" when x"A374",
			x"0000" when x"A375",
			x"0000" when x"A376",
			x"0000" when x"A377",
			x"0000" when x"A378",
			x"0000" when x"A379",
			x"0000" when x"A37A",
			x"0000" when x"A37B",
			x"0000" when x"A37C",
			x"0000" when x"A37D",
			x"0000" when x"A37E",
			x"0000" when x"A37F",
			x"0000" when x"A380",
			x"0000" when x"A381",
			x"0000" when x"A382",
			x"0000" when x"A383",
			x"0000" when x"A384",
			x"0000" when x"A385",
			x"0000" when x"A386",
			x"0000" when x"A387",
			x"0000" when x"A388",
			x"0000" when x"A389",
			x"0000" when x"A38A",
			x"0000" when x"A38B",
			x"0000" when x"A38C",
			x"0000" when x"A38D",
			x"0000" when x"A38E",
			x"0000" when x"A38F",
			x"0000" when x"A390",
			x"0000" when x"A391",
			x"0000" when x"A392",
			x"0000" when x"A393",
			x"0000" when x"A394",
			x"0000" when x"A395",
			x"0000" when x"A396",
			x"0000" when x"A397",
			x"0000" when x"A398",
			x"0000" when x"A399",
			x"0000" when x"A39A",
			x"0000" when x"A39B",
			x"0000" when x"A39C",
			x"0000" when x"A39D",
			x"0000" when x"A39E",
			x"0000" when x"A39F",
			x"0000" when x"A3A0",
			x"0000" when x"A3A1",
			x"0000" when x"A3A2",
			x"0000" when x"A3A3",
			x"0000" when x"A3A4",
			x"0000" when x"A3A5",
			x"0000" when x"A3A6",
			x"0000" when x"A3A7",
			x"0000" when x"A3A8",
			x"0000" when x"A3A9",
			x"0000" when x"A3AA",
			x"0000" when x"A3AB",
			x"0000" when x"A3AC",
			x"0000" when x"A3AD",
			x"0000" when x"A3AE",
			x"0000" when x"A3AF",
			x"0000" when x"A3B0",
			x"0000" when x"A3B1",
			x"0000" when x"A3B2",
			x"0000" when x"A3B3",
			x"0000" when x"A3B4",
			x"0000" when x"A3B5",
			x"0000" when x"A3B6",
			x"0000" when x"A3B7",
			x"0000" when x"A3B8",
			x"0000" when x"A3B9",
			x"0000" when x"A3BA",
			x"0000" when x"A3BB",
			x"0000" when x"A3BC",
			x"0000" when x"A3BD",
			x"0000" when x"A3BE",
			x"0000" when x"A3BF",
			x"0000" when x"A3C0",
			x"0000" when x"A3C1",
			x"0000" when x"A3C2",
			x"0000" when x"A3C3",
			x"0000" when x"A3C4",
			x"0000" when x"A3C5",
			x"0000" when x"A3C6",
			x"0000" when x"A3C7",
			x"0000" when x"A3C8",
			x"0000" when x"A3C9",
			x"0000" when x"A3CA",
			x"0000" when x"A3CB",
			x"0000" when x"A3CC",
			x"0000" when x"A3CD",
			x"0000" when x"A3CE",
			x"0000" when x"A3CF",
			x"0000" when x"A3D0",
			x"0000" when x"A3D1",
			x"0000" when x"A3D2",
			x"0000" when x"A3D3",
			x"0000" when x"A3D4",
			x"0000" when x"A3D5",
			x"0000" when x"A3D6",
			x"0000" when x"A3D7",
			x"0000" when x"A3D8",
			x"0000" when x"A3D9",
			x"0000" when x"A3DA",
			x"0000" when x"A3DB",
			x"0000" when x"A3DC",
			x"0000" when x"A3DD",
			x"0000" when x"A3DE",
			x"0000" when x"A3DF",
			x"0000" when x"A3E0",
			x"0000" when x"A3E1",
			x"0000" when x"A3E2",
			x"0000" when x"A3E3",
			x"0000" when x"A3E4",
			x"0000" when x"A3E5",
			x"0000" when x"A3E6",
			x"0000" when x"A3E7",
			x"0000" when x"A3E8",
			x"0000" when x"A3E9",
			x"0000" when x"A3EA",
			x"0000" when x"A3EB",
			x"0000" when x"A3EC",
			x"0000" when x"A3ED",
			x"0000" when x"A3EE",
			x"0000" when x"A3EF",
			x"0000" when x"A3F0",
			x"0000" when x"A3F1",
			x"0000" when x"A3F2",
			x"0000" when x"A3F3",
			x"0000" when x"A3F4",
			x"0000" when x"A3F5",
			x"0000" when x"A3F6",
			x"0000" when x"A3F7",
			x"0000" when x"A3F8",
			x"0000" when x"A3F9",
			x"0000" when x"A3FA",
			x"0000" when x"A3FB",
			x"0000" when x"A3FC",
			x"0000" when x"A3FD",
			x"0000" when x"A3FE",
			x"0000" when x"A3FF",
			x"0000" when x"A400",
			x"0000" when x"A401",
			x"0000" when x"A402",
			x"0000" when x"A403",
			x"0000" when x"A404",
			x"0000" when x"A405",
			x"0000" when x"A406",
			x"0000" when x"A407",
			x"0000" when x"A408",
			x"0000" when x"A409",
			x"0000" when x"A40A",
			x"0000" when x"A40B",
			x"0000" when x"A40C",
			x"0000" when x"A40D",
			x"0000" when x"A40E",
			x"0000" when x"A40F",
			x"0000" when x"A410",
			x"0000" when x"A411",
			x"0000" when x"A412",
			x"0000" when x"A413",
			x"0000" when x"A414",
			x"0000" when x"A415",
			x"0000" when x"A416",
			x"0000" when x"A417",
			x"0000" when x"A418",
			x"0000" when x"A419",
			x"0000" when x"A41A",
			x"0000" when x"A41B",
			x"0000" when x"A41C",
			x"0000" when x"A41D",
			x"0000" when x"A41E",
			x"0000" when x"A41F",
			x"0000" when x"A420",
			x"0000" when x"A421",
			x"0000" when x"A422",
			x"0000" when x"A423",
			x"0000" when x"A424",
			x"0000" when x"A425",
			x"0000" when x"A426",
			x"0000" when x"A427",
			x"0000" when x"A428",
			x"0000" when x"A429",
			x"0000" when x"A42A",
			x"0000" when x"A42B",
			x"0000" when x"A42C",
			x"0000" when x"A42D",
			x"0000" when x"A42E",
			x"0000" when x"A42F",
			x"0000" when x"A430",
			x"0000" when x"A431",
			x"0000" when x"A432",
			x"0000" when x"A433",
			x"0000" when x"A434",
			x"0000" when x"A435",
			x"0000" when x"A436",
			x"0000" when x"A437",
			x"0000" when x"A438",
			x"0000" when x"A439",
			x"0000" when x"A43A",
			x"0000" when x"A43B",
			x"0000" when x"A43C",
			x"0000" when x"A43D",
			x"0000" when x"A43E",
			x"0000" when x"A43F",
			x"0000" when x"A440",
			x"0000" when x"A441",
			x"0000" when x"A442",
			x"0000" when x"A443",
			x"0000" when x"A444",
			x"0000" when x"A445",
			x"0000" when x"A446",
			x"0000" when x"A447",
			x"0000" when x"A448",
			x"0000" when x"A449",
			x"0000" when x"A44A",
			x"0000" when x"A44B",
			x"0000" when x"A44C",
			x"0000" when x"A44D",
			x"0000" when x"A44E",
			x"0000" when x"A44F",
			x"0000" when x"A450",
			x"0000" when x"A451",
			x"0000" when x"A452",
			x"0000" when x"A453",
			x"0000" when x"A454",
			x"0000" when x"A455",
			x"0000" when x"A456",
			x"0000" when x"A457",
			x"0000" when x"A458",
			x"0000" when x"A459",
			x"0000" when x"A45A",
			x"0000" when x"A45B",
			x"0000" when x"A45C",
			x"0000" when x"A45D",
			x"0000" when x"A45E",
			x"0000" when x"A45F",
			x"0000" when x"A460",
			x"0000" when x"A461",
			x"0000" when x"A462",
			x"0000" when x"A463",
			x"0000" when x"A464",
			x"0000" when x"A465",
			x"0000" when x"A466",
			x"0000" when x"A467",
			x"0000" when x"A468",
			x"0000" when x"A469",
			x"0000" when x"A46A",
			x"0000" when x"A46B",
			x"0000" when x"A46C",
			x"0000" when x"A46D",
			x"0000" when x"A46E",
			x"0000" when x"A46F",
			x"0000" when x"A470",
			x"0000" when x"A471",
			x"0000" when x"A472",
			x"0000" when x"A473",
			x"0000" when x"A474",
			x"0000" when x"A475",
			x"0000" when x"A476",
			x"0000" when x"A477",
			x"0000" when x"A478",
			x"0000" when x"A479",
			x"0000" when x"A47A",
			x"0000" when x"A47B",
			x"0000" when x"A47C",
			x"0000" when x"A47D",
			x"0000" when x"A47E",
			x"0000" when x"A47F",
			x"0000" when x"A480",
			x"0000" when x"A481",
			x"0000" when x"A482",
			x"0000" when x"A483",
			x"0000" when x"A484",
			x"0000" when x"A485",
			x"0000" when x"A486",
			x"0000" when x"A487",
			x"0000" when x"A488",
			x"0000" when x"A489",
			x"0000" when x"A48A",
			x"0000" when x"A48B",
			x"0000" when x"A48C",
			x"0000" when x"A48D",
			x"0000" when x"A48E",
			x"0000" when x"A48F",
			x"0000" when x"A490",
			x"0000" when x"A491",
			x"0000" when x"A492",
			x"0000" when x"A493",
			x"0000" when x"A494",
			x"0000" when x"A495",
			x"0000" when x"A496",
			x"0000" when x"A497",
			x"0000" when x"A498",
			x"0000" when x"A499",
			x"0000" when x"A49A",
			x"0000" when x"A49B",
			x"0000" when x"A49C",
			x"0000" when x"A49D",
			x"0000" when x"A49E",
			x"0000" when x"A49F",
			x"0000" when x"A4A0",
			x"0000" when x"A4A1",
			x"0000" when x"A4A2",
			x"0000" when x"A4A3",
			x"0000" when x"A4A4",
			x"0000" when x"A4A5",
			x"0000" when x"A4A6",
			x"0000" when x"A4A7",
			x"0000" when x"A4A8",
			x"0000" when x"A4A9",
			x"0000" when x"A4AA",
			x"0000" when x"A4AB",
			x"0000" when x"A4AC",
			x"0000" when x"A4AD",
			x"0000" when x"A4AE",
			x"0000" when x"A4AF",
			x"0000" when x"A4B0",
			x"0000" when x"A4B1",
			x"0000" when x"A4B2",
			x"0000" when x"A4B3",
			x"0000" when x"A4B4",
			x"0000" when x"A4B5",
			x"0000" when x"A4B6",
			x"0000" when x"A4B7",
			x"0000" when x"A4B8",
			x"0000" when x"A4B9",
			x"0000" when x"A4BA",
			x"0000" when x"A4BB",
			x"0000" when x"A4BC",
			x"0000" when x"A4BD",
			x"0000" when x"A4BE",
			x"0000" when x"A4BF",
			x"0000" when x"A4C0",
			x"0000" when x"A4C1",
			x"0000" when x"A4C2",
			x"0000" when x"A4C3",
			x"0000" when x"A4C4",
			x"0000" when x"A4C5",
			x"0000" when x"A4C6",
			x"0000" when x"A4C7",
			x"0000" when x"A4C8",
			x"0000" when x"A4C9",
			x"0000" when x"A4CA",
			x"0000" when x"A4CB",
			x"0000" when x"A4CC",
			x"0000" when x"A4CD",
			x"0000" when x"A4CE",
			x"0000" when x"A4CF",
			x"0000" when x"A4D0",
			x"0000" when x"A4D1",
			x"0000" when x"A4D2",
			x"0000" when x"A4D3",
			x"0000" when x"A4D4",
			x"0000" when x"A4D5",
			x"0000" when x"A4D6",
			x"0000" when x"A4D7",
			x"0000" when x"A4D8",
			x"0000" when x"A4D9",
			x"0000" when x"A4DA",
			x"0000" when x"A4DB",
			x"0000" when x"A4DC",
			x"0000" when x"A4DD",
			x"0000" when x"A4DE",
			x"0000" when x"A4DF",
			x"0000" when x"A4E0",
			x"0000" when x"A4E1",
			x"0000" when x"A4E2",
			x"0000" when x"A4E3",
			x"0000" when x"A4E4",
			x"0000" when x"A4E5",
			x"0000" when x"A4E6",
			x"0000" when x"A4E7",
			x"0000" when x"A4E8",
			x"0000" when x"A4E9",
			x"0000" when x"A4EA",
			x"0000" when x"A4EB",
			x"0000" when x"A4EC",
			x"0000" when x"A4ED",
			x"0000" when x"A4EE",
			x"0000" when x"A4EF",
			x"0000" when x"A4F0",
			x"0000" when x"A4F1",
			x"0000" when x"A4F2",
			x"0000" when x"A4F3",
			x"0000" when x"A4F4",
			x"0000" when x"A4F5",
			x"0000" when x"A4F6",
			x"0000" when x"A4F7",
			x"0000" when x"A4F8",
			x"0000" when x"A4F9",
			x"0000" when x"A4FA",
			x"0000" when x"A4FB",
			x"0000" when x"A4FC",
			x"0000" when x"A4FD",
			x"0000" when x"A4FE",
			x"0000" when x"A4FF",
			x"0000" when x"A500",
			x"0000" when x"A501",
			x"0000" when x"A502",
			x"0000" when x"A503",
			x"0000" when x"A504",
			x"0000" when x"A505",
			x"0000" when x"A506",
			x"0000" when x"A507",
			x"0000" when x"A508",
			x"0000" when x"A509",
			x"0000" when x"A50A",
			x"0000" when x"A50B",
			x"0000" when x"A50C",
			x"0000" when x"A50D",
			x"0000" when x"A50E",
			x"0000" when x"A50F",
			x"0000" when x"A510",
			x"0000" when x"A511",
			x"0000" when x"A512",
			x"0000" when x"A513",
			x"0000" when x"A514",
			x"0000" when x"A515",
			x"0000" when x"A516",
			x"0000" when x"A517",
			x"0000" when x"A518",
			x"0000" when x"A519",
			x"0000" when x"A51A",
			x"0000" when x"A51B",
			x"0000" when x"A51C",
			x"0000" when x"A51D",
			x"0000" when x"A51E",
			x"0000" when x"A51F",
			x"0000" when x"A520",
			x"0000" when x"A521",
			x"0000" when x"A522",
			x"0000" when x"A523",
			x"0000" when x"A524",
			x"0000" when x"A525",
			x"0000" when x"A526",
			x"0000" when x"A527",
			x"0000" when x"A528",
			x"0000" when x"A529",
			x"0000" when x"A52A",
			x"0000" when x"A52B",
			x"0000" when x"A52C",
			x"0000" when x"A52D",
			x"0000" when x"A52E",
			x"0000" when x"A52F",
			x"0000" when x"A530",
			x"0000" when x"A531",
			x"0000" when x"A532",
			x"0000" when x"A533",
			x"0000" when x"A534",
			x"0000" when x"A535",
			x"0000" when x"A536",
			x"0000" when x"A537",
			x"0000" when x"A538",
			x"0000" when x"A539",
			x"0000" when x"A53A",
			x"0000" when x"A53B",
			x"0000" when x"A53C",
			x"0000" when x"A53D",
			x"0000" when x"A53E",
			x"0000" when x"A53F",
			x"0000" when x"A540",
			x"0000" when x"A541",
			x"0000" when x"A542",
			x"0000" when x"A543",
			x"0000" when x"A544",
			x"0000" when x"A545",
			x"0000" when x"A546",
			x"0000" when x"A547",
			x"0000" when x"A548",
			x"0000" when x"A549",
			x"0000" when x"A54A",
			x"0000" when x"A54B",
			x"0000" when x"A54C",
			x"0000" when x"A54D",
			x"0000" when x"A54E",
			x"0000" when x"A54F",
			x"0000" when x"A550",
			x"0000" when x"A551",
			x"0000" when x"A552",
			x"0000" when x"A553",
			x"0000" when x"A554",
			x"0000" when x"A555",
			x"0000" when x"A556",
			x"0000" when x"A557",
			x"0000" when x"A558",
			x"0000" when x"A559",
			x"0000" when x"A55A",
			x"0000" when x"A55B",
			x"0000" when x"A55C",
			x"0000" when x"A55D",
			x"0000" when x"A55E",
			x"0000" when x"A55F",
			x"0000" when x"A560",
			x"0000" when x"A561",
			x"0000" when x"A562",
			x"0000" when x"A563",
			x"0000" when x"A564",
			x"0000" when x"A565",
			x"0000" when x"A566",
			x"0000" when x"A567",
			x"0000" when x"A568",
			x"0000" when x"A569",
			x"0000" when x"A56A",
			x"0000" when x"A56B",
			x"0000" when x"A56C",
			x"0000" when x"A56D",
			x"0000" when x"A56E",
			x"0000" when x"A56F",
			x"0000" when x"A570",
			x"0000" when x"A571",
			x"0000" when x"A572",
			x"0000" when x"A573",
			x"0000" when x"A574",
			x"0000" when x"A575",
			x"0000" when x"A576",
			x"0000" when x"A577",
			x"0000" when x"A578",
			x"0000" when x"A579",
			x"0000" when x"A57A",
			x"0000" when x"A57B",
			x"0000" when x"A57C",
			x"0000" when x"A57D",
			x"0000" when x"A57E",
			x"0000" when x"A57F",
			x"0000" when x"A580",
			x"0000" when x"A581",
			x"0000" when x"A582",
			x"0000" when x"A583",
			x"0000" when x"A584",
			x"0000" when x"A585",
			x"0000" when x"A586",
			x"0000" when x"A587",
			x"0000" when x"A588",
			x"0000" when x"A589",
			x"0000" when x"A58A",
			x"0000" when x"A58B",
			x"0000" when x"A58C",
			x"0000" when x"A58D",
			x"0000" when x"A58E",
			x"0000" when x"A58F",
			x"0000" when x"A590",
			x"0000" when x"A591",
			x"0000" when x"A592",
			x"0000" when x"A593",
			x"0000" when x"A594",
			x"0000" when x"A595",
			x"0000" when x"A596",
			x"0000" when x"A597",
			x"0000" when x"A598",
			x"0000" when x"A599",
			x"0000" when x"A59A",
			x"0000" when x"A59B",
			x"0000" when x"A59C",
			x"0000" when x"A59D",
			x"0000" when x"A59E",
			x"0000" when x"A59F",
			x"0000" when x"A5A0",
			x"0000" when x"A5A1",
			x"0000" when x"A5A2",
			x"0000" when x"A5A3",
			x"0000" when x"A5A4",
			x"0000" when x"A5A5",
			x"0000" when x"A5A6",
			x"0000" when x"A5A7",
			x"0000" when x"A5A8",
			x"0000" when x"A5A9",
			x"0000" when x"A5AA",
			x"0000" when x"A5AB",
			x"0000" when x"A5AC",
			x"0000" when x"A5AD",
			x"0000" when x"A5AE",
			x"0000" when x"A5AF",
			x"0000" when x"A5B0",
			x"0000" when x"A5B1",
			x"0000" when x"A5B2",
			x"0000" when x"A5B3",
			x"0000" when x"A5B4",
			x"0000" when x"A5B5",
			x"0000" when x"A5B6",
			x"0000" when x"A5B7",
			x"0000" when x"A5B8",
			x"0000" when x"A5B9",
			x"0000" when x"A5BA",
			x"0000" when x"A5BB",
			x"0000" when x"A5BC",
			x"0000" when x"A5BD",
			x"0000" when x"A5BE",
			x"0000" when x"A5BF",
			x"0000" when x"A5C0",
			x"0000" when x"A5C1",
			x"0000" when x"A5C2",
			x"0000" when x"A5C3",
			x"0000" when x"A5C4",
			x"0000" when x"A5C5",
			x"0000" when x"A5C6",
			x"0000" when x"A5C7",
			x"0000" when x"A5C8",
			x"0000" when x"A5C9",
			x"0000" when x"A5CA",
			x"0000" when x"A5CB",
			x"0000" when x"A5CC",
			x"0000" when x"A5CD",
			x"0000" when x"A5CE",
			x"0000" when x"A5CF",
			x"0000" when x"A5D0",
			x"0000" when x"A5D1",
			x"0000" when x"A5D2",
			x"0000" when x"A5D3",
			x"0000" when x"A5D4",
			x"0000" when x"A5D5",
			x"0000" when x"A5D6",
			x"0000" when x"A5D7",
			x"0000" when x"A5D8",
			x"0000" when x"A5D9",
			x"0000" when x"A5DA",
			x"0000" when x"A5DB",
			x"0000" when x"A5DC",
			x"0000" when x"A5DD",
			x"0000" when x"A5DE",
			x"0000" when x"A5DF",
			x"0000" when x"A5E0",
			x"0000" when x"A5E1",
			x"0000" when x"A5E2",
			x"0000" when x"A5E3",
			x"0000" when x"A5E4",
			x"0000" when x"A5E5",
			x"0000" when x"A5E6",
			x"0000" when x"A5E7",
			x"0000" when x"A5E8",
			x"0000" when x"A5E9",
			x"0000" when x"A5EA",
			x"0000" when x"A5EB",
			x"0000" when x"A5EC",
			x"0000" when x"A5ED",
			x"0000" when x"A5EE",
			x"0000" when x"A5EF",
			x"0000" when x"A5F0",
			x"0000" when x"A5F1",
			x"0000" when x"A5F2",
			x"0000" when x"A5F3",
			x"0000" when x"A5F4",
			x"0000" when x"A5F5",
			x"0000" when x"A5F6",
			x"0000" when x"A5F7",
			x"0000" when x"A5F8",
			x"0000" when x"A5F9",
			x"0000" when x"A5FA",
			x"0000" when x"A5FB",
			x"0000" when x"A5FC",
			x"0000" when x"A5FD",
			x"0000" when x"A5FE",
			x"0000" when x"A5FF",
			x"0000" when x"A600",
			x"0000" when x"A601",
			x"0000" when x"A602",
			x"0000" when x"A603",
			x"0000" when x"A604",
			x"0000" when x"A605",
			x"0000" when x"A606",
			x"0000" when x"A607",
			x"0000" when x"A608",
			x"0000" when x"A609",
			x"0000" when x"A60A",
			x"0000" when x"A60B",
			x"0000" when x"A60C",
			x"0000" when x"A60D",
			x"0000" when x"A60E",
			x"0000" when x"A60F",
			x"0000" when x"A610",
			x"0000" when x"A611",
			x"0000" when x"A612",
			x"0000" when x"A613",
			x"0000" when x"A614",
			x"0000" when x"A615",
			x"0000" when x"A616",
			x"0000" when x"A617",
			x"0000" when x"A618",
			x"0000" when x"A619",
			x"0000" when x"A61A",
			x"0000" when x"A61B",
			x"0000" when x"A61C",
			x"0000" when x"A61D",
			x"0000" when x"A61E",
			x"0000" when x"A61F",
			x"0000" when x"A620",
			x"0000" when x"A621",
			x"0000" when x"A622",
			x"0000" when x"A623",
			x"0000" when x"A624",
			x"0000" when x"A625",
			x"0000" when x"A626",
			x"0000" when x"A627",
			x"0000" when x"A628",
			x"0000" when x"A629",
			x"0000" when x"A62A",
			x"0000" when x"A62B",
			x"0000" when x"A62C",
			x"0000" when x"A62D",
			x"0000" when x"A62E",
			x"0000" when x"A62F",
			x"0000" when x"A630",
			x"0000" when x"A631",
			x"0000" when x"A632",
			x"0000" when x"A633",
			x"0000" when x"A634",
			x"0000" when x"A635",
			x"0000" when x"A636",
			x"0000" when x"A637",
			x"0000" when x"A638",
			x"0000" when x"A639",
			x"0000" when x"A63A",
			x"0000" when x"A63B",
			x"0000" when x"A63C",
			x"0000" when x"A63D",
			x"0000" when x"A63E",
			x"0000" when x"A63F",
			x"0000" when x"A640",
			x"0000" when x"A641",
			x"0000" when x"A642",
			x"0000" when x"A643",
			x"0000" when x"A644",
			x"0000" when x"A645",
			x"0000" when x"A646",
			x"0000" when x"A647",
			x"0000" when x"A648",
			x"0000" when x"A649",
			x"0000" when x"A64A",
			x"0000" when x"A64B",
			x"0000" when x"A64C",
			x"0000" when x"A64D",
			x"0000" when x"A64E",
			x"0000" when x"A64F",
			x"0000" when x"A650",
			x"0000" when x"A651",
			x"0000" when x"A652",
			x"0000" when x"A653",
			x"0000" when x"A654",
			x"0000" when x"A655",
			x"0000" when x"A656",
			x"0000" when x"A657",
			x"0000" when x"A658",
			x"0000" when x"A659",
			x"0000" when x"A65A",
			x"0000" when x"A65B",
			x"0000" when x"A65C",
			x"0000" when x"A65D",
			x"0000" when x"A65E",
			x"0000" when x"A65F",
			x"0000" when x"A660",
			x"0000" when x"A661",
			x"0000" when x"A662",
			x"0000" when x"A663",
			x"0000" when x"A664",
			x"0000" when x"A665",
			x"0000" when x"A666",
			x"0000" when x"A667",
			x"0000" when x"A668",
			x"0000" when x"A669",
			x"0000" when x"A66A",
			x"0000" when x"A66B",
			x"0000" when x"A66C",
			x"0000" when x"A66D",
			x"0000" when x"A66E",
			x"0000" when x"A66F",
			x"0000" when x"A670",
			x"0000" when x"A671",
			x"0000" when x"A672",
			x"0000" when x"A673",
			x"0000" when x"A674",
			x"0000" when x"A675",
			x"0000" when x"A676",
			x"0000" when x"A677",
			x"0000" when x"A678",
			x"0000" when x"A679",
			x"0000" when x"A67A",
			x"0000" when x"A67B",
			x"0000" when x"A67C",
			x"0000" when x"A67D",
			x"0000" when x"A67E",
			x"0000" when x"A67F",
			x"0000" when x"A680",
			x"0000" when x"A681",
			x"0000" when x"A682",
			x"0000" when x"A683",
			x"0000" when x"A684",
			x"0000" when x"A685",
			x"0000" when x"A686",
			x"0000" when x"A687",
			x"0000" when x"A688",
			x"0000" when x"A689",
			x"0000" when x"A68A",
			x"0000" when x"A68B",
			x"0000" when x"A68C",
			x"0000" when x"A68D",
			x"0000" when x"A68E",
			x"0000" when x"A68F",
			x"0000" when x"A690",
			x"0000" when x"A691",
			x"0000" when x"A692",
			x"0000" when x"A693",
			x"0000" when x"A694",
			x"0000" when x"A695",
			x"0000" when x"A696",
			x"0000" when x"A697",
			x"0000" when x"A698",
			x"0000" when x"A699",
			x"0000" when x"A69A",
			x"0000" when x"A69B",
			x"0000" when x"A69C",
			x"0000" when x"A69D",
			x"0000" when x"A69E",
			x"0000" when x"A69F",
			x"0000" when x"A6A0",
			x"0000" when x"A6A1",
			x"0000" when x"A6A2",
			x"0000" when x"A6A3",
			x"0000" when x"A6A4",
			x"0000" when x"A6A5",
			x"0000" when x"A6A6",
			x"0000" when x"A6A7",
			x"0000" when x"A6A8",
			x"0000" when x"A6A9",
			x"0000" when x"A6AA",
			x"0000" when x"A6AB",
			x"0000" when x"A6AC",
			x"0000" when x"A6AD",
			x"0000" when x"A6AE",
			x"0000" when x"A6AF",
			x"0000" when x"A6B0",
			x"0000" when x"A6B1",
			x"0000" when x"A6B2",
			x"0000" when x"A6B3",
			x"0000" when x"A6B4",
			x"0000" when x"A6B5",
			x"0000" when x"A6B6",
			x"0000" when x"A6B7",
			x"0000" when x"A6B8",
			x"0000" when x"A6B9",
			x"0000" when x"A6BA",
			x"0000" when x"A6BB",
			x"0000" when x"A6BC",
			x"0000" when x"A6BD",
			x"0000" when x"A6BE",
			x"0000" when x"A6BF",
			x"0000" when x"A6C0",
			x"0000" when x"A6C1",
			x"0000" when x"A6C2",
			x"0000" when x"A6C3",
			x"0000" when x"A6C4",
			x"0000" when x"A6C5",
			x"0000" when x"A6C6",
			x"0000" when x"A6C7",
			x"0000" when x"A6C8",
			x"0000" when x"A6C9",
			x"0000" when x"A6CA",
			x"0000" when x"A6CB",
			x"0000" when x"A6CC",
			x"0000" when x"A6CD",
			x"0000" when x"A6CE",
			x"0000" when x"A6CF",
			x"0000" when x"A6D0",
			x"0000" when x"A6D1",
			x"0000" when x"A6D2",
			x"0000" when x"A6D3",
			x"0000" when x"A6D4",
			x"0000" when x"A6D5",
			x"0000" when x"A6D6",
			x"0000" when x"A6D7",
			x"0000" when x"A6D8",
			x"0000" when x"A6D9",
			x"0000" when x"A6DA",
			x"0000" when x"A6DB",
			x"0000" when x"A6DC",
			x"0000" when x"A6DD",
			x"0000" when x"A6DE",
			x"0000" when x"A6DF",
			x"0000" when x"A6E0",
			x"0000" when x"A6E1",
			x"0000" when x"A6E2",
			x"0000" when x"A6E3",
			x"0000" when x"A6E4",
			x"0000" when x"A6E5",
			x"0000" when x"A6E6",
			x"0000" when x"A6E7",
			x"0000" when x"A6E8",
			x"0000" when x"A6E9",
			x"0000" when x"A6EA",
			x"0000" when x"A6EB",
			x"0000" when x"A6EC",
			x"0000" when x"A6ED",
			x"0000" when x"A6EE",
			x"0000" when x"A6EF",
			x"0000" when x"A6F0",
			x"0000" when x"A6F1",
			x"0000" when x"A6F2",
			x"0000" when x"A6F3",
			x"0000" when x"A6F4",
			x"0000" when x"A6F5",
			x"0000" when x"A6F6",
			x"0000" when x"A6F7",
			x"0000" when x"A6F8",
			x"0000" when x"A6F9",
			x"0000" when x"A6FA",
			x"0000" when x"A6FB",
			x"0000" when x"A6FC",
			x"0000" when x"A6FD",
			x"0000" when x"A6FE",
			x"0000" when x"A6FF",
			x"0000" when x"A700",
			x"0000" when x"A701",
			x"0000" when x"A702",
			x"0000" when x"A703",
			x"0000" when x"A704",
			x"0000" when x"A705",
			x"0000" when x"A706",
			x"0000" when x"A707",
			x"0000" when x"A708",
			x"0000" when x"A709",
			x"0000" when x"A70A",
			x"0000" when x"A70B",
			x"0000" when x"A70C",
			x"0000" when x"A70D",
			x"0000" when x"A70E",
			x"0000" when x"A70F",
			x"0000" when x"A710",
			x"0000" when x"A711",
			x"0000" when x"A712",
			x"0000" when x"A713",
			x"0000" when x"A714",
			x"0000" when x"A715",
			x"0000" when x"A716",
			x"0000" when x"A717",
			x"0000" when x"A718",
			x"0000" when x"A719",
			x"0000" when x"A71A",
			x"0000" when x"A71B",
			x"0000" when x"A71C",
			x"0000" when x"A71D",
			x"0000" when x"A71E",
			x"0000" when x"A71F",
			x"0000" when x"A720",
			x"0000" when x"A721",
			x"0000" when x"A722",
			x"0000" when x"A723",
			x"0000" when x"A724",
			x"0000" when x"A725",
			x"0000" when x"A726",
			x"0000" when x"A727",
			x"0000" when x"A728",
			x"0000" when x"A729",
			x"0000" when x"A72A",
			x"0000" when x"A72B",
			x"0000" when x"A72C",
			x"0000" when x"A72D",
			x"0000" when x"A72E",
			x"0000" when x"A72F",
			x"0000" when x"A730",
			x"0000" when x"A731",
			x"0000" when x"A732",
			x"0000" when x"A733",
			x"0000" when x"A734",
			x"0000" when x"A735",
			x"0000" when x"A736",
			x"0000" when x"A737",
			x"0000" when x"A738",
			x"0000" when x"A739",
			x"0000" when x"A73A",
			x"0000" when x"A73B",
			x"0000" when x"A73C",
			x"0000" when x"A73D",
			x"0000" when x"A73E",
			x"0000" when x"A73F",
			x"0000" when x"A740",
			x"0000" when x"A741",
			x"0000" when x"A742",
			x"0000" when x"A743",
			x"0000" when x"A744",
			x"0000" when x"A745",
			x"0000" when x"A746",
			x"0000" when x"A747",
			x"0000" when x"A748",
			x"0000" when x"A749",
			x"0000" when x"A74A",
			x"0000" when x"A74B",
			x"0000" when x"A74C",
			x"0000" when x"A74D",
			x"0000" when x"A74E",
			x"0000" when x"A74F",
			x"0000" when x"A750",
			x"0000" when x"A751",
			x"0000" when x"A752",
			x"0000" when x"A753",
			x"0000" when x"A754",
			x"0000" when x"A755",
			x"0000" when x"A756",
			x"0000" when x"A757",
			x"0000" when x"A758",
			x"0000" when x"A759",
			x"0000" when x"A75A",
			x"0000" when x"A75B",
			x"0000" when x"A75C",
			x"0000" when x"A75D",
			x"0000" when x"A75E",
			x"0000" when x"A75F",
			x"0000" when x"A760",
			x"0000" when x"A761",
			x"0000" when x"A762",
			x"0000" when x"A763",
			x"0000" when x"A764",
			x"0000" when x"A765",
			x"0000" when x"A766",
			x"0000" when x"A767",
			x"0000" when x"A768",
			x"0000" when x"A769",
			x"0000" when x"A76A",
			x"0000" when x"A76B",
			x"0000" when x"A76C",
			x"0000" when x"A76D",
			x"0000" when x"A76E",
			x"0000" when x"A76F",
			x"0000" when x"A770",
			x"0000" when x"A771",
			x"0000" when x"A772",
			x"0000" when x"A773",
			x"0000" when x"A774",
			x"0000" when x"A775",
			x"0000" when x"A776",
			x"0000" when x"A777",
			x"0000" when x"A778",
			x"0000" when x"A779",
			x"0000" when x"A77A",
			x"0000" when x"A77B",
			x"0000" when x"A77C",
			x"0000" when x"A77D",
			x"0000" when x"A77E",
			x"0000" when x"A77F",
			x"0000" when x"A780",
			x"0000" when x"A781",
			x"0000" when x"A782",
			x"0000" when x"A783",
			x"0000" when x"A784",
			x"0000" when x"A785",
			x"0000" when x"A786",
			x"0000" when x"A787",
			x"0000" when x"A788",
			x"0000" when x"A789",
			x"0000" when x"A78A",
			x"0000" when x"A78B",
			x"0000" when x"A78C",
			x"0000" when x"A78D",
			x"0000" when x"A78E",
			x"0000" when x"A78F",
			x"0000" when x"A790",
			x"0000" when x"A791",
			x"0000" when x"A792",
			x"0000" when x"A793",
			x"0000" when x"A794",
			x"0000" when x"A795",
			x"0000" when x"A796",
			x"0000" when x"A797",
			x"0000" when x"A798",
			x"0000" when x"A799",
			x"0000" when x"A79A",
			x"0000" when x"A79B",
			x"0000" when x"A79C",
			x"0000" when x"A79D",
			x"0000" when x"A79E",
			x"0000" when x"A79F",
			x"0000" when x"A7A0",
			x"0000" when x"A7A1",
			x"0000" when x"A7A2",
			x"0000" when x"A7A3",
			x"0000" when x"A7A4",
			x"0000" when x"A7A5",
			x"0000" when x"A7A6",
			x"0000" when x"A7A7",
			x"0000" when x"A7A8",
			x"0000" when x"A7A9",
			x"0000" when x"A7AA",
			x"0000" when x"A7AB",
			x"0000" when x"A7AC",
			x"0000" when x"A7AD",
			x"0000" when x"A7AE",
			x"0000" when x"A7AF",
			x"0000" when x"A7B0",
			x"0000" when x"A7B1",
			x"0000" when x"A7B2",
			x"0000" when x"A7B3",
			x"0000" when x"A7B4",
			x"0000" when x"A7B5",
			x"0000" when x"A7B6",
			x"0000" when x"A7B7",
			x"0000" when x"A7B8",
			x"0000" when x"A7B9",
			x"0000" when x"A7BA",
			x"0000" when x"A7BB",
			x"0000" when x"A7BC",
			x"0000" when x"A7BD",
			x"0000" when x"A7BE",
			x"0000" when x"A7BF",
			x"0000" when x"A7C0",
			x"0000" when x"A7C1",
			x"0000" when x"A7C2",
			x"0000" when x"A7C3",
			x"0000" when x"A7C4",
			x"0000" when x"A7C5",
			x"0000" when x"A7C6",
			x"0000" when x"A7C7",
			x"0000" when x"A7C8",
			x"0000" when x"A7C9",
			x"0000" when x"A7CA",
			x"0000" when x"A7CB",
			x"0000" when x"A7CC",
			x"0000" when x"A7CD",
			x"0000" when x"A7CE",
			x"0000" when x"A7CF",
			x"0000" when x"A7D0",
			x"0000" when x"A7D1",
			x"0000" when x"A7D2",
			x"0000" when x"A7D3",
			x"0000" when x"A7D4",
			x"0000" when x"A7D5",
			x"0000" when x"A7D6",
			x"0000" when x"A7D7",
			x"0000" when x"A7D8",
			x"0000" when x"A7D9",
			x"0000" when x"A7DA",
			x"0000" when x"A7DB",
			x"0000" when x"A7DC",
			x"0000" when x"A7DD",
			x"0000" when x"A7DE",
			x"0000" when x"A7DF",
			x"0000" when x"A7E0",
			x"0000" when x"A7E1",
			x"0000" when x"A7E2",
			x"0000" when x"A7E3",
			x"0000" when x"A7E4",
			x"0000" when x"A7E5",
			x"0000" when x"A7E6",
			x"0000" when x"A7E7",
			x"0000" when x"A7E8",
			x"0000" when x"A7E9",
			x"0000" when x"A7EA",
			x"0000" when x"A7EB",
			x"0000" when x"A7EC",
			x"0000" when x"A7ED",
			x"0000" when x"A7EE",
			x"0000" when x"A7EF",
			x"0000" when x"A7F0",
			x"0000" when x"A7F1",
			x"0000" when x"A7F2",
			x"0000" when x"A7F3",
			x"0000" when x"A7F4",
			x"0000" when x"A7F5",
			x"0000" when x"A7F6",
			x"0000" when x"A7F7",
			x"0000" when x"A7F8",
			x"0000" when x"A7F9",
			x"0000" when x"A7FA",
			x"0000" when x"A7FB",
			x"0000" when x"A7FC",
			x"0000" when x"A7FD",
			x"0000" when x"A7FE",
			x"0000" when x"A7FF",
			x"0000" when x"A800",
			x"0000" when x"A801",
			x"0000" when x"A802",
			x"0000" when x"A803",
			x"0000" when x"A804",
			x"0000" when x"A805",
			x"0000" when x"A806",
			x"0000" when x"A807",
			x"0000" when x"A808",
			x"0000" when x"A809",
			x"0000" when x"A80A",
			x"0000" when x"A80B",
			x"0000" when x"A80C",
			x"0000" when x"A80D",
			x"0000" when x"A80E",
			x"0000" when x"A80F",
			x"0000" when x"A810",
			x"0000" when x"A811",
			x"0000" when x"A812",
			x"0000" when x"A813",
			x"0000" when x"A814",
			x"0000" when x"A815",
			x"0000" when x"A816",
			x"0000" when x"A817",
			x"0000" when x"A818",
			x"0000" when x"A819",
			x"0000" when x"A81A",
			x"0000" when x"A81B",
			x"0000" when x"A81C",
			x"0000" when x"A81D",
			x"0000" when x"A81E",
			x"0000" when x"A81F",
			x"0000" when x"A820",
			x"0000" when x"A821",
			x"0000" when x"A822",
			x"0000" when x"A823",
			x"0000" when x"A824",
			x"0000" when x"A825",
			x"0000" when x"A826",
			x"0000" when x"A827",
			x"0000" when x"A828",
			x"0000" when x"A829",
			x"0000" when x"A82A",
			x"0000" when x"A82B",
			x"0000" when x"A82C",
			x"0000" when x"A82D",
			x"0000" when x"A82E",
			x"0000" when x"A82F",
			x"0000" when x"A830",
			x"0000" when x"A831",
			x"0000" when x"A832",
			x"0000" when x"A833",
			x"0000" when x"A834",
			x"0000" when x"A835",
			x"0000" when x"A836",
			x"0000" when x"A837",
			x"0000" when x"A838",
			x"0000" when x"A839",
			x"0000" when x"A83A",
			x"0000" when x"A83B",
			x"0000" when x"A83C",
			x"0000" when x"A83D",
			x"0000" when x"A83E",
			x"0000" when x"A83F",
			x"0000" when x"A840",
			x"0000" when x"A841",
			x"0000" when x"A842",
			x"0000" when x"A843",
			x"0000" when x"A844",
			x"0000" when x"A845",
			x"0000" when x"A846",
			x"0000" when x"A847",
			x"0000" when x"A848",
			x"0000" when x"A849",
			x"0000" when x"A84A",
			x"0000" when x"A84B",
			x"0000" when x"A84C",
			x"0000" when x"A84D",
			x"0000" when x"A84E",
			x"0000" when x"A84F",
			x"0000" when x"A850",
			x"0000" when x"A851",
			x"0000" when x"A852",
			x"0000" when x"A853",
			x"0000" when x"A854",
			x"0000" when x"A855",
			x"0000" when x"A856",
			x"0000" when x"A857",
			x"0000" when x"A858",
			x"0000" when x"A859",
			x"0000" when x"A85A",
			x"0000" when x"A85B",
			x"0000" when x"A85C",
			x"0000" when x"A85D",
			x"0000" when x"A85E",
			x"0000" when x"A85F",
			x"0000" when x"A860",
			x"0000" when x"A861",
			x"0000" when x"A862",
			x"0000" when x"A863",
			x"0000" when x"A864",
			x"0000" when x"A865",
			x"0000" when x"A866",
			x"0000" when x"A867",
			x"0000" when x"A868",
			x"0000" when x"A869",
			x"0000" when x"A86A",
			x"0000" when x"A86B",
			x"0000" when x"A86C",
			x"0000" when x"A86D",
			x"0000" when x"A86E",
			x"0000" when x"A86F",
			x"0000" when x"A870",
			x"0000" when x"A871",
			x"0000" when x"A872",
			x"0000" when x"A873",
			x"0000" when x"A874",
			x"0000" when x"A875",
			x"0000" when x"A876",
			x"0000" when x"A877",
			x"0000" when x"A878",
			x"0000" when x"A879",
			x"0000" when x"A87A",
			x"0000" when x"A87B",
			x"0000" when x"A87C",
			x"0000" when x"A87D",
			x"0000" when x"A87E",
			x"0000" when x"A87F",
			x"0000" when x"A880",
			x"0000" when x"A881",
			x"0000" when x"A882",
			x"0000" when x"A883",
			x"0000" when x"A884",
			x"0000" when x"A885",
			x"0000" when x"A886",
			x"0000" when x"A887",
			x"0000" when x"A888",
			x"0000" when x"A889",
			x"0000" when x"A88A",
			x"0000" when x"A88B",
			x"0000" when x"A88C",
			x"0000" when x"A88D",
			x"0000" when x"A88E",
			x"0000" when x"A88F",
			x"0000" when x"A890",
			x"0000" when x"A891",
			x"0000" when x"A892",
			x"0000" when x"A893",
			x"0000" when x"A894",
			x"0000" when x"A895",
			x"0000" when x"A896",
			x"0000" when x"A897",
			x"0000" when x"A898",
			x"0000" when x"A899",
			x"0000" when x"A89A",
			x"0000" when x"A89B",
			x"0000" when x"A89C",
			x"0000" when x"A89D",
			x"0000" when x"A89E",
			x"0000" when x"A89F",
			x"0000" when x"A8A0",
			x"0000" when x"A8A1",
			x"0000" when x"A8A2",
			x"0000" when x"A8A3",
			x"0000" when x"A8A4",
			x"0000" when x"A8A5",
			x"0000" when x"A8A6",
			x"0000" when x"A8A7",
			x"0000" when x"A8A8",
			x"0000" when x"A8A9",
			x"0000" when x"A8AA",
			x"0000" when x"A8AB",
			x"0000" when x"A8AC",
			x"0000" when x"A8AD",
			x"0000" when x"A8AE",
			x"0000" when x"A8AF",
			x"0000" when x"A8B0",
			x"0000" when x"A8B1",
			x"0000" when x"A8B2",
			x"0000" when x"A8B3",
			x"0000" when x"A8B4",
			x"0000" when x"A8B5",
			x"0000" when x"A8B6",
			x"0000" when x"A8B7",
			x"0000" when x"A8B8",
			x"0000" when x"A8B9",
			x"0000" when x"A8BA",
			x"0000" when x"A8BB",
			x"0000" when x"A8BC",
			x"0000" when x"A8BD",
			x"0000" when x"A8BE",
			x"0000" when x"A8BF",
			x"0000" when x"A8C0",
			x"0000" when x"A8C1",
			x"0000" when x"A8C2",
			x"0000" when x"A8C3",
			x"0000" when x"A8C4",
			x"0000" when x"A8C5",
			x"0000" when x"A8C6",
			x"0000" when x"A8C7",
			x"0000" when x"A8C8",
			x"0000" when x"A8C9",
			x"0000" when x"A8CA",
			x"0000" when x"A8CB",
			x"0000" when x"A8CC",
			x"0000" when x"A8CD",
			x"0000" when x"A8CE",
			x"0000" when x"A8CF",
			x"0000" when x"A8D0",
			x"0000" when x"A8D1",
			x"0000" when x"A8D2",
			x"0000" when x"A8D3",
			x"0000" when x"A8D4",
			x"0000" when x"A8D5",
			x"0000" when x"A8D6",
			x"0000" when x"A8D7",
			x"0000" when x"A8D8",
			x"0000" when x"A8D9",
			x"0000" when x"A8DA",
			x"0000" when x"A8DB",
			x"0000" when x"A8DC",
			x"0000" when x"A8DD",
			x"0000" when x"A8DE",
			x"0000" when x"A8DF",
			x"0000" when x"A8E0",
			x"0000" when x"A8E1",
			x"0000" when x"A8E2",
			x"0000" when x"A8E3",
			x"0000" when x"A8E4",
			x"0000" when x"A8E5",
			x"0000" when x"A8E6",
			x"0000" when x"A8E7",
			x"0000" when x"A8E8",
			x"0000" when x"A8E9",
			x"0000" when x"A8EA",
			x"0000" when x"A8EB",
			x"0000" when x"A8EC",
			x"0000" when x"A8ED",
			x"0000" when x"A8EE",
			x"0000" when x"A8EF",
			x"0000" when x"A8F0",
			x"0000" when x"A8F1",
			x"0000" when x"A8F2",
			x"0000" when x"A8F3",
			x"0000" when x"A8F4",
			x"0000" when x"A8F5",
			x"0000" when x"A8F6",
			x"0000" when x"A8F7",
			x"0000" when x"A8F8",
			x"0000" when x"A8F9",
			x"0000" when x"A8FA",
			x"0000" when x"A8FB",
			x"0000" when x"A8FC",
			x"0000" when x"A8FD",
			x"0000" when x"A8FE",
			x"0000" when x"A8FF",
			x"0000" when x"A900",
			x"0000" when x"A901",
			x"0000" when x"A902",
			x"0000" when x"A903",
			x"0000" when x"A904",
			x"0000" when x"A905",
			x"0000" when x"A906",
			x"0000" when x"A907",
			x"0000" when x"A908",
			x"0000" when x"A909",
			x"0000" when x"A90A",
			x"0000" when x"A90B",
			x"0000" when x"A90C",
			x"0000" when x"A90D",
			x"0000" when x"A90E",
			x"0000" when x"A90F",
			x"0000" when x"A910",
			x"0000" when x"A911",
			x"0000" when x"A912",
			x"0000" when x"A913",
			x"0000" when x"A914",
			x"0000" when x"A915",
			x"0000" when x"A916",
			x"0000" when x"A917",
			x"0000" when x"A918",
			x"0000" when x"A919",
			x"0000" when x"A91A",
			x"0000" when x"A91B",
			x"0000" when x"A91C",
			x"0000" when x"A91D",
			x"0000" when x"A91E",
			x"0000" when x"A91F",
			x"0000" when x"A920",
			x"0000" when x"A921",
			x"0000" when x"A922",
			x"0000" when x"A923",
			x"0000" when x"A924",
			x"0000" when x"A925",
			x"0000" when x"A926",
			x"0000" when x"A927",
			x"0000" when x"A928",
			x"0000" when x"A929",
			x"0000" when x"A92A",
			x"0000" when x"A92B",
			x"0000" when x"A92C",
			x"0000" when x"A92D",
			x"0000" when x"A92E",
			x"0000" when x"A92F",
			x"0000" when x"A930",
			x"0000" when x"A931",
			x"0000" when x"A932",
			x"0000" when x"A933",
			x"0000" when x"A934",
			x"0000" when x"A935",
			x"0000" when x"A936",
			x"0000" when x"A937",
			x"0000" when x"A938",
			x"0000" when x"A939",
			x"0000" when x"A93A",
			x"0000" when x"A93B",
			x"0000" when x"A93C",
			x"0000" when x"A93D",
			x"0000" when x"A93E",
			x"0000" when x"A93F",
			x"0000" when x"A940",
			x"0000" when x"A941",
			x"0000" when x"A942",
			x"0000" when x"A943",
			x"0000" when x"A944",
			x"0000" when x"A945",
			x"0000" when x"A946",
			x"0000" when x"A947",
			x"0000" when x"A948",
			x"0000" when x"A949",
			x"0000" when x"A94A",
			x"0000" when x"A94B",
			x"0000" when x"A94C",
			x"0000" when x"A94D",
			x"0000" when x"A94E",
			x"0000" when x"A94F",
			x"0000" when x"A950",
			x"0000" when x"A951",
			x"0000" when x"A952",
			x"0000" when x"A953",
			x"0000" when x"A954",
			x"0000" when x"A955",
			x"0000" when x"A956",
			x"0000" when x"A957",
			x"0000" when x"A958",
			x"0000" when x"A959",
			x"0000" when x"A95A",
			x"0000" when x"A95B",
			x"0000" when x"A95C",
			x"0000" when x"A95D",
			x"0000" when x"A95E",
			x"0000" when x"A95F",
			x"0000" when x"A960",
			x"0000" when x"A961",
			x"0000" when x"A962",
			x"0000" when x"A963",
			x"0000" when x"A964",
			x"0000" when x"A965",
			x"0000" when x"A966",
			x"0000" when x"A967",
			x"0000" when x"A968",
			x"0000" when x"A969",
			x"0000" when x"A96A",
			x"0000" when x"A96B",
			x"0000" when x"A96C",
			x"0000" when x"A96D",
			x"0000" when x"A96E",
			x"0000" when x"A96F",
			x"0000" when x"A970",
			x"0000" when x"A971",
			x"0000" when x"A972",
			x"0000" when x"A973",
			x"0000" when x"A974",
			x"0000" when x"A975",
			x"0000" when x"A976",
			x"0000" when x"A977",
			x"0000" when x"A978",
			x"0000" when x"A979",
			x"0000" when x"A97A",
			x"0000" when x"A97B",
			x"0000" when x"A97C",
			x"0000" when x"A97D",
			x"0000" when x"A97E",
			x"0000" when x"A97F",
			x"0000" when x"A980",
			x"0000" when x"A981",
			x"0000" when x"A982",
			x"0000" when x"A983",
			x"0000" when x"A984",
			x"0000" when x"A985",
			x"0000" when x"A986",
			x"0000" when x"A987",
			x"0000" when x"A988",
			x"0000" when x"A989",
			x"0000" when x"A98A",
			x"0000" when x"A98B",
			x"0000" when x"A98C",
			x"0000" when x"A98D",
			x"0000" when x"A98E",
			x"0000" when x"A98F",
			x"0000" when x"A990",
			x"0000" when x"A991",
			x"0000" when x"A992",
			x"0000" when x"A993",
			x"0000" when x"A994",
			x"0000" when x"A995",
			x"0000" when x"A996",
			x"0000" when x"A997",
			x"0000" when x"A998",
			x"0000" when x"A999",
			x"0000" when x"A99A",
			x"0000" when x"A99B",
			x"0000" when x"A99C",
			x"0000" when x"A99D",
			x"0000" when x"A99E",
			x"0000" when x"A99F",
			x"0000" when x"A9A0",
			x"0000" when x"A9A1",
			x"0000" when x"A9A2",
			x"0000" when x"A9A3",
			x"0000" when x"A9A4",
			x"0000" when x"A9A5",
			x"0000" when x"A9A6",
			x"0000" when x"A9A7",
			x"0000" when x"A9A8",
			x"0000" when x"A9A9",
			x"0000" when x"A9AA",
			x"0000" when x"A9AB",
			x"0000" when x"A9AC",
			x"0000" when x"A9AD",
			x"0000" when x"A9AE",
			x"0000" when x"A9AF",
			x"0000" when x"A9B0",
			x"0000" when x"A9B1",
			x"0000" when x"A9B2",
			x"0000" when x"A9B3",
			x"0000" when x"A9B4",
			x"0000" when x"A9B5",
			x"0000" when x"A9B6",
			x"0000" when x"A9B7",
			x"0000" when x"A9B8",
			x"0000" when x"A9B9",
			x"0000" when x"A9BA",
			x"0000" when x"A9BB",
			x"0000" when x"A9BC",
			x"0000" when x"A9BD",
			x"0000" when x"A9BE",
			x"0000" when x"A9BF",
			x"0000" when x"A9C0",
			x"0000" when x"A9C1",
			x"0000" when x"A9C2",
			x"0000" when x"A9C3",
			x"0000" when x"A9C4",
			x"0000" when x"A9C5",
			x"0000" when x"A9C6",
			x"0000" when x"A9C7",
			x"0000" when x"A9C8",
			x"0000" when x"A9C9",
			x"0000" when x"A9CA",
			x"0000" when x"A9CB",
			x"0000" when x"A9CC",
			x"0000" when x"A9CD",
			x"0000" when x"A9CE",
			x"0000" when x"A9CF",
			x"0000" when x"A9D0",
			x"0000" when x"A9D1",
			x"0000" when x"A9D2",
			x"0000" when x"A9D3",
			x"0000" when x"A9D4",
			x"0000" when x"A9D5",
			x"0000" when x"A9D6",
			x"0000" when x"A9D7",
			x"0000" when x"A9D8",
			x"0000" when x"A9D9",
			x"0000" when x"A9DA",
			x"0000" when x"A9DB",
			x"0000" when x"A9DC",
			x"0000" when x"A9DD",
			x"0000" when x"A9DE",
			x"0000" when x"A9DF",
			x"0000" when x"A9E0",
			x"0000" when x"A9E1",
			x"0000" when x"A9E2",
			x"0000" when x"A9E3",
			x"0000" when x"A9E4",
			x"0000" when x"A9E5",
			x"0000" when x"A9E6",
			x"0000" when x"A9E7",
			x"0000" when x"A9E8",
			x"0000" when x"A9E9",
			x"0000" when x"A9EA",
			x"0000" when x"A9EB",
			x"0000" when x"A9EC",
			x"0000" when x"A9ED",
			x"0000" when x"A9EE",
			x"0000" when x"A9EF",
			x"0000" when x"A9F0",
			x"0000" when x"A9F1",
			x"0000" when x"A9F2",
			x"0000" when x"A9F3",
			x"0000" when x"A9F4",
			x"0000" when x"A9F5",
			x"0000" when x"A9F6",
			x"0000" when x"A9F7",
			x"0000" when x"A9F8",
			x"0000" when x"A9F9",
			x"0000" when x"A9FA",
			x"0000" when x"A9FB",
			x"0000" when x"A9FC",
			x"0000" when x"A9FD",
			x"0000" when x"A9FE",
			x"0000" when x"A9FF",
			x"0000" when x"AA00",
			x"0000" when x"AA01",
			x"0000" when x"AA02",
			x"0000" when x"AA03",
			x"0000" when x"AA04",
			x"0000" when x"AA05",
			x"0000" when x"AA06",
			x"0000" when x"AA07",
			x"0000" when x"AA08",
			x"0000" when x"AA09",
			x"0000" when x"AA0A",
			x"0000" when x"AA0B",
			x"0000" when x"AA0C",
			x"0000" when x"AA0D",
			x"0000" when x"AA0E",
			x"0000" when x"AA0F",
			x"0000" when x"AA10",
			x"0000" when x"AA11",
			x"0000" when x"AA12",
			x"0000" when x"AA13",
			x"0000" when x"AA14",
			x"0000" when x"AA15",
			x"0000" when x"AA16",
			x"0000" when x"AA17",
			x"0000" when x"AA18",
			x"0000" when x"AA19",
			x"0000" when x"AA1A",
			x"0000" when x"AA1B",
			x"0000" when x"AA1C",
			x"0000" when x"AA1D",
			x"0000" when x"AA1E",
			x"0000" when x"AA1F",
			x"0000" when x"AA20",
			x"0000" when x"AA21",
			x"0000" when x"AA22",
			x"0000" when x"AA23",
			x"0000" when x"AA24",
			x"0000" when x"AA25",
			x"0000" when x"AA26",
			x"0000" when x"AA27",
			x"0000" when x"AA28",
			x"0000" when x"AA29",
			x"0000" when x"AA2A",
			x"0000" when x"AA2B",
			x"0000" when x"AA2C",
			x"0000" when x"AA2D",
			x"0000" when x"AA2E",
			x"0000" when x"AA2F",
			x"0000" when x"AA30",
			x"0000" when x"AA31",
			x"0000" when x"AA32",
			x"0000" when x"AA33",
			x"0000" when x"AA34",
			x"0000" when x"AA35",
			x"0000" when x"AA36",
			x"0000" when x"AA37",
			x"0000" when x"AA38",
			x"0000" when x"AA39",
			x"0000" when x"AA3A",
			x"0000" when x"AA3B",
			x"0000" when x"AA3C",
			x"0000" when x"AA3D",
			x"0000" when x"AA3E",
			x"0000" when x"AA3F",
			x"0000" when x"AA40",
			x"0000" when x"AA41",
			x"0000" when x"AA42",
			x"0000" when x"AA43",
			x"0000" when x"AA44",
			x"0000" when x"AA45",
			x"0000" when x"AA46",
			x"0000" when x"AA47",
			x"0000" when x"AA48",
			x"0000" when x"AA49",
			x"0000" when x"AA4A",
			x"0000" when x"AA4B",
			x"0000" when x"AA4C",
			x"0000" when x"AA4D",
			x"0000" when x"AA4E",
			x"0000" when x"AA4F",
			x"0000" when x"AA50",
			x"0000" when x"AA51",
			x"0000" when x"AA52",
			x"0000" when x"AA53",
			x"0000" when x"AA54",
			x"0000" when x"AA55",
			x"0000" when x"AA56",
			x"0000" when x"AA57",
			x"0000" when x"AA58",
			x"0000" when x"AA59",
			x"0000" when x"AA5A",
			x"0000" when x"AA5B",
			x"0000" when x"AA5C",
			x"0000" when x"AA5D",
			x"0000" when x"AA5E",
			x"0000" when x"AA5F",
			x"0000" when x"AA60",
			x"0000" when x"AA61",
			x"0000" when x"AA62",
			x"0000" when x"AA63",
			x"0000" when x"AA64",
			x"0000" when x"AA65",
			x"0000" when x"AA66",
			x"0000" when x"AA67",
			x"0000" when x"AA68",
			x"0000" when x"AA69",
			x"0000" when x"AA6A",
			x"0000" when x"AA6B",
			x"0000" when x"AA6C",
			x"0000" when x"AA6D",
			x"0000" when x"AA6E",
			x"0000" when x"AA6F",
			x"0000" when x"AA70",
			x"0000" when x"AA71",
			x"0000" when x"AA72",
			x"0000" when x"AA73",
			x"0000" when x"AA74",
			x"0000" when x"AA75",
			x"0000" when x"AA76",
			x"0000" when x"AA77",
			x"0000" when x"AA78",
			x"0000" when x"AA79",
			x"0000" when x"AA7A",
			x"0000" when x"AA7B",
			x"0000" when x"AA7C",
			x"0000" when x"AA7D",
			x"0000" when x"AA7E",
			x"0000" when x"AA7F",
			x"0000" when x"AA80",
			x"0000" when x"AA81",
			x"0000" when x"AA82",
			x"0000" when x"AA83",
			x"0000" when x"AA84",
			x"0000" when x"AA85",
			x"0000" when x"AA86",
			x"0000" when x"AA87",
			x"0000" when x"AA88",
			x"0000" when x"AA89",
			x"0000" when x"AA8A",
			x"0000" when x"AA8B",
			x"0000" when x"AA8C",
			x"0000" when x"AA8D",
			x"0000" when x"AA8E",
			x"0000" when x"AA8F",
			x"0000" when x"AA90",
			x"0000" when x"AA91",
			x"0000" when x"AA92",
			x"0000" when x"AA93",
			x"0000" when x"AA94",
			x"0000" when x"AA95",
			x"0000" when x"AA96",
			x"0000" when x"AA97",
			x"0000" when x"AA98",
			x"0000" when x"AA99",
			x"0000" when x"AA9A",
			x"0000" when x"AA9B",
			x"0000" when x"AA9C",
			x"0000" when x"AA9D",
			x"0000" when x"AA9E",
			x"0000" when x"AA9F",
			x"0000" when x"AAA0",
			x"0000" when x"AAA1",
			x"0000" when x"AAA2",
			x"0000" when x"AAA3",
			x"0000" when x"AAA4",
			x"0000" when x"AAA5",
			x"0000" when x"AAA6",
			x"0000" when x"AAA7",
			x"0000" when x"AAA8",
			x"0000" when x"AAA9",
			x"0000" when x"AAAA",
			x"0000" when x"AAAB",
			x"0000" when x"AAAC",
			x"0000" when x"AAAD",
			x"0000" when x"AAAE",
			x"0000" when x"AAAF",
			x"0000" when x"AAB0",
			x"0000" when x"AAB1",
			x"0000" when x"AAB2",
			x"0000" when x"AAB3",
			x"0000" when x"AAB4",
			x"0000" when x"AAB5",
			x"0000" when x"AAB6",
			x"0000" when x"AAB7",
			x"0000" when x"AAB8",
			x"0000" when x"AAB9",
			x"0000" when x"AABA",
			x"0000" when x"AABB",
			x"0000" when x"AABC",
			x"0000" when x"AABD",
			x"0000" when x"AABE",
			x"0000" when x"AABF",
			x"0000" when x"AAC0",
			x"0000" when x"AAC1",
			x"0000" when x"AAC2",
			x"0000" when x"AAC3",
			x"0000" when x"AAC4",
			x"0000" when x"AAC5",
			x"0000" when x"AAC6",
			x"0000" when x"AAC7",
			x"0000" when x"AAC8",
			x"0000" when x"AAC9",
			x"0000" when x"AACA",
			x"0000" when x"AACB",
			x"0000" when x"AACC",
			x"0000" when x"AACD",
			x"0000" when x"AACE",
			x"0000" when x"AACF",
			x"0000" when x"AAD0",
			x"0000" when x"AAD1",
			x"0000" when x"AAD2",
			x"0000" when x"AAD3",
			x"0000" when x"AAD4",
			x"0000" when x"AAD5",
			x"0000" when x"AAD6",
			x"0000" when x"AAD7",
			x"0000" when x"AAD8",
			x"0000" when x"AAD9",
			x"0000" when x"AADA",
			x"0000" when x"AADB",
			x"0000" when x"AADC",
			x"0000" when x"AADD",
			x"0000" when x"AADE",
			x"0000" when x"AADF",
			x"0000" when x"AAE0",
			x"0000" when x"AAE1",
			x"0000" when x"AAE2",
			x"0000" when x"AAE3",
			x"0000" when x"AAE4",
			x"0000" when x"AAE5",
			x"0000" when x"AAE6",
			x"0000" when x"AAE7",
			x"0000" when x"AAE8",
			x"0000" when x"AAE9",
			x"0000" when x"AAEA",
			x"0000" when x"AAEB",
			x"0000" when x"AAEC",
			x"0000" when x"AAED",
			x"0000" when x"AAEE",
			x"0000" when x"AAEF",
			x"0000" when x"AAF0",
			x"0000" when x"AAF1",
			x"0000" when x"AAF2",
			x"0000" when x"AAF3",
			x"0000" when x"AAF4",
			x"0000" when x"AAF5",
			x"0000" when x"AAF6",
			x"0000" when x"AAF7",
			x"0000" when x"AAF8",
			x"0000" when x"AAF9",
			x"0000" when x"AAFA",
			x"0000" when x"AAFB",
			x"0000" when x"AAFC",
			x"0000" when x"AAFD",
			x"0000" when x"AAFE",
			x"0000" when x"AAFF",
			x"0000" when x"AB00",
			x"0000" when x"AB01",
			x"0000" when x"AB02",
			x"0000" when x"AB03",
			x"0000" when x"AB04",
			x"0000" when x"AB05",
			x"0000" when x"AB06",
			x"0000" when x"AB07",
			x"0000" when x"AB08",
			x"0000" when x"AB09",
			x"0000" when x"AB0A",
			x"0000" when x"AB0B",
			x"0000" when x"AB0C",
			x"0000" when x"AB0D",
			x"0000" when x"AB0E",
			x"0000" when x"AB0F",
			x"0000" when x"AB10",
			x"0000" when x"AB11",
			x"0000" when x"AB12",
			x"0000" when x"AB13",
			x"0000" when x"AB14",
			x"0000" when x"AB15",
			x"0000" when x"AB16",
			x"0000" when x"AB17",
			x"0000" when x"AB18",
			x"0000" when x"AB19",
			x"0000" when x"AB1A",
			x"0000" when x"AB1B",
			x"0000" when x"AB1C",
			x"0000" when x"AB1D",
			x"0000" when x"AB1E",
			x"0000" when x"AB1F",
			x"0000" when x"AB20",
			x"0000" when x"AB21",
			x"0000" when x"AB22",
			x"0000" when x"AB23",
			x"0000" when x"AB24",
			x"0000" when x"AB25",
			x"0000" when x"AB26",
			x"0000" when x"AB27",
			x"0000" when x"AB28",
			x"0000" when x"AB29",
			x"0000" when x"AB2A",
			x"0000" when x"AB2B",
			x"0000" when x"AB2C",
			x"0000" when x"AB2D",
			x"0000" when x"AB2E",
			x"0000" when x"AB2F",
			x"0000" when x"AB30",
			x"0000" when x"AB31",
			x"0000" when x"AB32",
			x"0000" when x"AB33",
			x"0000" when x"AB34",
			x"0000" when x"AB35",
			x"0000" when x"AB36",
			x"0000" when x"AB37",
			x"0000" when x"AB38",
			x"0000" when x"AB39",
			x"0000" when x"AB3A",
			x"0000" when x"AB3B",
			x"0000" when x"AB3C",
			x"0000" when x"AB3D",
			x"0000" when x"AB3E",
			x"0000" when x"AB3F",
			x"0000" when x"AB40",
			x"0000" when x"AB41",
			x"0000" when x"AB42",
			x"0000" when x"AB43",
			x"0000" when x"AB44",
			x"0000" when x"AB45",
			x"0000" when x"AB46",
			x"0000" when x"AB47",
			x"0000" when x"AB48",
			x"0000" when x"AB49",
			x"0000" when x"AB4A",
			x"0000" when x"AB4B",
			x"0000" when x"AB4C",
			x"0000" when x"AB4D",
			x"0000" when x"AB4E",
			x"0000" when x"AB4F",
			x"0000" when x"AB50",
			x"0000" when x"AB51",
			x"0000" when x"AB52",
			x"0000" when x"AB53",
			x"0000" when x"AB54",
			x"0000" when x"AB55",
			x"0000" when x"AB56",
			x"0000" when x"AB57",
			x"0000" when x"AB58",
			x"0000" when x"AB59",
			x"0000" when x"AB5A",
			x"0000" when x"AB5B",
			x"0000" when x"AB5C",
			x"0000" when x"AB5D",
			x"0000" when x"AB5E",
			x"0000" when x"AB5F",
			x"0000" when x"AB60",
			x"0000" when x"AB61",
			x"0000" when x"AB62",
			x"0000" when x"AB63",
			x"0000" when x"AB64",
			x"0000" when x"AB65",
			x"0000" when x"AB66",
			x"0000" when x"AB67",
			x"0000" when x"AB68",
			x"0000" when x"AB69",
			x"0000" when x"AB6A",
			x"0000" when x"AB6B",
			x"0000" when x"AB6C",
			x"0000" when x"AB6D",
			x"0000" when x"AB6E",
			x"0000" when x"AB6F",
			x"0000" when x"AB70",
			x"0000" when x"AB71",
			x"0000" when x"AB72",
			x"0000" when x"AB73",
			x"0000" when x"AB74",
			x"0000" when x"AB75",
			x"0000" when x"AB76",
			x"0000" when x"AB77",
			x"0000" when x"AB78",
			x"0000" when x"AB79",
			x"0000" when x"AB7A",
			x"0000" when x"AB7B",
			x"0000" when x"AB7C",
			x"0000" when x"AB7D",
			x"0000" when x"AB7E",
			x"0000" when x"AB7F",
			x"0000" when x"AB80",
			x"0000" when x"AB81",
			x"0000" when x"AB82",
			x"0000" when x"AB83",
			x"0000" when x"AB84",
			x"0000" when x"AB85",
			x"0000" when x"AB86",
			x"0000" when x"AB87",
			x"0000" when x"AB88",
			x"0000" when x"AB89",
			x"0000" when x"AB8A",
			x"0000" when x"AB8B",
			x"0000" when x"AB8C",
			x"0000" when x"AB8D",
			x"0000" when x"AB8E",
			x"0000" when x"AB8F",
			x"0000" when x"AB90",
			x"0000" when x"AB91",
			x"0000" when x"AB92",
			x"0000" when x"AB93",
			x"0000" when x"AB94",
			x"0000" when x"AB95",
			x"0000" when x"AB96",
			x"0000" when x"AB97",
			x"0000" when x"AB98",
			x"0000" when x"AB99",
			x"0000" when x"AB9A",
			x"0000" when x"AB9B",
			x"0000" when x"AB9C",
			x"0000" when x"AB9D",
			x"0000" when x"AB9E",
			x"0000" when x"AB9F",
			x"0000" when x"ABA0",
			x"0000" when x"ABA1",
			x"0000" when x"ABA2",
			x"0000" when x"ABA3",
			x"0000" when x"ABA4",
			x"0000" when x"ABA5",
			x"0000" when x"ABA6",
			x"0000" when x"ABA7",
			x"0000" when x"ABA8",
			x"0000" when x"ABA9",
			x"0000" when x"ABAA",
			x"0000" when x"ABAB",
			x"0000" when x"ABAC",
			x"0000" when x"ABAD",
			x"0000" when x"ABAE",
			x"0000" when x"ABAF",
			x"0000" when x"ABB0",
			x"0000" when x"ABB1",
			x"0000" when x"ABB2",
			x"0000" when x"ABB3",
			x"0000" when x"ABB4",
			x"0000" when x"ABB5",
			x"0000" when x"ABB6",
			x"0000" when x"ABB7",
			x"0000" when x"ABB8",
			x"0000" when x"ABB9",
			x"0000" when x"ABBA",
			x"0000" when x"ABBB",
			x"0000" when x"ABBC",
			x"0000" when x"ABBD",
			x"0000" when x"ABBE",
			x"0000" when x"ABBF",
			x"0000" when x"ABC0",
			x"0000" when x"ABC1",
			x"0000" when x"ABC2",
			x"0000" when x"ABC3",
			x"0000" when x"ABC4",
			x"0000" when x"ABC5",
			x"0000" when x"ABC6",
			x"0000" when x"ABC7",
			x"0000" when x"ABC8",
			x"0000" when x"ABC9",
			x"0000" when x"ABCA",
			x"0000" when x"ABCB",
			x"0000" when x"ABCC",
			x"0000" when x"ABCD",
			x"0000" when x"ABCE",
			x"0000" when x"ABCF",
			x"0000" when x"ABD0",
			x"0000" when x"ABD1",
			x"0000" when x"ABD2",
			x"0000" when x"ABD3",
			x"0000" when x"ABD4",
			x"0000" when x"ABD5",
			x"0000" when x"ABD6",
			x"0000" when x"ABD7",
			x"0000" when x"ABD8",
			x"0000" when x"ABD9",
			x"0000" when x"ABDA",
			x"0000" when x"ABDB",
			x"0000" when x"ABDC",
			x"0000" when x"ABDD",
			x"0000" when x"ABDE",
			x"0000" when x"ABDF",
			x"0000" when x"ABE0",
			x"0000" when x"ABE1",
			x"0000" when x"ABE2",
			x"0000" when x"ABE3",
			x"0000" when x"ABE4",
			x"0000" when x"ABE5",
			x"0000" when x"ABE6",
			x"0000" when x"ABE7",
			x"0000" when x"ABE8",
			x"0000" when x"ABE9",
			x"0000" when x"ABEA",
			x"0000" when x"ABEB",
			x"0000" when x"ABEC",
			x"0000" when x"ABED",
			x"0000" when x"ABEE",
			x"0000" when x"ABEF",
			x"0000" when x"ABF0",
			x"0000" when x"ABF1",
			x"0000" when x"ABF2",
			x"0000" when x"ABF3",
			x"0000" when x"ABF4",
			x"0000" when x"ABF5",
			x"0000" when x"ABF6",
			x"0000" when x"ABF7",
			x"0000" when x"ABF8",
			x"0000" when x"ABF9",
			x"0000" when x"ABFA",
			x"0000" when x"ABFB",
			x"0000" when x"ABFC",
			x"0000" when x"ABFD",
			x"0000" when x"ABFE",
			x"0000" when x"ABFF",
			x"0000" when x"AC00",
			x"0000" when x"AC01",
			x"0000" when x"AC02",
			x"0000" when x"AC03",
			x"0000" when x"AC04",
			x"0000" when x"AC05",
			x"0000" when x"AC06",
			x"0000" when x"AC07",
			x"0000" when x"AC08",
			x"0000" when x"AC09",
			x"0000" when x"AC0A",
			x"0000" when x"AC0B",
			x"0000" when x"AC0C",
			x"0000" when x"AC0D",
			x"0000" when x"AC0E",
			x"0000" when x"AC0F",
			x"0000" when x"AC10",
			x"0000" when x"AC11",
			x"0000" when x"AC12",
			x"0000" when x"AC13",
			x"0000" when x"AC14",
			x"0000" when x"AC15",
			x"0000" when x"AC16",
			x"0000" when x"AC17",
			x"0000" when x"AC18",
			x"0000" when x"AC19",
			x"0000" when x"AC1A",
			x"0000" when x"AC1B",
			x"0000" when x"AC1C",
			x"0000" when x"AC1D",
			x"0000" when x"AC1E",
			x"0000" when x"AC1F",
			x"0000" when x"AC20",
			x"0000" when x"AC21",
			x"0000" when x"AC22",
			x"0000" when x"AC23",
			x"0000" when x"AC24",
			x"0000" when x"AC25",
			x"0000" when x"AC26",
			x"0000" when x"AC27",
			x"0000" when x"AC28",
			x"0000" when x"AC29",
			x"0000" when x"AC2A",
			x"0000" when x"AC2B",
			x"0000" when x"AC2C",
			x"0000" when x"AC2D",
			x"0000" when x"AC2E",
			x"0000" when x"AC2F",
			x"0000" when x"AC30",
			x"0000" when x"AC31",
			x"0000" when x"AC32",
			x"0000" when x"AC33",
			x"0000" when x"AC34",
			x"0000" when x"AC35",
			x"0000" when x"AC36",
			x"0000" when x"AC37",
			x"0000" when x"AC38",
			x"0000" when x"AC39",
			x"0000" when x"AC3A",
			x"0000" when x"AC3B",
			x"0000" when x"AC3C",
			x"0000" when x"AC3D",
			x"0000" when x"AC3E",
			x"0000" when x"AC3F",
			x"0000" when x"AC40",
			x"0000" when x"AC41",
			x"0000" when x"AC42",
			x"0000" when x"AC43",
			x"0000" when x"AC44",
			x"0000" when x"AC45",
			x"0000" when x"AC46",
			x"0000" when x"AC47",
			x"0000" when x"AC48",
			x"0000" when x"AC49",
			x"0000" when x"AC4A",
			x"0000" when x"AC4B",
			x"0000" when x"AC4C",
			x"0000" when x"AC4D",
			x"0000" when x"AC4E",
			x"0000" when x"AC4F",
			x"0000" when x"AC50",
			x"0000" when x"AC51",
			x"0000" when x"AC52",
			x"0000" when x"AC53",
			x"0000" when x"AC54",
			x"0000" when x"AC55",
			x"0000" when x"AC56",
			x"0000" when x"AC57",
			x"0000" when x"AC58",
			x"0000" when x"AC59",
			x"0000" when x"AC5A",
			x"0000" when x"AC5B",
			x"0000" when x"AC5C",
			x"0000" when x"AC5D",
			x"0000" when x"AC5E",
			x"0000" when x"AC5F",
			x"0000" when x"AC60",
			x"0000" when x"AC61",
			x"0000" when x"AC62",
			x"0000" when x"AC63",
			x"0000" when x"AC64",
			x"0000" when x"AC65",
			x"0000" when x"AC66",
			x"0000" when x"AC67",
			x"0000" when x"AC68",
			x"0000" when x"AC69",
			x"0000" when x"AC6A",
			x"0000" when x"AC6B",
			x"0000" when x"AC6C",
			x"0000" when x"AC6D",
			x"0000" when x"AC6E",
			x"0000" when x"AC6F",
			x"0000" when x"AC70",
			x"0000" when x"AC71",
			x"0000" when x"AC72",
			x"0000" when x"AC73",
			x"0000" when x"AC74",
			x"0000" when x"AC75",
			x"0000" when x"AC76",
			x"0000" when x"AC77",
			x"0000" when x"AC78",
			x"0000" when x"AC79",
			x"0000" when x"AC7A",
			x"0000" when x"AC7B",
			x"0000" when x"AC7C",
			x"0000" when x"AC7D",
			x"0000" when x"AC7E",
			x"0000" when x"AC7F",
			x"0000" when x"AC80",
			x"0000" when x"AC81",
			x"0000" when x"AC82",
			x"0000" when x"AC83",
			x"0000" when x"AC84",
			x"0000" when x"AC85",
			x"0000" when x"AC86",
			x"0000" when x"AC87",
			x"0000" when x"AC88",
			x"0000" when x"AC89",
			x"0000" when x"AC8A",
			x"0000" when x"AC8B",
			x"0000" when x"AC8C",
			x"0000" when x"AC8D",
			x"0000" when x"AC8E",
			x"0000" when x"AC8F",
			x"0000" when x"AC90",
			x"0000" when x"AC91",
			x"0000" when x"AC92",
			x"0000" when x"AC93",
			x"0000" when x"AC94",
			x"0000" when x"AC95",
			x"0000" when x"AC96",
			x"0000" when x"AC97",
			x"0000" when x"AC98",
			x"0000" when x"AC99",
			x"0000" when x"AC9A",
			x"0000" when x"AC9B",
			x"0000" when x"AC9C",
			x"0000" when x"AC9D",
			x"0000" when x"AC9E",
			x"0000" when x"AC9F",
			x"0000" when x"ACA0",
			x"0000" when x"ACA1",
			x"0000" when x"ACA2",
			x"0000" when x"ACA3",
			x"0000" when x"ACA4",
			x"0000" when x"ACA5",
			x"0000" when x"ACA6",
			x"0000" when x"ACA7",
			x"0000" when x"ACA8",
			x"0000" when x"ACA9",
			x"0000" when x"ACAA",
			x"0000" when x"ACAB",
			x"0000" when x"ACAC",
			x"0000" when x"ACAD",
			x"0000" when x"ACAE",
			x"0000" when x"ACAF",
			x"0000" when x"ACB0",
			x"0000" when x"ACB1",
			x"0000" when x"ACB2",
			x"0000" when x"ACB3",
			x"0000" when x"ACB4",
			x"0000" when x"ACB5",
			x"0000" when x"ACB6",
			x"0000" when x"ACB7",
			x"0000" when x"ACB8",
			x"0000" when x"ACB9",
			x"0000" when x"ACBA",
			x"0000" when x"ACBB",
			x"0000" when x"ACBC",
			x"0000" when x"ACBD",
			x"0000" when x"ACBE",
			x"0000" when x"ACBF",
			x"0000" when x"ACC0",
			x"0000" when x"ACC1",
			x"0000" when x"ACC2",
			x"0000" when x"ACC3",
			x"0000" when x"ACC4",
			x"0000" when x"ACC5",
			x"0000" when x"ACC6",
			x"0000" when x"ACC7",
			x"0000" when x"ACC8",
			x"0000" when x"ACC9",
			x"0000" when x"ACCA",
			x"0000" when x"ACCB",
			x"0000" when x"ACCC",
			x"0000" when x"ACCD",
			x"0000" when x"ACCE",
			x"0000" when x"ACCF",
			x"0000" when x"ACD0",
			x"0000" when x"ACD1",
			x"0000" when x"ACD2",
			x"0000" when x"ACD3",
			x"0000" when x"ACD4",
			x"0000" when x"ACD5",
			x"0000" when x"ACD6",
			x"0000" when x"ACD7",
			x"0000" when x"ACD8",
			x"0000" when x"ACD9",
			x"0000" when x"ACDA",
			x"0000" when x"ACDB",
			x"0000" when x"ACDC",
			x"0000" when x"ACDD",
			x"0000" when x"ACDE",
			x"0000" when x"ACDF",
			x"0000" when x"ACE0",
			x"0000" when x"ACE1",
			x"0000" when x"ACE2",
			x"0000" when x"ACE3",
			x"0000" when x"ACE4",
			x"0000" when x"ACE5",
			x"0000" when x"ACE6",
			x"0000" when x"ACE7",
			x"0000" when x"ACE8",
			x"0000" when x"ACE9",
			x"0000" when x"ACEA",
			x"0000" when x"ACEB",
			x"0000" when x"ACEC",
			x"0000" when x"ACED",
			x"0000" when x"ACEE",
			x"0000" when x"ACEF",
			x"0000" when x"ACF0",
			x"0000" when x"ACF1",
			x"0000" when x"ACF2",
			x"0000" when x"ACF3",
			x"0000" when x"ACF4",
			x"0000" when x"ACF5",
			x"0000" when x"ACF6",
			x"0000" when x"ACF7",
			x"0000" when x"ACF8",
			x"0000" when x"ACF9",
			x"0000" when x"ACFA",
			x"0000" when x"ACFB",
			x"0000" when x"ACFC",
			x"0000" when x"ACFD",
			x"0000" when x"ACFE",
			x"0000" when x"ACFF",
			x"0000" when x"AD00",
			x"0000" when x"AD01",
			x"0000" when x"AD02",
			x"0000" when x"AD03",
			x"0000" when x"AD04",
			x"0000" when x"AD05",
			x"0000" when x"AD06",
			x"0000" when x"AD07",
			x"0000" when x"AD08",
			x"0000" when x"AD09",
			x"0000" when x"AD0A",
			x"0000" when x"AD0B",
			x"0000" when x"AD0C",
			x"0000" when x"AD0D",
			x"0000" when x"AD0E",
			x"0000" when x"AD0F",
			x"0000" when x"AD10",
			x"0000" when x"AD11",
			x"0000" when x"AD12",
			x"0000" when x"AD13",
			x"0000" when x"AD14",
			x"0000" when x"AD15",
			x"0000" when x"AD16",
			x"0000" when x"AD17",
			x"0000" when x"AD18",
			x"0000" when x"AD19",
			x"0000" when x"AD1A",
			x"0000" when x"AD1B",
			x"0000" when x"AD1C",
			x"0000" when x"AD1D",
			x"0000" when x"AD1E",
			x"0000" when x"AD1F",
			x"0000" when x"AD20",
			x"0000" when x"AD21",
			x"0000" when x"AD22",
			x"0000" when x"AD23",
			x"0000" when x"AD24",
			x"0000" when x"AD25",
			x"0000" when x"AD26",
			x"0000" when x"AD27",
			x"0000" when x"AD28",
			x"0000" when x"AD29",
			x"0000" when x"AD2A",
			x"0000" when x"AD2B",
			x"0000" when x"AD2C",
			x"0000" when x"AD2D",
			x"0000" when x"AD2E",
			x"0000" when x"AD2F",
			x"0000" when x"AD30",
			x"0000" when x"AD31",
			x"0000" when x"AD32",
			x"0000" when x"AD33",
			x"0000" when x"AD34",
			x"0000" when x"AD35",
			x"0000" when x"AD36",
			x"0000" when x"AD37",
			x"0000" when x"AD38",
			x"0000" when x"AD39",
			x"0000" when x"AD3A",
			x"0000" when x"AD3B",
			x"0000" when x"AD3C",
			x"0000" when x"AD3D",
			x"0000" when x"AD3E",
			x"0000" when x"AD3F",
			x"0000" when x"AD40",
			x"0000" when x"AD41",
			x"0000" when x"AD42",
			x"0000" when x"AD43",
			x"0000" when x"AD44",
			x"0000" when x"AD45",
			x"0000" when x"AD46",
			x"0000" when x"AD47",
			x"0000" when x"AD48",
			x"0000" when x"AD49",
			x"0000" when x"AD4A",
			x"0000" when x"AD4B",
			x"0000" when x"AD4C",
			x"0000" when x"AD4D",
			x"0000" when x"AD4E",
			x"0000" when x"AD4F",
			x"0000" when x"AD50",
			x"0000" when x"AD51",
			x"0000" when x"AD52",
			x"0000" when x"AD53",
			x"0000" when x"AD54",
			x"0000" when x"AD55",
			x"0000" when x"AD56",
			x"0000" when x"AD57",
			x"0000" when x"AD58",
			x"0000" when x"AD59",
			x"0000" when x"AD5A",
			x"0000" when x"AD5B",
			x"0000" when x"AD5C",
			x"0000" when x"AD5D",
			x"0000" when x"AD5E",
			x"0000" when x"AD5F",
			x"0000" when x"AD60",
			x"0000" when x"AD61",
			x"0000" when x"AD62",
			x"0000" when x"AD63",
			x"0000" when x"AD64",
			x"0000" when x"AD65",
			x"0000" when x"AD66",
			x"0000" when x"AD67",
			x"0000" when x"AD68",
			x"0000" when x"AD69",
			x"0000" when x"AD6A",
			x"0000" when x"AD6B",
			x"0000" when x"AD6C",
			x"0000" when x"AD6D",
			x"0000" when x"AD6E",
			x"0000" when x"AD6F",
			x"0000" when x"AD70",
			x"0000" when x"AD71",
			x"0000" when x"AD72",
			x"0000" when x"AD73",
			x"0000" when x"AD74",
			x"0000" when x"AD75",
			x"0000" when x"AD76",
			x"0000" when x"AD77",
			x"0000" when x"AD78",
			x"0000" when x"AD79",
			x"0000" when x"AD7A",
			x"0000" when x"AD7B",
			x"0000" when x"AD7C",
			x"0000" when x"AD7D",
			x"0000" when x"AD7E",
			x"0000" when x"AD7F",
			x"0000" when x"AD80",
			x"0000" when x"AD81",
			x"0000" when x"AD82",
			x"0000" when x"AD83",
			x"0000" when x"AD84",
			x"0000" when x"AD85",
			x"0000" when x"AD86",
			x"0000" when x"AD87",
			x"0000" when x"AD88",
			x"0000" when x"AD89",
			x"0000" when x"AD8A",
			x"0000" when x"AD8B",
			x"0000" when x"AD8C",
			x"0000" when x"AD8D",
			x"0000" when x"AD8E",
			x"0000" when x"AD8F",
			x"0000" when x"AD90",
			x"0000" when x"AD91",
			x"0000" when x"AD92",
			x"0000" when x"AD93",
			x"0000" when x"AD94",
			x"0000" when x"AD95",
			x"0000" when x"AD96",
			x"0000" when x"AD97",
			x"0000" when x"AD98",
			x"0000" when x"AD99",
			x"0000" when x"AD9A",
			x"0000" when x"AD9B",
			x"0000" when x"AD9C",
			x"0000" when x"AD9D",
			x"0000" when x"AD9E",
			x"0000" when x"AD9F",
			x"0000" when x"ADA0",
			x"0000" when x"ADA1",
			x"0000" when x"ADA2",
			x"0000" when x"ADA3",
			x"0000" when x"ADA4",
			x"0000" when x"ADA5",
			x"0000" when x"ADA6",
			x"0000" when x"ADA7",
			x"0000" when x"ADA8",
			x"0000" when x"ADA9",
			x"0000" when x"ADAA",
			x"0000" when x"ADAB",
			x"0000" when x"ADAC",
			x"0000" when x"ADAD",
			x"0000" when x"ADAE",
			x"0000" when x"ADAF",
			x"0000" when x"ADB0",
			x"0000" when x"ADB1",
			x"0000" when x"ADB2",
			x"0000" when x"ADB3",
			x"0000" when x"ADB4",
			x"0000" when x"ADB5",
			x"0000" when x"ADB6",
			x"0000" when x"ADB7",
			x"0000" when x"ADB8",
			x"0000" when x"ADB9",
			x"0000" when x"ADBA",
			x"0000" when x"ADBB",
			x"0000" when x"ADBC",
			x"0000" when x"ADBD",
			x"0000" when x"ADBE",
			x"0000" when x"ADBF",
			x"0000" when x"ADC0",
			x"0000" when x"ADC1",
			x"0000" when x"ADC2",
			x"0000" when x"ADC3",
			x"0000" when x"ADC4",
			x"0000" when x"ADC5",
			x"0000" when x"ADC6",
			x"0000" when x"ADC7",
			x"0000" when x"ADC8",
			x"0000" when x"ADC9",
			x"0000" when x"ADCA",
			x"0000" when x"ADCB",
			x"0000" when x"ADCC",
			x"0000" when x"ADCD",
			x"0000" when x"ADCE",
			x"0000" when x"ADCF",
			x"0000" when x"ADD0",
			x"0000" when x"ADD1",
			x"0000" when x"ADD2",
			x"0000" when x"ADD3",
			x"0000" when x"ADD4",
			x"0000" when x"ADD5",
			x"0000" when x"ADD6",
			x"0000" when x"ADD7",
			x"0000" when x"ADD8",
			x"0000" when x"ADD9",
			x"0000" when x"ADDA",
			x"0000" when x"ADDB",
			x"0000" when x"ADDC",
			x"0000" when x"ADDD",
			x"0000" when x"ADDE",
			x"0000" when x"ADDF",
			x"0000" when x"ADE0",
			x"0000" when x"ADE1",
			x"0000" when x"ADE2",
			x"0000" when x"ADE3",
			x"0000" when x"ADE4",
			x"0000" when x"ADE5",
			x"0000" when x"ADE6",
			x"0000" when x"ADE7",
			x"0000" when x"ADE8",
			x"0000" when x"ADE9",
			x"0000" when x"ADEA",
			x"0000" when x"ADEB",
			x"0000" when x"ADEC",
			x"0000" when x"ADED",
			x"0000" when x"ADEE",
			x"0000" when x"ADEF",
			x"0000" when x"ADF0",
			x"0000" when x"ADF1",
			x"0000" when x"ADF2",
			x"0000" when x"ADF3",
			x"0000" when x"ADF4",
			x"0000" when x"ADF5",
			x"0000" when x"ADF6",
			x"0000" when x"ADF7",
			x"0000" when x"ADF8",
			x"0000" when x"ADF9",
			x"0000" when x"ADFA",
			x"0000" when x"ADFB",
			x"0000" when x"ADFC",
			x"0000" when x"ADFD",
			x"0000" when x"ADFE",
			x"0000" when x"ADFF",
			x"0000" when x"AE00",
			x"0000" when x"AE01",
			x"0000" when x"AE02",
			x"0000" when x"AE03",
			x"0000" when x"AE04",
			x"0000" when x"AE05",
			x"0000" when x"AE06",
			x"0000" when x"AE07",
			x"0000" when x"AE08",
			x"0000" when x"AE09",
			x"0000" when x"AE0A",
			x"0000" when x"AE0B",
			x"0000" when x"AE0C",
			x"0000" when x"AE0D",
			x"0000" when x"AE0E",
			x"0000" when x"AE0F",
			x"0000" when x"AE10",
			x"0000" when x"AE11",
			x"0000" when x"AE12",
			x"0000" when x"AE13",
			x"0000" when x"AE14",
			x"0000" when x"AE15",
			x"0000" when x"AE16",
			x"0000" when x"AE17",
			x"0000" when x"AE18",
			x"0000" when x"AE19",
			x"0000" when x"AE1A",
			x"0000" when x"AE1B",
			x"0000" when x"AE1C",
			x"0000" when x"AE1D",
			x"0000" when x"AE1E",
			x"0000" when x"AE1F",
			x"0000" when x"AE20",
			x"0000" when x"AE21",
			x"0000" when x"AE22",
			x"0000" when x"AE23",
			x"0000" when x"AE24",
			x"0000" when x"AE25",
			x"0000" when x"AE26",
			x"0000" when x"AE27",
			x"0000" when x"AE28",
			x"0000" when x"AE29",
			x"0000" when x"AE2A",
			x"0000" when x"AE2B",
			x"0000" when x"AE2C",
			x"0000" when x"AE2D",
			x"0000" when x"AE2E",
			x"0000" when x"AE2F",
			x"0000" when x"AE30",
			x"0000" when x"AE31",
			x"0000" when x"AE32",
			x"0000" when x"AE33",
			x"0000" when x"AE34",
			x"0000" when x"AE35",
			x"0000" when x"AE36",
			x"0000" when x"AE37",
			x"0000" when x"AE38",
			x"0000" when x"AE39",
			x"0000" when x"AE3A",
			x"0000" when x"AE3B",
			x"0000" when x"AE3C",
			x"0000" when x"AE3D",
			x"0000" when x"AE3E",
			x"0000" when x"AE3F",
			x"0000" when x"AE40",
			x"0000" when x"AE41",
			x"0000" when x"AE42",
			x"0000" when x"AE43",
			x"0000" when x"AE44",
			x"0000" when x"AE45",
			x"0000" when x"AE46",
			x"0000" when x"AE47",
			x"0000" when x"AE48",
			x"0000" when x"AE49",
			x"0000" when x"AE4A",
			x"0000" when x"AE4B",
			x"0000" when x"AE4C",
			x"0000" when x"AE4D",
			x"0000" when x"AE4E",
			x"0000" when x"AE4F",
			x"0000" when x"AE50",
			x"0000" when x"AE51",
			x"0000" when x"AE52",
			x"0000" when x"AE53",
			x"0000" when x"AE54",
			x"0000" when x"AE55",
			x"0000" when x"AE56",
			x"0000" when x"AE57",
			x"0000" when x"AE58",
			x"0000" when x"AE59",
			x"0000" when x"AE5A",
			x"0000" when x"AE5B",
			x"0000" when x"AE5C",
			x"0000" when x"AE5D",
			x"0000" when x"AE5E",
			x"0000" when x"AE5F",
			x"0000" when x"AE60",
			x"0000" when x"AE61",
			x"0000" when x"AE62",
			x"0000" when x"AE63",
			x"0000" when x"AE64",
			x"0000" when x"AE65",
			x"0000" when x"AE66",
			x"0000" when x"AE67",
			x"0000" when x"AE68",
			x"0000" when x"AE69",
			x"0000" when x"AE6A",
			x"0000" when x"AE6B",
			x"0000" when x"AE6C",
			x"0000" when x"AE6D",
			x"0000" when x"AE6E",
			x"0000" when x"AE6F",
			x"0000" when x"AE70",
			x"0000" when x"AE71",
			x"0000" when x"AE72",
			x"0000" when x"AE73",
			x"0000" when x"AE74",
			x"0000" when x"AE75",
			x"0000" when x"AE76",
			x"0000" when x"AE77",
			x"0000" when x"AE78",
			x"0000" when x"AE79",
			x"0000" when x"AE7A",
			x"0000" when x"AE7B",
			x"0000" when x"AE7C",
			x"0000" when x"AE7D",
			x"0000" when x"AE7E",
			x"0000" when x"AE7F",
			x"0000" when x"AE80",
			x"0000" when x"AE81",
			x"0000" when x"AE82",
			x"0000" when x"AE83",
			x"0000" when x"AE84",
			x"0000" when x"AE85",
			x"0000" when x"AE86",
			x"0000" when x"AE87",
			x"0000" when x"AE88",
			x"0000" when x"AE89",
			x"0000" when x"AE8A",
			x"0000" when x"AE8B",
			x"0000" when x"AE8C",
			x"0000" when x"AE8D",
			x"0000" when x"AE8E",
			x"0000" when x"AE8F",
			x"0000" when x"AE90",
			x"0000" when x"AE91",
			x"0000" when x"AE92",
			x"0000" when x"AE93",
			x"0000" when x"AE94",
			x"0000" when x"AE95",
			x"0000" when x"AE96",
			x"0000" when x"AE97",
			x"0000" when x"AE98",
			x"0000" when x"AE99",
			x"0000" when x"AE9A",
			x"0000" when x"AE9B",
			x"0000" when x"AE9C",
			x"0000" when x"AE9D",
			x"0000" when x"AE9E",
			x"0000" when x"AE9F",
			x"0000" when x"AEA0",
			x"0000" when x"AEA1",
			x"0000" when x"AEA2",
			x"0000" when x"AEA3",
			x"0000" when x"AEA4",
			x"0000" when x"AEA5",
			x"0000" when x"AEA6",
			x"0000" when x"AEA7",
			x"0000" when x"AEA8",
			x"0000" when x"AEA9",
			x"0000" when x"AEAA",
			x"0000" when x"AEAB",
			x"0000" when x"AEAC",
			x"0000" when x"AEAD",
			x"0000" when x"AEAE",
			x"0000" when x"AEAF",
			x"0000" when x"AEB0",
			x"0000" when x"AEB1",
			x"0000" when x"AEB2",
			x"0000" when x"AEB3",
			x"0000" when x"AEB4",
			x"0000" when x"AEB5",
			x"0000" when x"AEB6",
			x"0000" when x"AEB7",
			x"0000" when x"AEB8",
			x"0000" when x"AEB9",
			x"0000" when x"AEBA",
			x"0000" when x"AEBB",
			x"0000" when x"AEBC",
			x"0000" when x"AEBD",
			x"0000" when x"AEBE",
			x"0000" when x"AEBF",
			x"0000" when x"AEC0",
			x"0000" when x"AEC1",
			x"0000" when x"AEC2",
			x"0000" when x"AEC3",
			x"0000" when x"AEC4",
			x"0000" when x"AEC5",
			x"0000" when x"AEC6",
			x"0000" when x"AEC7",
			x"0000" when x"AEC8",
			x"0000" when x"AEC9",
			x"0000" when x"AECA",
			x"0000" when x"AECB",
			x"0000" when x"AECC",
			x"0000" when x"AECD",
			x"0000" when x"AECE",
			x"0000" when x"AECF",
			x"0000" when x"AED0",
			x"0000" when x"AED1",
			x"0000" when x"AED2",
			x"0000" when x"AED3",
			x"0000" when x"AED4",
			x"0000" when x"AED5",
			x"0000" when x"AED6",
			x"0000" when x"AED7",
			x"0000" when x"AED8",
			x"0000" when x"AED9",
			x"0000" when x"AEDA",
			x"0000" when x"AEDB",
			x"0000" when x"AEDC",
			x"0000" when x"AEDD",
			x"0000" when x"AEDE",
			x"0000" when x"AEDF",
			x"0000" when x"AEE0",
			x"0000" when x"AEE1",
			x"0000" when x"AEE2",
			x"0000" when x"AEE3",
			x"0000" when x"AEE4",
			x"0000" when x"AEE5",
			x"0000" when x"AEE6",
			x"0000" when x"AEE7",
			x"0000" when x"AEE8",
			x"0000" when x"AEE9",
			x"0000" when x"AEEA",
			x"0000" when x"AEEB",
			x"0000" when x"AEEC",
			x"0000" when x"AEED",
			x"0000" when x"AEEE",
			x"0000" when x"AEEF",
			x"0000" when x"AEF0",
			x"0000" when x"AEF1",
			x"0000" when x"AEF2",
			x"0000" when x"AEF3",
			x"0000" when x"AEF4",
			x"0000" when x"AEF5",
			x"0000" when x"AEF6",
			x"0000" when x"AEF7",
			x"0000" when x"AEF8",
			x"0000" when x"AEF9",
			x"0000" when x"AEFA",
			x"0000" when x"AEFB",
			x"0000" when x"AEFC",
			x"0000" when x"AEFD",
			x"0000" when x"AEFE",
			x"0000" when x"AEFF",
			x"0000" when x"AF00",
			x"0000" when x"AF01",
			x"0000" when x"AF02",
			x"0000" when x"AF03",
			x"0000" when x"AF04",
			x"0000" when x"AF05",
			x"0000" when x"AF06",
			x"0000" when x"AF07",
			x"0000" when x"AF08",
			x"0000" when x"AF09",
			x"0000" when x"AF0A",
			x"0000" when x"AF0B",
			x"0000" when x"AF0C",
			x"0000" when x"AF0D",
			x"0000" when x"AF0E",
			x"0000" when x"AF0F",
			x"0000" when x"AF10",
			x"0000" when x"AF11",
			x"0000" when x"AF12",
			x"0000" when x"AF13",
			x"0000" when x"AF14",
			x"0000" when x"AF15",
			x"0000" when x"AF16",
			x"0000" when x"AF17",
			x"0000" when x"AF18",
			x"0000" when x"AF19",
			x"0000" when x"AF1A",
			x"0000" when x"AF1B",
			x"0000" when x"AF1C",
			x"0000" when x"AF1D",
			x"0000" when x"AF1E",
			x"0000" when x"AF1F",
			x"0000" when x"AF20",
			x"0000" when x"AF21",
			x"0000" when x"AF22",
			x"0000" when x"AF23",
			x"0000" when x"AF24",
			x"0000" when x"AF25",
			x"0000" when x"AF26",
			x"0000" when x"AF27",
			x"0000" when x"AF28",
			x"0000" when x"AF29",
			x"0000" when x"AF2A",
			x"0000" when x"AF2B",
			x"0000" when x"AF2C",
			x"0000" when x"AF2D",
			x"0000" when x"AF2E",
			x"0000" when x"AF2F",
			x"0000" when x"AF30",
			x"0000" when x"AF31",
			x"0000" when x"AF32",
			x"0000" when x"AF33",
			x"0000" when x"AF34",
			x"0000" when x"AF35",
			x"0000" when x"AF36",
			x"0000" when x"AF37",
			x"0000" when x"AF38",
			x"0000" when x"AF39",
			x"0000" when x"AF3A",
			x"0000" when x"AF3B",
			x"0000" when x"AF3C",
			x"0000" when x"AF3D",
			x"0000" when x"AF3E",
			x"0000" when x"AF3F",
			x"0000" when x"AF40",
			x"0000" when x"AF41",
			x"0000" when x"AF42",
			x"0000" when x"AF43",
			x"0000" when x"AF44",
			x"0000" when x"AF45",
			x"0000" when x"AF46",
			x"0000" when x"AF47",
			x"0000" when x"AF48",
			x"0000" when x"AF49",
			x"0000" when x"AF4A",
			x"0000" when x"AF4B",
			x"0000" when x"AF4C",
			x"0000" when x"AF4D",
			x"0000" when x"AF4E",
			x"0000" when x"AF4F",
			x"0000" when x"AF50",
			x"0000" when x"AF51",
			x"0000" when x"AF52",
			x"0000" when x"AF53",
			x"0000" when x"AF54",
			x"0000" when x"AF55",
			x"0000" when x"AF56",
			x"0000" when x"AF57",
			x"0000" when x"AF58",
			x"0000" when x"AF59",
			x"0000" when x"AF5A",
			x"0000" when x"AF5B",
			x"0000" when x"AF5C",
			x"0000" when x"AF5D",
			x"0000" when x"AF5E",
			x"0000" when x"AF5F",
			x"0000" when x"AF60",
			x"0000" when x"AF61",
			x"0000" when x"AF62",
			x"0000" when x"AF63",
			x"0000" when x"AF64",
			x"0000" when x"AF65",
			x"0000" when x"AF66",
			x"0000" when x"AF67",
			x"0000" when x"AF68",
			x"0000" when x"AF69",
			x"0000" when x"AF6A",
			x"0000" when x"AF6B",
			x"0000" when x"AF6C",
			x"0000" when x"AF6D",
			x"0000" when x"AF6E",
			x"0000" when x"AF6F",
			x"0000" when x"AF70",
			x"0000" when x"AF71",
			x"0000" when x"AF72",
			x"0000" when x"AF73",
			x"0000" when x"AF74",
			x"0000" when x"AF75",
			x"0000" when x"AF76",
			x"0000" when x"AF77",
			x"0000" when x"AF78",
			x"0000" when x"AF79",
			x"0000" when x"AF7A",
			x"0000" when x"AF7B",
			x"0000" when x"AF7C",
			x"0000" when x"AF7D",
			x"0000" when x"AF7E",
			x"0000" when x"AF7F",
			x"0000" when x"AF80",
			x"0000" when x"AF81",
			x"0000" when x"AF82",
			x"0000" when x"AF83",
			x"0000" when x"AF84",
			x"0000" when x"AF85",
			x"0000" when x"AF86",
			x"0000" when x"AF87",
			x"0000" when x"AF88",
			x"0000" when x"AF89",
			x"0000" when x"AF8A",
			x"0000" when x"AF8B",
			x"0000" when x"AF8C",
			x"0000" when x"AF8D",
			x"0000" when x"AF8E",
			x"0000" when x"AF8F",
			x"0000" when x"AF90",
			x"0000" when x"AF91",
			x"0000" when x"AF92",
			x"0000" when x"AF93",
			x"0000" when x"AF94",
			x"0000" when x"AF95",
			x"0000" when x"AF96",
			x"0000" when x"AF97",
			x"0000" when x"AF98",
			x"0000" when x"AF99",
			x"0000" when x"AF9A",
			x"0000" when x"AF9B",
			x"0000" when x"AF9C",
			x"0000" when x"AF9D",
			x"0000" when x"AF9E",
			x"0000" when x"AF9F",
			x"0000" when x"AFA0",
			x"0000" when x"AFA1",
			x"0000" when x"AFA2",
			x"0000" when x"AFA3",
			x"0000" when x"AFA4",
			x"0000" when x"AFA5",
			x"0000" when x"AFA6",
			x"0000" when x"AFA7",
			x"0000" when x"AFA8",
			x"0000" when x"AFA9",
			x"0000" when x"AFAA",
			x"0000" when x"AFAB",
			x"0000" when x"AFAC",
			x"0000" when x"AFAD",
			x"0000" when x"AFAE",
			x"0000" when x"AFAF",
			x"0000" when x"AFB0",
			x"0000" when x"AFB1",
			x"0000" when x"AFB2",
			x"0000" when x"AFB3",
			x"0000" when x"AFB4",
			x"0000" when x"AFB5",
			x"0000" when x"AFB6",
			x"0000" when x"AFB7",
			x"0000" when x"AFB8",
			x"0000" when x"AFB9",
			x"0000" when x"AFBA",
			x"0000" when x"AFBB",
			x"0000" when x"AFBC",
			x"0000" when x"AFBD",
			x"0000" when x"AFBE",
			x"0000" when x"AFBF",
			x"0000" when x"AFC0",
			x"0000" when x"AFC1",
			x"0000" when x"AFC2",
			x"0000" when x"AFC3",
			x"0000" when x"AFC4",
			x"0000" when x"AFC5",
			x"0000" when x"AFC6",
			x"0000" when x"AFC7",
			x"0000" when x"AFC8",
			x"0000" when x"AFC9",
			x"0000" when x"AFCA",
			x"0000" when x"AFCB",
			x"0000" when x"AFCC",
			x"0000" when x"AFCD",
			x"0000" when x"AFCE",
			x"0000" when x"AFCF",
			x"0000" when x"AFD0",
			x"0000" when x"AFD1",
			x"0000" when x"AFD2",
			x"0000" when x"AFD3",
			x"0000" when x"AFD4",
			x"0000" when x"AFD5",
			x"0000" when x"AFD6",
			x"0000" when x"AFD7",
			x"0000" when x"AFD8",
			x"0000" when x"AFD9",
			x"0000" when x"AFDA",
			x"0000" when x"AFDB",
			x"0000" when x"AFDC",
			x"0000" when x"AFDD",
			x"0000" when x"AFDE",
			x"0000" when x"AFDF",
			x"0000" when x"AFE0",
			x"0000" when x"AFE1",
			x"0000" when x"AFE2",
			x"0000" when x"AFE3",
			x"0000" when x"AFE4",
			x"0000" when x"AFE5",
			x"0000" when x"AFE6",
			x"0000" when x"AFE7",
			x"0000" when x"AFE8",
			x"0000" when x"AFE9",
			x"0000" when x"AFEA",
			x"0000" when x"AFEB",
			x"0000" when x"AFEC",
			x"0000" when x"AFED",
			x"0000" when x"AFEE",
			x"0000" when x"AFEF",
			x"0000" when x"AFF0",
			x"0000" when x"AFF1",
			x"0000" when x"AFF2",
			x"0000" when x"AFF3",
			x"0000" when x"AFF4",
			x"0000" when x"AFF5",
			x"0000" when x"AFF6",
			x"0000" when x"AFF7",
			x"0000" when x"AFF8",
			x"0000" when x"AFF9",
			x"0000" when x"AFFA",
			x"0000" when x"AFFB",
			x"0000" when x"AFFC",
			x"0000" when x"AFFD",
			x"0000" when x"AFFE",
			x"0000" when x"AFFF",
			x"0000" when x"B000",
			x"0000" when x"B001",
			x"0000" when x"B002",
			x"0000" when x"B003",
			x"0000" when x"B004",
			x"0000" when x"B005",
			x"0000" when x"B006",
			x"0000" when x"B007",
			x"0000" when x"B008",
			x"0000" when x"B009",
			x"0000" when x"B00A",
			x"0000" when x"B00B",
			x"0000" when x"B00C",
			x"0000" when x"B00D",
			x"0000" when x"B00E",
			x"0000" when x"B00F",
			x"0000" when x"B010",
			x"0000" when x"B011",
			x"0000" when x"B012",
			x"0000" when x"B013",
			x"0000" when x"B014",
			x"0000" when x"B015",
			x"0000" when x"B016",
			x"0000" when x"B017",
			x"0000" when x"B018",
			x"0000" when x"B019",
			x"0000" when x"B01A",
			x"0000" when x"B01B",
			x"0000" when x"B01C",
			x"0000" when x"B01D",
			x"0000" when x"B01E",
			x"0000" when x"B01F",
			x"0000" when x"B020",
			x"0000" when x"B021",
			x"0000" when x"B022",
			x"0000" when x"B023",
			x"0000" when x"B024",
			x"0000" when x"B025",
			x"0000" when x"B026",
			x"0000" when x"B027",
			x"0000" when x"B028",
			x"0000" when x"B029",
			x"0000" when x"B02A",
			x"0000" when x"B02B",
			x"0000" when x"B02C",
			x"0000" when x"B02D",
			x"0000" when x"B02E",
			x"0000" when x"B02F",
			x"0000" when x"B030",
			x"0000" when x"B031",
			x"0000" when x"B032",
			x"0000" when x"B033",
			x"0000" when x"B034",
			x"0000" when x"B035",
			x"0000" when x"B036",
			x"0000" when x"B037",
			x"0000" when x"B038",
			x"0000" when x"B039",
			x"0000" when x"B03A",
			x"0000" when x"B03B",
			x"0000" when x"B03C",
			x"0000" when x"B03D",
			x"0000" when x"B03E",
			x"0000" when x"B03F",
			x"0000" when x"B040",
			x"0000" when x"B041",
			x"0000" when x"B042",
			x"0000" when x"B043",
			x"0000" when x"B044",
			x"0000" when x"B045",
			x"0000" when x"B046",
			x"0000" when x"B047",
			x"0000" when x"B048",
			x"0000" when x"B049",
			x"0000" when x"B04A",
			x"0000" when x"B04B",
			x"0000" when x"B04C",
			x"0000" when x"B04D",
			x"0000" when x"B04E",
			x"0000" when x"B04F",
			x"0000" when x"B050",
			x"0000" when x"B051",
			x"0000" when x"B052",
			x"0000" when x"B053",
			x"0000" when x"B054",
			x"0000" when x"B055",
			x"0000" when x"B056",
			x"0000" when x"B057",
			x"0000" when x"B058",
			x"0000" when x"B059",
			x"0000" when x"B05A",
			x"0000" when x"B05B",
			x"0000" when x"B05C",
			x"0000" when x"B05D",
			x"0000" when x"B05E",
			x"0000" when x"B05F",
			x"0000" when x"B060",
			x"0000" when x"B061",
			x"0000" when x"B062",
			x"0000" when x"B063",
			x"0000" when x"B064",
			x"0000" when x"B065",
			x"0000" when x"B066",
			x"0000" when x"B067",
			x"0000" when x"B068",
			x"0000" when x"B069",
			x"0000" when x"B06A",
			x"0000" when x"B06B",
			x"0000" when x"B06C",
			x"0000" when x"B06D",
			x"0000" when x"B06E",
			x"0000" when x"B06F",
			x"0000" when x"B070",
			x"0000" when x"B071",
			x"0000" when x"B072",
			x"0000" when x"B073",
			x"0000" when x"B074",
			x"0000" when x"B075",
			x"0000" when x"B076",
			x"0000" when x"B077",
			x"0000" when x"B078",
			x"0000" when x"B079",
			x"0000" when x"B07A",
			x"0000" when x"B07B",
			x"0000" when x"B07C",
			x"0000" when x"B07D",
			x"0000" when x"B07E",
			x"0000" when x"B07F",
			x"0000" when x"B080",
			x"0000" when x"B081",
			x"0000" when x"B082",
			x"0000" when x"B083",
			x"0000" when x"B084",
			x"0000" when x"B085",
			x"0000" when x"B086",
			x"0000" when x"B087",
			x"0000" when x"B088",
			x"0000" when x"B089",
			x"0000" when x"B08A",
			x"0000" when x"B08B",
			x"0000" when x"B08C",
			x"0000" when x"B08D",
			x"0000" when x"B08E",
			x"0000" when x"B08F",
			x"0000" when x"B090",
			x"0000" when x"B091",
			x"0000" when x"B092",
			x"0000" when x"B093",
			x"0000" when x"B094",
			x"0000" when x"B095",
			x"0000" when x"B096",
			x"0000" when x"B097",
			x"0000" when x"B098",
			x"0000" when x"B099",
			x"0000" when x"B09A",
			x"0000" when x"B09B",
			x"0000" when x"B09C",
			x"0000" when x"B09D",
			x"0000" when x"B09E",
			x"0000" when x"B09F",
			x"0000" when x"B0A0",
			x"0000" when x"B0A1",
			x"0000" when x"B0A2",
			x"0000" when x"B0A3",
			x"0000" when x"B0A4",
			x"0000" when x"B0A5",
			x"0000" when x"B0A6",
			x"0000" when x"B0A7",
			x"0000" when x"B0A8",
			x"0000" when x"B0A9",
			x"0000" when x"B0AA",
			x"0000" when x"B0AB",
			x"0000" when x"B0AC",
			x"0000" when x"B0AD",
			x"0000" when x"B0AE",
			x"0000" when x"B0AF",
			x"0000" when x"B0B0",
			x"0000" when x"B0B1",
			x"0000" when x"B0B2",
			x"0000" when x"B0B3",
			x"0000" when x"B0B4",
			x"0000" when x"B0B5",
			x"0000" when x"B0B6",
			x"0000" when x"B0B7",
			x"0000" when x"B0B8",
			x"0000" when x"B0B9",
			x"0000" when x"B0BA",
			x"0000" when x"B0BB",
			x"0000" when x"B0BC",
			x"0000" when x"B0BD",
			x"0000" when x"B0BE",
			x"0000" when x"B0BF",
			x"0000" when x"B0C0",
			x"0000" when x"B0C1",
			x"0000" when x"B0C2",
			x"0000" when x"B0C3",
			x"0000" when x"B0C4",
			x"0000" when x"B0C5",
			x"0000" when x"B0C6",
			x"0000" when x"B0C7",
			x"0000" when x"B0C8",
			x"0000" when x"B0C9",
			x"0000" when x"B0CA",
			x"0000" when x"B0CB",
			x"0000" when x"B0CC",
			x"0000" when x"B0CD",
			x"0000" when x"B0CE",
			x"0000" when x"B0CF",
			x"0000" when x"B0D0",
			x"0000" when x"B0D1",
			x"0000" when x"B0D2",
			x"0000" when x"B0D3",
			x"0000" when x"B0D4",
			x"0000" when x"B0D5",
			x"0000" when x"B0D6",
			x"0000" when x"B0D7",
			x"0000" when x"B0D8",
			x"0000" when x"B0D9",
			x"0000" when x"B0DA",
			x"0000" when x"B0DB",
			x"0000" when x"B0DC",
			x"0000" when x"B0DD",
			x"0000" when x"B0DE",
			x"0000" when x"B0DF",
			x"0000" when x"B0E0",
			x"0000" when x"B0E1",
			x"0000" when x"B0E2",
			x"0000" when x"B0E3",
			x"0000" when x"B0E4",
			x"0000" when x"B0E5",
			x"0000" when x"B0E6",
			x"0000" when x"B0E7",
			x"0000" when x"B0E8",
			x"0000" when x"B0E9",
			x"0000" when x"B0EA",
			x"0000" when x"B0EB",
			x"0000" when x"B0EC",
			x"0000" when x"B0ED",
			x"0000" when x"B0EE",
			x"0000" when x"B0EF",
			x"0000" when x"B0F0",
			x"0000" when x"B0F1",
			x"0000" when x"B0F2",
			x"0000" when x"B0F3",
			x"0000" when x"B0F4",
			x"0000" when x"B0F5",
			x"0000" when x"B0F6",
			x"0000" when x"B0F7",
			x"0000" when x"B0F8",
			x"0000" when x"B0F9",
			x"0000" when x"B0FA",
			x"0000" when x"B0FB",
			x"0000" when x"B0FC",
			x"0000" when x"B0FD",
			x"0000" when x"B0FE",
			x"0000" when x"B0FF",
			x"0000" when x"B100",
			x"0000" when x"B101",
			x"0000" when x"B102",
			x"0000" when x"B103",
			x"0000" when x"B104",
			x"0000" when x"B105",
			x"0000" when x"B106",
			x"0000" when x"B107",
			x"0000" when x"B108",
			x"0000" when x"B109",
			x"0000" when x"B10A",
			x"0000" when x"B10B",
			x"0000" when x"B10C",
			x"0000" when x"B10D",
			x"0000" when x"B10E",
			x"0000" when x"B10F",
			x"0000" when x"B110",
			x"0000" when x"B111",
			x"0000" when x"B112",
			x"0000" when x"B113",
			x"0000" when x"B114",
			x"0000" when x"B115",
			x"0000" when x"B116",
			x"0000" when x"B117",
			x"0000" when x"B118",
			x"0000" when x"B119",
			x"0000" when x"B11A",
			x"0000" when x"B11B",
			x"0000" when x"B11C",
			x"0000" when x"B11D",
			x"0000" when x"B11E",
			x"0000" when x"B11F",
			x"0000" when x"B120",
			x"0000" when x"B121",
			x"0000" when x"B122",
			x"0000" when x"B123",
			x"0000" when x"B124",
			x"0000" when x"B125",
			x"0000" when x"B126",
			x"0000" when x"B127",
			x"0000" when x"B128",
			x"0000" when x"B129",
			x"0000" when x"B12A",
			x"0000" when x"B12B",
			x"0000" when x"B12C",
			x"0000" when x"B12D",
			x"0000" when x"B12E",
			x"0000" when x"B12F",
			x"0000" when x"B130",
			x"0000" when x"B131",
			x"0000" when x"B132",
			x"0000" when x"B133",
			x"0000" when x"B134",
			x"0000" when x"B135",
			x"0000" when x"B136",
			x"0000" when x"B137",
			x"0000" when x"B138",
			x"0000" when x"B139",
			x"0000" when x"B13A",
			x"0000" when x"B13B",
			x"0000" when x"B13C",
			x"0000" when x"B13D",
			x"0000" when x"B13E",
			x"0000" when x"B13F",
			x"0000" when x"B140",
			x"0000" when x"B141",
			x"0000" when x"B142",
			x"0000" when x"B143",
			x"0000" when x"B144",
			x"0000" when x"B145",
			x"0000" when x"B146",
			x"0000" when x"B147",
			x"0000" when x"B148",
			x"0000" when x"B149",
			x"0000" when x"B14A",
			x"0000" when x"B14B",
			x"0000" when x"B14C",
			x"0000" when x"B14D",
			x"0000" when x"B14E",
			x"0000" when x"B14F",
			x"0000" when x"B150",
			x"0000" when x"B151",
			x"0000" when x"B152",
			x"0000" when x"B153",
			x"0000" when x"B154",
			x"0000" when x"B155",
			x"0000" when x"B156",
			x"0000" when x"B157",
			x"0000" when x"B158",
			x"0000" when x"B159",
			x"0000" when x"B15A",
			x"0000" when x"B15B",
			x"0000" when x"B15C",
			x"0000" when x"B15D",
			x"0000" when x"B15E",
			x"0000" when x"B15F",
			x"0000" when x"B160",
			x"0000" when x"B161",
			x"0000" when x"B162",
			x"0000" when x"B163",
			x"0000" when x"B164",
			x"0000" when x"B165",
			x"0000" when x"B166",
			x"0000" when x"B167",
			x"0000" when x"B168",
			x"0000" when x"B169",
			x"0000" when x"B16A",
			x"0000" when x"B16B",
			x"0000" when x"B16C",
			x"0000" when x"B16D",
			x"0000" when x"B16E",
			x"0000" when x"B16F",
			x"0000" when x"B170",
			x"0000" when x"B171",
			x"0000" when x"B172",
			x"0000" when x"B173",
			x"0000" when x"B174",
			x"0000" when x"B175",
			x"0000" when x"B176",
			x"0000" when x"B177",
			x"0000" when x"B178",
			x"0000" when x"B179",
			x"0000" when x"B17A",
			x"0000" when x"B17B",
			x"0000" when x"B17C",
			x"0000" when x"B17D",
			x"0000" when x"B17E",
			x"0000" when x"B17F",
			x"0000" when x"B180",
			x"0000" when x"B181",
			x"0000" when x"B182",
			x"0000" when x"B183",
			x"0000" when x"B184",
			x"0000" when x"B185",
			x"0000" when x"B186",
			x"0000" when x"B187",
			x"0000" when x"B188",
			x"0000" when x"B189",
			x"0000" when x"B18A",
			x"0000" when x"B18B",
			x"0000" when x"B18C",
			x"0000" when x"B18D",
			x"0000" when x"B18E",
			x"0000" when x"B18F",
			x"0000" when x"B190",
			x"0000" when x"B191",
			x"0000" when x"B192",
			x"0000" when x"B193",
			x"0000" when x"B194",
			x"0000" when x"B195",
			x"0000" when x"B196",
			x"0000" when x"B197",
			x"0000" when x"B198",
			x"0000" when x"B199",
			x"0000" when x"B19A",
			x"0000" when x"B19B",
			x"0000" when x"B19C",
			x"0000" when x"B19D",
			x"0000" when x"B19E",
			x"0000" when x"B19F",
			x"0000" when x"B1A0",
			x"0000" when x"B1A1",
			x"0000" when x"B1A2",
			x"0000" when x"B1A3",
			x"0000" when x"B1A4",
			x"0000" when x"B1A5",
			x"0000" when x"B1A6",
			x"0000" when x"B1A7",
			x"0000" when x"B1A8",
			x"0000" when x"B1A9",
			x"0000" when x"B1AA",
			x"0000" when x"B1AB",
			x"0000" when x"B1AC",
			x"0000" when x"B1AD",
			x"0000" when x"B1AE",
			x"0000" when x"B1AF",
			x"0000" when x"B1B0",
			x"0000" when x"B1B1",
			x"0000" when x"B1B2",
			x"0000" when x"B1B3",
			x"0000" when x"B1B4",
			x"0000" when x"B1B5",
			x"0000" when x"B1B6",
			x"0000" when x"B1B7",
			x"0000" when x"B1B8",
			x"0000" when x"B1B9",
			x"0000" when x"B1BA",
			x"0000" when x"B1BB",
			x"0000" when x"B1BC",
			x"0000" when x"B1BD",
			x"0000" when x"B1BE",
			x"0000" when x"B1BF",
			x"0000" when x"B1C0",
			x"0000" when x"B1C1",
			x"0000" when x"B1C2",
			x"0000" when x"B1C3",
			x"0000" when x"B1C4",
			x"0000" when x"B1C5",
			x"0000" when x"B1C6",
			x"0000" when x"B1C7",
			x"0000" when x"B1C8",
			x"0000" when x"B1C9",
			x"0000" when x"B1CA",
			x"0000" when x"B1CB",
			x"0000" when x"B1CC",
			x"0000" when x"B1CD",
			x"0000" when x"B1CE",
			x"0000" when x"B1CF",
			x"0000" when x"B1D0",
			x"0000" when x"B1D1",
			x"0000" when x"B1D2",
			x"0000" when x"B1D3",
			x"0000" when x"B1D4",
			x"0000" when x"B1D5",
			x"0000" when x"B1D6",
			x"0000" when x"B1D7",
			x"0000" when x"B1D8",
			x"0000" when x"B1D9",
			x"0000" when x"B1DA",
			x"0000" when x"B1DB",
			x"0000" when x"B1DC",
			x"0000" when x"B1DD",
			x"0000" when x"B1DE",
			x"0000" when x"B1DF",
			x"0000" when x"B1E0",
			x"0000" when x"B1E1",
			x"0000" when x"B1E2",
			x"0000" when x"B1E3",
			x"0000" when x"B1E4",
			x"0000" when x"B1E5",
			x"0000" when x"B1E6",
			x"0000" when x"B1E7",
			x"0000" when x"B1E8",
			x"0000" when x"B1E9",
			x"0000" when x"B1EA",
			x"0000" when x"B1EB",
			x"0000" when x"B1EC",
			x"0000" when x"B1ED",
			x"0000" when x"B1EE",
			x"0000" when x"B1EF",
			x"0000" when x"B1F0",
			x"0000" when x"B1F1",
			x"0000" when x"B1F2",
			x"0000" when x"B1F3",
			x"0000" when x"B1F4",
			x"0000" when x"B1F5",
			x"0000" when x"B1F6",
			x"0000" when x"B1F7",
			x"0000" when x"B1F8",
			x"0000" when x"B1F9",
			x"0000" when x"B1FA",
			x"0000" when x"B1FB",
			x"0000" when x"B1FC",
			x"0000" when x"B1FD",
			x"0000" when x"B1FE",
			x"0000" when x"B1FF",
			x"0000" when x"B200",
			x"0000" when x"B201",
			x"0000" when x"B202",
			x"0000" when x"B203",
			x"0000" when x"B204",
			x"0000" when x"B205",
			x"0000" when x"B206",
			x"0000" when x"B207",
			x"0000" when x"B208",
			x"0000" when x"B209",
			x"0000" when x"B20A",
			x"0000" when x"B20B",
			x"0000" when x"B20C",
			x"0000" when x"B20D",
			x"0000" when x"B20E",
			x"0000" when x"B20F",
			x"0000" when x"B210",
			x"0000" when x"B211",
			x"0000" when x"B212",
			x"0000" when x"B213",
			x"0000" when x"B214",
			x"0000" when x"B215",
			x"0000" when x"B216",
			x"0000" when x"B217",
			x"0000" when x"B218",
			x"0000" when x"B219",
			x"0000" when x"B21A",
			x"0000" when x"B21B",
			x"0000" when x"B21C",
			x"0000" when x"B21D",
			x"0000" when x"B21E",
			x"0000" when x"B21F",
			x"0000" when x"B220",
			x"0000" when x"B221",
			x"0000" when x"B222",
			x"0000" when x"B223",
			x"0000" when x"B224",
			x"0000" when x"B225",
			x"0000" when x"B226",
			x"0000" when x"B227",
			x"0000" when x"B228",
			x"0000" when x"B229",
			x"0000" when x"B22A",
			x"0000" when x"B22B",
			x"0000" when x"B22C",
			x"0000" when x"B22D",
			x"0000" when x"B22E",
			x"0000" when x"B22F",
			x"0000" when x"B230",
			x"0000" when x"B231",
			x"0000" when x"B232",
			x"0000" when x"B233",
			x"0000" when x"B234",
			x"0000" when x"B235",
			x"0000" when x"B236",
			x"0000" when x"B237",
			x"0000" when x"B238",
			x"0000" when x"B239",
			x"0000" when x"B23A",
			x"0000" when x"B23B",
			x"0000" when x"B23C",
			x"0000" when x"B23D",
			x"0000" when x"B23E",
			x"0000" when x"B23F",
			x"0000" when x"B240",
			x"0000" when x"B241",
			x"0000" when x"B242",
			x"0000" when x"B243",
			x"0000" when x"B244",
			x"0000" when x"B245",
			x"0000" when x"B246",
			x"0000" when x"B247",
			x"0000" when x"B248",
			x"0000" when x"B249",
			x"0000" when x"B24A",
			x"0000" when x"B24B",
			x"0000" when x"B24C",
			x"0000" when x"B24D",
			x"0000" when x"B24E",
			x"0000" when x"B24F",
			x"0000" when x"B250",
			x"0000" when x"B251",
			x"0000" when x"B252",
			x"0000" when x"B253",
			x"0000" when x"B254",
			x"0000" when x"B255",
			x"0000" when x"B256",
			x"0000" when x"B257",
			x"0000" when x"B258",
			x"0000" when x"B259",
			x"0000" when x"B25A",
			x"0000" when x"B25B",
			x"0000" when x"B25C",
			x"0000" when x"B25D",
			x"0000" when x"B25E",
			x"0000" when x"B25F",
			x"0000" when x"B260",
			x"0000" when x"B261",
			x"0000" when x"B262",
			x"0000" when x"B263",
			x"0000" when x"B264",
			x"0000" when x"B265",
			x"0000" when x"B266",
			x"0000" when x"B267",
			x"0000" when x"B268",
			x"0000" when x"B269",
			x"0000" when x"B26A",
			x"0000" when x"B26B",
			x"0000" when x"B26C",
			x"0000" when x"B26D",
			x"0000" when x"B26E",
			x"0000" when x"B26F",
			x"0000" when x"B270",
			x"0000" when x"B271",
			x"0000" when x"B272",
			x"0000" when x"B273",
			x"0000" when x"B274",
			x"0000" when x"B275",
			x"0000" when x"B276",
			x"0000" when x"B277",
			x"0000" when x"B278",
			x"0000" when x"B279",
			x"0000" when x"B27A",
			x"0000" when x"B27B",
			x"0000" when x"B27C",
			x"0000" when x"B27D",
			x"0000" when x"B27E",
			x"0000" when x"B27F",
			x"0000" when x"B280",
			x"0000" when x"B281",
			x"0000" when x"B282",
			x"0000" when x"B283",
			x"0000" when x"B284",
			x"0000" when x"B285",
			x"0000" when x"B286",
			x"0000" when x"B287",
			x"0000" when x"B288",
			x"0000" when x"B289",
			x"0000" when x"B28A",
			x"0000" when x"B28B",
			x"0000" when x"B28C",
			x"0000" when x"B28D",
			x"0000" when x"B28E",
			x"0000" when x"B28F",
			x"0000" when x"B290",
			x"0000" when x"B291",
			x"0000" when x"B292",
			x"0000" when x"B293",
			x"0000" when x"B294",
			x"0000" when x"B295",
			x"0000" when x"B296",
			x"0000" when x"B297",
			x"0000" when x"B298",
			x"0000" when x"B299",
			x"0000" when x"B29A",
			x"0000" when x"B29B",
			x"0000" when x"B29C",
			x"0000" when x"B29D",
			x"0000" when x"B29E",
			x"0000" when x"B29F",
			x"0000" when x"B2A0",
			x"0000" when x"B2A1",
			x"0000" when x"B2A2",
			x"0000" when x"B2A3",
			x"0000" when x"B2A4",
			x"0000" when x"B2A5",
			x"0000" when x"B2A6",
			x"0000" when x"B2A7",
			x"0000" when x"B2A8",
			x"0000" when x"B2A9",
			x"0000" when x"B2AA",
			x"0000" when x"B2AB",
			x"0000" when x"B2AC",
			x"0000" when x"B2AD",
			x"0000" when x"B2AE",
			x"0000" when x"B2AF",
			x"0000" when x"B2B0",
			x"0000" when x"B2B1",
			x"0000" when x"B2B2",
			x"0000" when x"B2B3",
			x"0000" when x"B2B4",
			x"0000" when x"B2B5",
			x"0000" when x"B2B6",
			x"0000" when x"B2B7",
			x"0000" when x"B2B8",
			x"0000" when x"B2B9",
			x"0000" when x"B2BA",
			x"0000" when x"B2BB",
			x"0000" when x"B2BC",
			x"0000" when x"B2BD",
			x"0000" when x"B2BE",
			x"0000" when x"B2BF",
			x"0000" when x"B2C0",
			x"0000" when x"B2C1",
			x"0000" when x"B2C2",
			x"0000" when x"B2C3",
			x"0000" when x"B2C4",
			x"0000" when x"B2C5",
			x"0000" when x"B2C6",
			x"0000" when x"B2C7",
			x"0000" when x"B2C8",
			x"0000" when x"B2C9",
			x"0000" when x"B2CA",
			x"0000" when x"B2CB",
			x"0000" when x"B2CC",
			x"0000" when x"B2CD",
			x"0000" when x"B2CE",
			x"0000" when x"B2CF",
			x"0000" when x"B2D0",
			x"0000" when x"B2D1",
			x"0000" when x"B2D2",
			x"0000" when x"B2D3",
			x"0000" when x"B2D4",
			x"0000" when x"B2D5",
			x"0000" when x"B2D6",
			x"0000" when x"B2D7",
			x"0000" when x"B2D8",
			x"0000" when x"B2D9",
			x"0000" when x"B2DA",
			x"0000" when x"B2DB",
			x"0000" when x"B2DC",
			x"0000" when x"B2DD",
			x"0000" when x"B2DE",
			x"0000" when x"B2DF",
			x"0000" when x"B2E0",
			x"0000" when x"B2E1",
			x"0000" when x"B2E2",
			x"0000" when x"B2E3",
			x"0000" when x"B2E4",
			x"0000" when x"B2E5",
			x"0000" when x"B2E6",
			x"0000" when x"B2E7",
			x"0000" when x"B2E8",
			x"0000" when x"B2E9",
			x"0000" when x"B2EA",
			x"0000" when x"B2EB",
			x"0000" when x"B2EC",
			x"0000" when x"B2ED",
			x"0000" when x"B2EE",
			x"0000" when x"B2EF",
			x"0000" when x"B2F0",
			x"0000" when x"B2F1",
			x"0000" when x"B2F2",
			x"0000" when x"B2F3",
			x"0000" when x"B2F4",
			x"0000" when x"B2F5",
			x"0000" when x"B2F6",
			x"0000" when x"B2F7",
			x"0000" when x"B2F8",
			x"0000" when x"B2F9",
			x"0000" when x"B2FA",
			x"0000" when x"B2FB",
			x"0000" when x"B2FC",
			x"0000" when x"B2FD",
			x"0000" when x"B2FE",
			x"0000" when x"B2FF",
			x"0000" when x"B300",
			x"0000" when x"B301",
			x"0000" when x"B302",
			x"0000" when x"B303",
			x"0000" when x"B304",
			x"0000" when x"B305",
			x"0000" when x"B306",
			x"0000" when x"B307",
			x"0000" when x"B308",
			x"0000" when x"B309",
			x"0000" when x"B30A",
			x"0000" when x"B30B",
			x"0000" when x"B30C",
			x"0000" when x"B30D",
			x"0000" when x"B30E",
			x"0000" when x"B30F",
			x"0000" when x"B310",
			x"0000" when x"B311",
			x"0000" when x"B312",
			x"0000" when x"B313",
			x"0000" when x"B314",
			x"0000" when x"B315",
			x"0000" when x"B316",
			x"0000" when x"B317",
			x"0000" when x"B318",
			x"0000" when x"B319",
			x"0000" when x"B31A",
			x"0000" when x"B31B",
			x"0000" when x"B31C",
			x"0000" when x"B31D",
			x"0000" when x"B31E",
			x"0000" when x"B31F",
			x"0000" when x"B320",
			x"0000" when x"B321",
			x"0000" when x"B322",
			x"0000" when x"B323",
			x"0000" when x"B324",
			x"0000" when x"B325",
			x"0000" when x"B326",
			x"0000" when x"B327",
			x"0000" when x"B328",
			x"0000" when x"B329",
			x"0000" when x"B32A",
			x"0000" when x"B32B",
			x"0000" when x"B32C",
			x"0000" when x"B32D",
			x"0000" when x"B32E",
			x"0000" when x"B32F",
			x"0000" when x"B330",
			x"0000" when x"B331",
			x"0000" when x"B332",
			x"0000" when x"B333",
			x"0000" when x"B334",
			x"0000" when x"B335",
			x"0000" when x"B336",
			x"0000" when x"B337",
			x"0000" when x"B338",
			x"0000" when x"B339",
			x"0000" when x"B33A",
			x"0000" when x"B33B",
			x"0000" when x"B33C",
			x"0000" when x"B33D",
			x"0000" when x"B33E",
			x"0000" when x"B33F",
			x"0000" when x"B340",
			x"0000" when x"B341",
			x"0000" when x"B342",
			x"0000" when x"B343",
			x"0000" when x"B344",
			x"0000" when x"B345",
			x"0000" when x"B346",
			x"0000" when x"B347",
			x"0000" when x"B348",
			x"0000" when x"B349",
			x"0000" when x"B34A",
			x"0000" when x"B34B",
			x"0000" when x"B34C",
			x"0000" when x"B34D",
			x"0000" when x"B34E",
			x"0000" when x"B34F",
			x"0000" when x"B350",
			x"0000" when x"B351",
			x"0000" when x"B352",
			x"0000" when x"B353",
			x"0000" when x"B354",
			x"0000" when x"B355",
			x"0000" when x"B356",
			x"0000" when x"B357",
			x"0000" when x"B358",
			x"0000" when x"B359",
			x"0000" when x"B35A",
			x"0000" when x"B35B",
			x"0000" when x"B35C",
			x"0000" when x"B35D",
			x"0000" when x"B35E",
			x"0000" when x"B35F",
			x"0000" when x"B360",
			x"0000" when x"B361",
			x"0000" when x"B362",
			x"0000" when x"B363",
			x"0000" when x"B364",
			x"0000" when x"B365",
			x"0000" when x"B366",
			x"0000" when x"B367",
			x"0000" when x"B368",
			x"0000" when x"B369",
			x"0000" when x"B36A",
			x"0000" when x"B36B",
			x"0000" when x"B36C",
			x"0000" when x"B36D",
			x"0000" when x"B36E",
			x"0000" when x"B36F",
			x"0000" when x"B370",
			x"0000" when x"B371",
			x"0000" when x"B372",
			x"0000" when x"B373",
			x"0000" when x"B374",
			x"0000" when x"B375",
			x"0000" when x"B376",
			x"0000" when x"B377",
			x"0000" when x"B378",
			x"0000" when x"B379",
			x"0000" when x"B37A",
			x"0000" when x"B37B",
			x"0000" when x"B37C",
			x"0000" when x"B37D",
			x"0000" when x"B37E",
			x"0000" when x"B37F",
			x"0000" when x"B380",
			x"0000" when x"B381",
			x"0000" when x"B382",
			x"0000" when x"B383",
			x"0000" when x"B384",
			x"0000" when x"B385",
			x"0000" when x"B386",
			x"0000" when x"B387",
			x"0000" when x"B388",
			x"0000" when x"B389",
			x"0000" when x"B38A",
			x"0000" when x"B38B",
			x"0000" when x"B38C",
			x"0000" when x"B38D",
			x"0000" when x"B38E",
			x"0000" when x"B38F",
			x"0000" when x"B390",
			x"0000" when x"B391",
			x"0000" when x"B392",
			x"0000" when x"B393",
			x"0000" when x"B394",
			x"0000" when x"B395",
			x"0000" when x"B396",
			x"0000" when x"B397",
			x"0000" when x"B398",
			x"0000" when x"B399",
			x"0000" when x"B39A",
			x"0000" when x"B39B",
			x"0000" when x"B39C",
			x"0000" when x"B39D",
			x"0000" when x"B39E",
			x"0000" when x"B39F",
			x"0000" when x"B3A0",
			x"0000" when x"B3A1",
			x"0000" when x"B3A2",
			x"0000" when x"B3A3",
			x"0000" when x"B3A4",
			x"0000" when x"B3A5",
			x"0000" when x"B3A6",
			x"0000" when x"B3A7",
			x"0000" when x"B3A8",
			x"0000" when x"B3A9",
			x"0000" when x"B3AA",
			x"0000" when x"B3AB",
			x"0000" when x"B3AC",
			x"0000" when x"B3AD",
			x"0000" when x"B3AE",
			x"0000" when x"B3AF",
			x"0000" when x"B3B0",
			x"0000" when x"B3B1",
			x"0000" when x"B3B2",
			x"0000" when x"B3B3",
			x"0000" when x"B3B4",
			x"0000" when x"B3B5",
			x"0000" when x"B3B6",
			x"0000" when x"B3B7",
			x"0000" when x"B3B8",
			x"0000" when x"B3B9",
			x"0000" when x"B3BA",
			x"0000" when x"B3BB",
			x"0000" when x"B3BC",
			x"0000" when x"B3BD",
			x"0000" when x"B3BE",
			x"0000" when x"B3BF",
			x"0000" when x"B3C0",
			x"0000" when x"B3C1",
			x"0000" when x"B3C2",
			x"0000" when x"B3C3",
			x"0000" when x"B3C4",
			x"0000" when x"B3C5",
			x"0000" when x"B3C6",
			x"0000" when x"B3C7",
			x"0000" when x"B3C8",
			x"0000" when x"B3C9",
			x"0000" when x"B3CA",
			x"0000" when x"B3CB",
			x"0000" when x"B3CC",
			x"0000" when x"B3CD",
			x"0000" when x"B3CE",
			x"0000" when x"B3CF",
			x"0000" when x"B3D0",
			x"0000" when x"B3D1",
			x"0000" when x"B3D2",
			x"0000" when x"B3D3",
			x"0000" when x"B3D4",
			x"0000" when x"B3D5",
			x"0000" when x"B3D6",
			x"0000" when x"B3D7",
			x"0000" when x"B3D8",
			x"0000" when x"B3D9",
			x"0000" when x"B3DA",
			x"0000" when x"B3DB",
			x"0000" when x"B3DC",
			x"0000" when x"B3DD",
			x"0000" when x"B3DE",
			x"0000" when x"B3DF",
			x"0000" when x"B3E0",
			x"0000" when x"B3E1",
			x"0000" when x"B3E2",
			x"0000" when x"B3E3",
			x"0000" when x"B3E4",
			x"0000" when x"B3E5",
			x"0000" when x"B3E6",
			x"0000" when x"B3E7",
			x"0000" when x"B3E8",
			x"0000" when x"B3E9",
			x"0000" when x"B3EA",
			x"0000" when x"B3EB",
			x"0000" when x"B3EC",
			x"0000" when x"B3ED",
			x"0000" when x"B3EE",
			x"0000" when x"B3EF",
			x"0000" when x"B3F0",
			x"0000" when x"B3F1",
			x"0000" when x"B3F2",
			x"0000" when x"B3F3",
			x"0000" when x"B3F4",
			x"0000" when x"B3F5",
			x"0000" when x"B3F6",
			x"0000" when x"B3F7",
			x"0000" when x"B3F8",
			x"0000" when x"B3F9",
			x"0000" when x"B3FA",
			x"0000" when x"B3FB",
			x"0000" when x"B3FC",
			x"0000" when x"B3FD",
			x"0000" when x"B3FE",
			x"0000" when x"B3FF",
			x"0000" when x"B400",
			x"0000" when x"B401",
			x"0000" when x"B402",
			x"0000" when x"B403",
			x"0000" when x"B404",
			x"0000" when x"B405",
			x"0000" when x"B406",
			x"0000" when x"B407",
			x"0000" when x"B408",
			x"0000" when x"B409",
			x"0000" when x"B40A",
			x"0000" when x"B40B",
			x"0000" when x"B40C",
			x"0000" when x"B40D",
			x"0000" when x"B40E",
			x"0000" when x"B40F",
			x"0000" when x"B410",
			x"0000" when x"B411",
			x"0000" when x"B412",
			x"0000" when x"B413",
			x"0000" when x"B414",
			x"0000" when x"B415",
			x"0000" when x"B416",
			x"0000" when x"B417",
			x"0000" when x"B418",
			x"0000" when x"B419",
			x"0000" when x"B41A",
			x"0000" when x"B41B",
			x"0000" when x"B41C",
			x"0000" when x"B41D",
			x"0000" when x"B41E",
			x"0000" when x"B41F",
			x"0000" when x"B420",
			x"0000" when x"B421",
			x"0000" when x"B422",
			x"0000" when x"B423",
			x"0000" when x"B424",
			x"0000" when x"B425",
			x"0000" when x"B426",
			x"0000" when x"B427",
			x"0000" when x"B428",
			x"0000" when x"B429",
			x"0000" when x"B42A",
			x"0000" when x"B42B",
			x"0000" when x"B42C",
			x"0000" when x"B42D",
			x"0000" when x"B42E",
			x"0000" when x"B42F",
			x"0000" when x"B430",
			x"0000" when x"B431",
			x"0000" when x"B432",
			x"0000" when x"B433",
			x"0000" when x"B434",
			x"0000" when x"B435",
			x"0000" when x"B436",
			x"0000" when x"B437",
			x"0000" when x"B438",
			x"0000" when x"B439",
			x"0000" when x"B43A",
			x"0000" when x"B43B",
			x"0000" when x"B43C",
			x"0000" when x"B43D",
			x"0000" when x"B43E",
			x"0000" when x"B43F",
			x"0000" when x"B440",
			x"0000" when x"B441",
			x"0000" when x"B442",
			x"0000" when x"B443",
			x"0000" when x"B444",
			x"0000" when x"B445",
			x"0000" when x"B446",
			x"0000" when x"B447",
			x"0000" when x"B448",
			x"0000" when x"B449",
			x"0000" when x"B44A",
			x"0000" when x"B44B",
			x"0000" when x"B44C",
			x"0000" when x"B44D",
			x"0000" when x"B44E",
			x"0000" when x"B44F",
			x"0000" when x"B450",
			x"0000" when x"B451",
			x"0000" when x"B452",
			x"0000" when x"B453",
			x"0000" when x"B454",
			x"0000" when x"B455",
			x"0000" when x"B456",
			x"0000" when x"B457",
			x"0000" when x"B458",
			x"0000" when x"B459",
			x"0000" when x"B45A",
			x"0000" when x"B45B",
			x"0000" when x"B45C",
			x"0000" when x"B45D",
			x"0000" when x"B45E",
			x"0000" when x"B45F",
			x"0000" when x"B460",
			x"0000" when x"B461",
			x"0000" when x"B462",
			x"0000" when x"B463",
			x"0000" when x"B464",
			x"0000" when x"B465",
			x"0000" when x"B466",
			x"0000" when x"B467",
			x"0000" when x"B468",
			x"0000" when x"B469",
			x"0000" when x"B46A",
			x"0000" when x"B46B",
			x"0000" when x"B46C",
			x"0000" when x"B46D",
			x"0000" when x"B46E",
			x"0000" when x"B46F",
			x"0000" when x"B470",
			x"0000" when x"B471",
			x"0000" when x"B472",
			x"0000" when x"B473",
			x"0000" when x"B474",
			x"0000" when x"B475",
			x"0000" when x"B476",
			x"0000" when x"B477",
			x"0000" when x"B478",
			x"0000" when x"B479",
			x"0000" when x"B47A",
			x"0000" when x"B47B",
			x"0000" when x"B47C",
			x"0000" when x"B47D",
			x"0000" when x"B47E",
			x"0000" when x"B47F",
			x"0000" when x"B480",
			x"0000" when x"B481",
			x"0000" when x"B482",
			x"0000" when x"B483",
			x"0000" when x"B484",
			x"0000" when x"B485",
			x"0000" when x"B486",
			x"0000" when x"B487",
			x"0000" when x"B488",
			x"0000" when x"B489",
			x"0000" when x"B48A",
			x"0000" when x"B48B",
			x"0000" when x"B48C",
			x"0000" when x"B48D",
			x"0000" when x"B48E",
			x"0000" when x"B48F",
			x"0000" when x"B490",
			x"0000" when x"B491",
			x"0000" when x"B492",
			x"0000" when x"B493",
			x"0000" when x"B494",
			x"0000" when x"B495",
			x"0000" when x"B496",
			x"0000" when x"B497",
			x"0000" when x"B498",
			x"0000" when x"B499",
			x"0000" when x"B49A",
			x"0000" when x"B49B",
			x"0000" when x"B49C",
			x"0000" when x"B49D",
			x"0000" when x"B49E",
			x"0000" when x"B49F",
			x"0000" when x"B4A0",
			x"0000" when x"B4A1",
			x"0000" when x"B4A2",
			x"0000" when x"B4A3",
			x"0000" when x"B4A4",
			x"0000" when x"B4A5",
			x"0000" when x"B4A6",
			x"0000" when x"B4A7",
			x"0000" when x"B4A8",
			x"0000" when x"B4A9",
			x"0000" when x"B4AA",
			x"0000" when x"B4AB",
			x"0000" when x"B4AC",
			x"0000" when x"B4AD",
			x"0000" when x"B4AE",
			x"0000" when x"B4AF",
			x"0000" when x"B4B0",
			x"0000" when x"B4B1",
			x"0000" when x"B4B2",
			x"0000" when x"B4B3",
			x"0000" when x"B4B4",
			x"0000" when x"B4B5",
			x"0000" when x"B4B6",
			x"0000" when x"B4B7",
			x"0000" when x"B4B8",
			x"0000" when x"B4B9",
			x"0000" when x"B4BA",
			x"0000" when x"B4BB",
			x"0000" when x"B4BC",
			x"0000" when x"B4BD",
			x"0000" when x"B4BE",
			x"0000" when x"B4BF",
			x"0000" when x"B4C0",
			x"0000" when x"B4C1",
			x"0000" when x"B4C2",
			x"0000" when x"B4C3",
			x"0000" when x"B4C4",
			x"0000" when x"B4C5",
			x"0000" when x"B4C6",
			x"0000" when x"B4C7",
			x"0000" when x"B4C8",
			x"0000" when x"B4C9",
			x"0000" when x"B4CA",
			x"0000" when x"B4CB",
			x"0000" when x"B4CC",
			x"0000" when x"B4CD",
			x"0000" when x"B4CE",
			x"0000" when x"B4CF",
			x"0000" when x"B4D0",
			x"0000" when x"B4D1",
			x"0000" when x"B4D2",
			x"0000" when x"B4D3",
			x"0000" when x"B4D4",
			x"0000" when x"B4D5",
			x"0000" when x"B4D6",
			x"0000" when x"B4D7",
			x"0000" when x"B4D8",
			x"0000" when x"B4D9",
			x"0000" when x"B4DA",
			x"0000" when x"B4DB",
			x"0000" when x"B4DC",
			x"0000" when x"B4DD",
			x"0000" when x"B4DE",
			x"0000" when x"B4DF",
			x"0000" when x"B4E0",
			x"0000" when x"B4E1",
			x"0000" when x"B4E2",
			x"0000" when x"B4E3",
			x"0000" when x"B4E4",
			x"0000" when x"B4E5",
			x"0000" when x"B4E6",
			x"0000" when x"B4E7",
			x"0000" when x"B4E8",
			x"0000" when x"B4E9",
			x"0000" when x"B4EA",
			x"0000" when x"B4EB",
			x"0000" when x"B4EC",
			x"0000" when x"B4ED",
			x"0000" when x"B4EE",
			x"0000" when x"B4EF",
			x"0000" when x"B4F0",
			x"0000" when x"B4F1",
			x"0000" when x"B4F2",
			x"0000" when x"B4F3",
			x"0000" when x"B4F4",
			x"0000" when x"B4F5",
			x"0000" when x"B4F6",
			x"0000" when x"B4F7",
			x"0000" when x"B4F8",
			x"0000" when x"B4F9",
			x"0000" when x"B4FA",
			x"0000" when x"B4FB",
			x"0000" when x"B4FC",
			x"0000" when x"B4FD",
			x"0000" when x"B4FE",
			x"0000" when x"B4FF",
			x"0000" when x"B500",
			x"0000" when x"B501",
			x"0000" when x"B502",
			x"0000" when x"B503",
			x"0000" when x"B504",
			x"0000" when x"B505",
			x"0000" when x"B506",
			x"0000" when x"B507",
			x"0000" when x"B508",
			x"0000" when x"B509",
			x"0000" when x"B50A",
			x"0000" when x"B50B",
			x"0000" when x"B50C",
			x"0000" when x"B50D",
			x"0000" when x"B50E",
			x"0000" when x"B50F",
			x"0000" when x"B510",
			x"0000" when x"B511",
			x"0000" when x"B512",
			x"0000" when x"B513",
			x"0000" when x"B514",
			x"0000" when x"B515",
			x"0000" when x"B516",
			x"0000" when x"B517",
			x"0000" when x"B518",
			x"0000" when x"B519",
			x"0000" when x"B51A",
			x"0000" when x"B51B",
			x"0000" when x"B51C",
			x"0000" when x"B51D",
			x"0000" when x"B51E",
			x"0000" when x"B51F",
			x"0000" when x"B520",
			x"0000" when x"B521",
			x"0000" when x"B522",
			x"0000" when x"B523",
			x"0000" when x"B524",
			x"0000" when x"B525",
			x"0000" when x"B526",
			x"0000" when x"B527",
			x"0000" when x"B528",
			x"0000" when x"B529",
			x"0000" when x"B52A",
			x"0000" when x"B52B",
			x"0000" when x"B52C",
			x"0000" when x"B52D",
			x"0000" when x"B52E",
			x"0000" when x"B52F",
			x"0000" when x"B530",
			x"0000" when x"B531",
			x"0000" when x"B532",
			x"0000" when x"B533",
			x"0000" when x"B534",
			x"0000" when x"B535",
			x"0000" when x"B536",
			x"0000" when x"B537",
			x"0000" when x"B538",
			x"0000" when x"B539",
			x"0000" when x"B53A",
			x"0000" when x"B53B",
			x"0000" when x"B53C",
			x"0000" when x"B53D",
			x"0000" when x"B53E",
			x"0000" when x"B53F",
			x"0000" when x"B540",
			x"0000" when x"B541",
			x"0000" when x"B542",
			x"0000" when x"B543",
			x"0000" when x"B544",
			x"0000" when x"B545",
			x"0000" when x"B546",
			x"0000" when x"B547",
			x"0000" when x"B548",
			x"0000" when x"B549",
			x"0000" when x"B54A",
			x"0000" when x"B54B",
			x"0000" when x"B54C",
			x"0000" when x"B54D",
			x"0000" when x"B54E",
			x"0000" when x"B54F",
			x"0000" when x"B550",
			x"0000" when x"B551",
			x"0000" when x"B552",
			x"0000" when x"B553",
			x"0000" when x"B554",
			x"0000" when x"B555",
			x"0000" when x"B556",
			x"0000" when x"B557",
			x"0000" when x"B558",
			x"0000" when x"B559",
			x"0000" when x"B55A",
			x"0000" when x"B55B",
			x"0000" when x"B55C",
			x"0000" when x"B55D",
			x"0000" when x"B55E",
			x"0000" when x"B55F",
			x"0000" when x"B560",
			x"0000" when x"B561",
			x"0000" when x"B562",
			x"0000" when x"B563",
			x"0000" when x"B564",
			x"0000" when x"B565",
			x"0000" when x"B566",
			x"0000" when x"B567",
			x"0000" when x"B568",
			x"0000" when x"B569",
			x"0000" when x"B56A",
			x"0000" when x"B56B",
			x"0000" when x"B56C",
			x"0000" when x"B56D",
			x"0000" when x"B56E",
			x"0000" when x"B56F",
			x"0000" when x"B570",
			x"0000" when x"B571",
			x"0000" when x"B572",
			x"0000" when x"B573",
			x"0000" when x"B574",
			x"0000" when x"B575",
			x"0000" when x"B576",
			x"0000" when x"B577",
			x"0000" when x"B578",
			x"0000" when x"B579",
			x"0000" when x"B57A",
			x"0000" when x"B57B",
			x"0000" when x"B57C",
			x"0000" when x"B57D",
			x"0000" when x"B57E",
			x"0000" when x"B57F",
			x"0000" when x"B580",
			x"0000" when x"B581",
			x"0000" when x"B582",
			x"0000" when x"B583",
			x"0000" when x"B584",
			x"0000" when x"B585",
			x"0000" when x"B586",
			x"0000" when x"B587",
			x"0000" when x"B588",
			x"0000" when x"B589",
			x"0000" when x"B58A",
			x"0000" when x"B58B",
			x"0000" when x"B58C",
			x"0000" when x"B58D",
			x"0000" when x"B58E",
			x"0000" when x"B58F",
			x"0000" when x"B590",
			x"0000" when x"B591",
			x"0000" when x"B592",
			x"0000" when x"B593",
			x"0000" when x"B594",
			x"0000" when x"B595",
			x"0000" when x"B596",
			x"0000" when x"B597",
			x"0000" when x"B598",
			x"0000" when x"B599",
			x"0000" when x"B59A",
			x"0000" when x"B59B",
			x"0000" when x"B59C",
			x"0000" when x"B59D",
			x"0000" when x"B59E",
			x"0000" when x"B59F",
			x"0000" when x"B5A0",
			x"0000" when x"B5A1",
			x"0000" when x"B5A2",
			x"0000" when x"B5A3",
			x"0000" when x"B5A4",
			x"0000" when x"B5A5",
			x"0000" when x"B5A6",
			x"0000" when x"B5A7",
			x"0000" when x"B5A8",
			x"0000" when x"B5A9",
			x"0000" when x"B5AA",
			x"0000" when x"B5AB",
			x"0000" when x"B5AC",
			x"0000" when x"B5AD",
			x"0000" when x"B5AE",
			x"0000" when x"B5AF",
			x"0000" when x"B5B0",
			x"0000" when x"B5B1",
			x"0000" when x"B5B2",
			x"0000" when x"B5B3",
			x"0000" when x"B5B4",
			x"0000" when x"B5B5",
			x"0000" when x"B5B6",
			x"0000" when x"B5B7",
			x"0000" when x"B5B8",
			x"0000" when x"B5B9",
			x"0000" when x"B5BA",
			x"0000" when x"B5BB",
			x"0000" when x"B5BC",
			x"0000" when x"B5BD",
			x"0000" when x"B5BE",
			x"0000" when x"B5BF",
			x"0000" when x"B5C0",
			x"0000" when x"B5C1",
			x"0000" when x"B5C2",
			x"0000" when x"B5C3",
			x"0000" when x"B5C4",
			x"0000" when x"B5C5",
			x"0000" when x"B5C6",
			x"0000" when x"B5C7",
			x"0000" when x"B5C8",
			x"0000" when x"B5C9",
			x"0000" when x"B5CA",
			x"0000" when x"B5CB",
			x"0000" when x"B5CC",
			x"0000" when x"B5CD",
			x"0000" when x"B5CE",
			x"0000" when x"B5CF",
			x"0000" when x"B5D0",
			x"0000" when x"B5D1",
			x"0000" when x"B5D2",
			x"0000" when x"B5D3",
			x"0000" when x"B5D4",
			x"0000" when x"B5D5",
			x"0000" when x"B5D6",
			x"0000" when x"B5D7",
			x"0000" when x"B5D8",
			x"0000" when x"B5D9",
			x"0000" when x"B5DA",
			x"0000" when x"B5DB",
			x"0000" when x"B5DC",
			x"0000" when x"B5DD",
			x"0000" when x"B5DE",
			x"0000" when x"B5DF",
			x"0000" when x"B5E0",
			x"0000" when x"B5E1",
			x"0000" when x"B5E2",
			x"0000" when x"B5E3",
			x"0000" when x"B5E4",
			x"0000" when x"B5E5",
			x"0000" when x"B5E6",
			x"0000" when x"B5E7",
			x"0000" when x"B5E8",
			x"0000" when x"B5E9",
			x"0000" when x"B5EA",
			x"0000" when x"B5EB",
			x"0000" when x"B5EC",
			x"0000" when x"B5ED",
			x"0000" when x"B5EE",
			x"0000" when x"B5EF",
			x"0000" when x"B5F0",
			x"0000" when x"B5F1",
			x"0000" when x"B5F2",
			x"0000" when x"B5F3",
			x"0000" when x"B5F4",
			x"0000" when x"B5F5",
			x"0000" when x"B5F6",
			x"0000" when x"B5F7",
			x"0000" when x"B5F8",
			x"0000" when x"B5F9",
			x"0000" when x"B5FA",
			x"0000" when x"B5FB",
			x"0000" when x"B5FC",
			x"0000" when x"B5FD",
			x"0000" when x"B5FE",
			x"0000" when x"B5FF",
			x"0000" when x"B600",
			x"0000" when x"B601",
			x"0000" when x"B602",
			x"0000" when x"B603",
			x"0000" when x"B604",
			x"0000" when x"B605",
			x"0000" when x"B606",
			x"0000" when x"B607",
			x"0000" when x"B608",
			x"0000" when x"B609",
			x"0000" when x"B60A",
			x"0000" when x"B60B",
			x"0000" when x"B60C",
			x"0000" when x"B60D",
			x"0000" when x"B60E",
			x"0000" when x"B60F",
			x"0000" when x"B610",
			x"0000" when x"B611",
			x"0000" when x"B612",
			x"0000" when x"B613",
			x"0000" when x"B614",
			x"0000" when x"B615",
			x"0000" when x"B616",
			x"0000" when x"B617",
			x"0000" when x"B618",
			x"0000" when x"B619",
			x"0000" when x"B61A",
			x"0000" when x"B61B",
			x"0000" when x"B61C",
			x"0000" when x"B61D",
			x"0000" when x"B61E",
			x"0000" when x"B61F",
			x"0000" when x"B620",
			x"0000" when x"B621",
			x"0000" when x"B622",
			x"0000" when x"B623",
			x"0000" when x"B624",
			x"0000" when x"B625",
			x"0000" when x"B626",
			x"0000" when x"B627",
			x"0000" when x"B628",
			x"0000" when x"B629",
			x"0000" when x"B62A",
			x"0000" when x"B62B",
			x"0000" when x"B62C",
			x"0000" when x"B62D",
			x"0000" when x"B62E",
			x"0000" when x"B62F",
			x"0000" when x"B630",
			x"0000" when x"B631",
			x"0000" when x"B632",
			x"0000" when x"B633",
			x"0000" when x"B634",
			x"0000" when x"B635",
			x"0000" when x"B636",
			x"0000" when x"B637",
			x"0000" when x"B638",
			x"0000" when x"B639",
			x"0000" when x"B63A",
			x"0000" when x"B63B",
			x"0000" when x"B63C",
			x"0000" when x"B63D",
			x"0000" when x"B63E",
			x"0000" when x"B63F",
			x"0000" when x"B640",
			x"0000" when x"B641",
			x"0000" when x"B642",
			x"0000" when x"B643",
			x"0000" when x"B644",
			x"0000" when x"B645",
			x"0000" when x"B646",
			x"0000" when x"B647",
			x"0000" when x"B648",
			x"0000" when x"B649",
			x"0000" when x"B64A",
			x"0000" when x"B64B",
			x"0000" when x"B64C",
			x"0000" when x"B64D",
			x"0000" when x"B64E",
			x"0000" when x"B64F",
			x"0000" when x"B650",
			x"0000" when x"B651",
			x"0000" when x"B652",
			x"0000" when x"B653",
			x"0000" when x"B654",
			x"0000" when x"B655",
			x"0000" when x"B656",
			x"0000" when x"B657",
			x"0000" when x"B658",
			x"0000" when x"B659",
			x"0000" when x"B65A",
			x"0000" when x"B65B",
			x"0000" when x"B65C",
			x"0000" when x"B65D",
			x"0000" when x"B65E",
			x"0000" when x"B65F",
			x"0000" when x"B660",
			x"0000" when x"B661",
			x"0000" when x"B662",
			x"0000" when x"B663",
			x"0000" when x"B664",
			x"0000" when x"B665",
			x"0000" when x"B666",
			x"0000" when x"B667",
			x"0000" when x"B668",
			x"0000" when x"B669",
			x"0000" when x"B66A",
			x"0000" when x"B66B",
			x"0000" when x"B66C",
			x"0000" when x"B66D",
			x"0000" when x"B66E",
			x"0000" when x"B66F",
			x"0000" when x"B670",
			x"0000" when x"B671",
			x"0000" when x"B672",
			x"0000" when x"B673",
			x"0000" when x"B674",
			x"0000" when x"B675",
			x"0000" when x"B676",
			x"0000" when x"B677",
			x"0000" when x"B678",
			x"0000" when x"B679",
			x"0000" when x"B67A",
			x"0000" when x"B67B",
			x"0000" when x"B67C",
			x"0000" when x"B67D",
			x"0000" when x"B67E",
			x"0000" when x"B67F",
			x"0000" when x"B680",
			x"0000" when x"B681",
			x"0000" when x"B682",
			x"0000" when x"B683",
			x"0000" when x"B684",
			x"0000" when x"B685",
			x"0000" when x"B686",
			x"0000" when x"B687",
			x"0000" when x"B688",
			x"0000" when x"B689",
			x"0000" when x"B68A",
			x"0000" when x"B68B",
			x"0000" when x"B68C",
			x"0000" when x"B68D",
			x"0000" when x"B68E",
			x"0000" when x"B68F",
			x"0000" when x"B690",
			x"0000" when x"B691",
			x"0000" when x"B692",
			x"0000" when x"B693",
			x"0000" when x"B694",
			x"0000" when x"B695",
			x"0000" when x"B696",
			x"0000" when x"B697",
			x"0000" when x"B698",
			x"0000" when x"B699",
			x"0000" when x"B69A",
			x"0000" when x"B69B",
			x"0000" when x"B69C",
			x"0000" when x"B69D",
			x"0000" when x"B69E",
			x"0000" when x"B69F",
			x"0000" when x"B6A0",
			x"0000" when x"B6A1",
			x"0000" when x"B6A2",
			x"0000" when x"B6A3",
			x"0000" when x"B6A4",
			x"0000" when x"B6A5",
			x"0000" when x"B6A6",
			x"0000" when x"B6A7",
			x"0000" when x"B6A8",
			x"0000" when x"B6A9",
			x"0000" when x"B6AA",
			x"0000" when x"B6AB",
			x"0000" when x"B6AC",
			x"0000" when x"B6AD",
			x"0000" when x"B6AE",
			x"0000" when x"B6AF",
			x"0000" when x"B6B0",
			x"0000" when x"B6B1",
			x"0000" when x"B6B2",
			x"0000" when x"B6B3",
			x"0000" when x"B6B4",
			x"0000" when x"B6B5",
			x"0000" when x"B6B6",
			x"0000" when x"B6B7",
			x"0000" when x"B6B8",
			x"0000" when x"B6B9",
			x"0000" when x"B6BA",
			x"0000" when x"B6BB",
			x"0000" when x"B6BC",
			x"0000" when x"B6BD",
			x"0000" when x"B6BE",
			x"0000" when x"B6BF",
			x"0000" when x"B6C0",
			x"0000" when x"B6C1",
			x"0000" when x"B6C2",
			x"0000" when x"B6C3",
			x"0000" when x"B6C4",
			x"0000" when x"B6C5",
			x"0000" when x"B6C6",
			x"0000" when x"B6C7",
			x"0000" when x"B6C8",
			x"0000" when x"B6C9",
			x"0000" when x"B6CA",
			x"0000" when x"B6CB",
			x"0000" when x"B6CC",
			x"0000" when x"B6CD",
			x"0000" when x"B6CE",
			x"0000" when x"B6CF",
			x"0000" when x"B6D0",
			x"0000" when x"B6D1",
			x"0000" when x"B6D2",
			x"0000" when x"B6D3",
			x"0000" when x"B6D4",
			x"0000" when x"B6D5",
			x"0000" when x"B6D6",
			x"0000" when x"B6D7",
			x"0000" when x"B6D8",
			x"0000" when x"B6D9",
			x"0000" when x"B6DA",
			x"0000" when x"B6DB",
			x"0000" when x"B6DC",
			x"0000" when x"B6DD",
			x"0000" when x"B6DE",
			x"0000" when x"B6DF",
			x"0000" when x"B6E0",
			x"0000" when x"B6E1",
			x"0000" when x"B6E2",
			x"0000" when x"B6E3",
			x"0000" when x"B6E4",
			x"0000" when x"B6E5",
			x"0000" when x"B6E6",
			x"0000" when x"B6E7",
			x"0000" when x"B6E8",
			x"0000" when x"B6E9",
			x"0000" when x"B6EA",
			x"0000" when x"B6EB",
			x"0000" when x"B6EC",
			x"0000" when x"B6ED",
			x"0000" when x"B6EE",
			x"0000" when x"B6EF",
			x"0000" when x"B6F0",
			x"0000" when x"B6F1",
			x"0000" when x"B6F2",
			x"0000" when x"B6F3",
			x"0000" when x"B6F4",
			x"0000" when x"B6F5",
			x"0000" when x"B6F6",
			x"0000" when x"B6F7",
			x"0000" when x"B6F8",
			x"0000" when x"B6F9",
			x"0000" when x"B6FA",
			x"0000" when x"B6FB",
			x"0000" when x"B6FC",
			x"0000" when x"B6FD",
			x"0000" when x"B6FE",
			x"0000" when x"B6FF",
			x"0000" when x"B700",
			x"0000" when x"B701",
			x"0000" when x"B702",
			x"0000" when x"B703",
			x"0000" when x"B704",
			x"0000" when x"B705",
			x"0000" when x"B706",
			x"0000" when x"B707",
			x"0000" when x"B708",
			x"0000" when x"B709",
			x"0000" when x"B70A",
			x"0000" when x"B70B",
			x"0000" when x"B70C",
			x"0000" when x"B70D",
			x"0000" when x"B70E",
			x"0000" when x"B70F",
			x"0000" when x"B710",
			x"0000" when x"B711",
			x"0000" when x"B712",
			x"0000" when x"B713",
			x"0000" when x"B714",
			x"0000" when x"B715",
			x"0000" when x"B716",
			x"0000" when x"B717",
			x"0000" when x"B718",
			x"0000" when x"B719",
			x"0000" when x"B71A",
			x"0000" when x"B71B",
			x"0000" when x"B71C",
			x"0000" when x"B71D",
			x"0000" when x"B71E",
			x"0000" when x"B71F",
			x"0000" when x"B720",
			x"0000" when x"B721",
			x"0000" when x"B722",
			x"0000" when x"B723",
			x"0000" when x"B724",
			x"0000" when x"B725",
			x"0000" when x"B726",
			x"0000" when x"B727",
			x"0000" when x"B728",
			x"0000" when x"B729",
			x"0000" when x"B72A",
			x"0000" when x"B72B",
			x"0000" when x"B72C",
			x"0000" when x"B72D",
			x"0000" when x"B72E",
			x"0000" when x"B72F",
			x"0000" when x"B730",
			x"0000" when x"B731",
			x"0000" when x"B732",
			x"0000" when x"B733",
			x"0000" when x"B734",
			x"0000" when x"B735",
			x"0000" when x"B736",
			x"0000" when x"B737",
			x"0000" when x"B738",
			x"0000" when x"B739",
			x"0000" when x"B73A",
			x"0000" when x"B73B",
			x"0000" when x"B73C",
			x"0000" when x"B73D",
			x"0000" when x"B73E",
			x"0000" when x"B73F",
			x"0000" when x"B740",
			x"0000" when x"B741",
			x"0000" when x"B742",
			x"0000" when x"B743",
			x"0000" when x"B744",
			x"0000" when x"B745",
			x"0000" when x"B746",
			x"0000" when x"B747",
			x"0000" when x"B748",
			x"0000" when x"B749",
			x"0000" when x"B74A",
			x"0000" when x"B74B",
			x"0000" when x"B74C",
			x"0000" when x"B74D",
			x"0000" when x"B74E",
			x"0000" when x"B74F",
			x"0000" when x"B750",
			x"0000" when x"B751",
			x"0000" when x"B752",
			x"0000" when x"B753",
			x"0000" when x"B754",
			x"0000" when x"B755",
			x"0000" when x"B756",
			x"0000" when x"B757",
			x"0000" when x"B758",
			x"0000" when x"B759",
			x"0000" when x"B75A",
			x"0000" when x"B75B",
			x"0000" when x"B75C",
			x"0000" when x"B75D",
			x"0000" when x"B75E",
			x"0000" when x"B75F",
			x"0000" when x"B760",
			x"0000" when x"B761",
			x"0000" when x"B762",
			x"0000" when x"B763",
			x"0000" when x"B764",
			x"0000" when x"B765",
			x"0000" when x"B766",
			x"0000" when x"B767",
			x"0000" when x"B768",
			x"0000" when x"B769",
			x"0000" when x"B76A",
			x"0000" when x"B76B",
			x"0000" when x"B76C",
			x"0000" when x"B76D",
			x"0000" when x"B76E",
			x"0000" when x"B76F",
			x"0000" when x"B770",
			x"0000" when x"B771",
			x"0000" when x"B772",
			x"0000" when x"B773",
			x"0000" when x"B774",
			x"0000" when x"B775",
			x"0000" when x"B776",
			x"0000" when x"B777",
			x"0000" when x"B778",
			x"0000" when x"B779",
			x"0000" when x"B77A",
			x"0000" when x"B77B",
			x"0000" when x"B77C",
			x"0000" when x"B77D",
			x"0000" when x"B77E",
			x"0000" when x"B77F",
			x"0000" when x"B780",
			x"0000" when x"B781",
			x"0000" when x"B782",
			x"0000" when x"B783",
			x"0000" when x"B784",
			x"0000" when x"B785",
			x"0000" when x"B786",
			x"0000" when x"B787",
			x"0000" when x"B788",
			x"0000" when x"B789",
			x"0000" when x"B78A",
			x"0000" when x"B78B",
			x"0000" when x"B78C",
			x"0000" when x"B78D",
			x"0000" when x"B78E",
			x"0000" when x"B78F",
			x"0000" when x"B790",
			x"0000" when x"B791",
			x"0000" when x"B792",
			x"0000" when x"B793",
			x"0000" when x"B794",
			x"0000" when x"B795",
			x"0000" when x"B796",
			x"0000" when x"B797",
			x"0000" when x"B798",
			x"0000" when x"B799",
			x"0000" when x"B79A",
			x"0000" when x"B79B",
			x"0000" when x"B79C",
			x"0000" when x"B79D",
			x"0000" when x"B79E",
			x"0000" when x"B79F",
			x"0000" when x"B7A0",
			x"0000" when x"B7A1",
			x"0000" when x"B7A2",
			x"0000" when x"B7A3",
			x"0000" when x"B7A4",
			x"0000" when x"B7A5",
			x"0000" when x"B7A6",
			x"0000" when x"B7A7",
			x"0000" when x"B7A8",
			x"0000" when x"B7A9",
			x"0000" when x"B7AA",
			x"0000" when x"B7AB",
			x"0000" when x"B7AC",
			x"0000" when x"B7AD",
			x"0000" when x"B7AE",
			x"0000" when x"B7AF",
			x"0000" when x"B7B0",
			x"0000" when x"B7B1",
			x"0000" when x"B7B2",
			x"0000" when x"B7B3",
			x"0000" when x"B7B4",
			x"0000" when x"B7B5",
			x"0000" when x"B7B6",
			x"0000" when x"B7B7",
			x"0000" when x"B7B8",
			x"0000" when x"B7B9",
			x"0000" when x"B7BA",
			x"0000" when x"B7BB",
			x"0000" when x"B7BC",
			x"0000" when x"B7BD",
			x"0000" when x"B7BE",
			x"0000" when x"B7BF",
			x"0000" when x"B7C0",
			x"0000" when x"B7C1",
			x"0000" when x"B7C2",
			x"0000" when x"B7C3",
			x"0000" when x"B7C4",
			x"0000" when x"B7C5",
			x"0000" when x"B7C6",
			x"0000" when x"B7C7",
			x"0000" when x"B7C8",
			x"0000" when x"B7C9",
			x"0000" when x"B7CA",
			x"0000" when x"B7CB",
			x"0000" when x"B7CC",
			x"0000" when x"B7CD",
			x"0000" when x"B7CE",
			x"0000" when x"B7CF",
			x"0000" when x"B7D0",
			x"0000" when x"B7D1",
			x"0000" when x"B7D2",
			x"0000" when x"B7D3",
			x"0000" when x"B7D4",
			x"0000" when x"B7D5",
			x"0000" when x"B7D6",
			x"0000" when x"B7D7",
			x"0000" when x"B7D8",
			x"0000" when x"B7D9",
			x"0000" when x"B7DA",
			x"0000" when x"B7DB",
			x"0000" when x"B7DC",
			x"0000" when x"B7DD",
			x"0000" when x"B7DE",
			x"0000" when x"B7DF",
			x"0000" when x"B7E0",
			x"0000" when x"B7E1",
			x"0000" when x"B7E2",
			x"0000" when x"B7E3",
			x"0000" when x"B7E4",
			x"0000" when x"B7E5",
			x"0000" when x"B7E6",
			x"0000" when x"B7E7",
			x"0000" when x"B7E8",
			x"0000" when x"B7E9",
			x"0000" when x"B7EA",
			x"0000" when x"B7EB",
			x"0000" when x"B7EC",
			x"0000" when x"B7ED",
			x"0000" when x"B7EE",
			x"0000" when x"B7EF",
			x"0000" when x"B7F0",
			x"0000" when x"B7F1",
			x"0000" when x"B7F2",
			x"0000" when x"B7F3",
			x"0000" when x"B7F4",
			x"0000" when x"B7F5",
			x"0000" when x"B7F6",
			x"0000" when x"B7F7",
			x"0000" when x"B7F8",
			x"0000" when x"B7F9",
			x"0000" when x"B7FA",
			x"0000" when x"B7FB",
			x"0000" when x"B7FC",
			x"0000" when x"B7FD",
			x"0000" when x"B7FE",
			x"0000" when x"B7FF",
			x"0000" when x"B800",
			x"0000" when x"B801",
			x"0000" when x"B802",
			x"0000" when x"B803",
			x"0000" when x"B804",
			x"0000" when x"B805",
			x"0000" when x"B806",
			x"0000" when x"B807",
			x"0000" when x"B808",
			x"0000" when x"B809",
			x"0000" when x"B80A",
			x"0000" when x"B80B",
			x"0000" when x"B80C",
			x"0000" when x"B80D",
			x"0000" when x"B80E",
			x"0000" when x"B80F",
			x"0000" when x"B810",
			x"0000" when x"B811",
			x"0000" when x"B812",
			x"0000" when x"B813",
			x"0000" when x"B814",
			x"0000" when x"B815",
			x"0000" when x"B816",
			x"0000" when x"B817",
			x"0000" when x"B818",
			x"0000" when x"B819",
			x"0000" when x"B81A",
			x"0000" when x"B81B",
			x"0000" when x"B81C",
			x"0000" when x"B81D",
			x"0000" when x"B81E",
			x"0000" when x"B81F",
			x"0000" when x"B820",
			x"0000" when x"B821",
			x"0000" when x"B822",
			x"0000" when x"B823",
			x"0000" when x"B824",
			x"0000" when x"B825",
			x"0000" when x"B826",
			x"0000" when x"B827",
			x"0000" when x"B828",
			x"0000" when x"B829",
			x"0000" when x"B82A",
			x"0000" when x"B82B",
			x"0000" when x"B82C",
			x"0000" when x"B82D",
			x"0000" when x"B82E",
			x"0000" when x"B82F",
			x"0000" when x"B830",
			x"0000" when x"B831",
			x"0000" when x"B832",
			x"0000" when x"B833",
			x"0000" when x"B834",
			x"0000" when x"B835",
			x"0000" when x"B836",
			x"0000" when x"B837",
			x"0000" when x"B838",
			x"0000" when x"B839",
			x"0000" when x"B83A",
			x"0000" when x"B83B",
			x"0000" when x"B83C",
			x"0000" when x"B83D",
			x"0000" when x"B83E",
			x"0000" when x"B83F",
			x"0000" when x"B840",
			x"0000" when x"B841",
			x"0000" when x"B842",
			x"0000" when x"B843",
			x"0000" when x"B844",
			x"0000" when x"B845",
			x"0000" when x"B846",
			x"0000" when x"B847",
			x"0000" when x"B848",
			x"0000" when x"B849",
			x"0000" when x"B84A",
			x"0000" when x"B84B",
			x"0000" when x"B84C",
			x"0000" when x"B84D",
			x"0000" when x"B84E",
			x"0000" when x"B84F",
			x"0000" when x"B850",
			x"0000" when x"B851",
			x"0000" when x"B852",
			x"0000" when x"B853",
			x"0000" when x"B854",
			x"0000" when x"B855",
			x"0000" when x"B856",
			x"0000" when x"B857",
			x"0000" when x"B858",
			x"0000" when x"B859",
			x"0000" when x"B85A",
			x"0000" when x"B85B",
			x"0000" when x"B85C",
			x"0000" when x"B85D",
			x"0000" when x"B85E",
			x"0000" when x"B85F",
			x"0000" when x"B860",
			x"0000" when x"B861",
			x"0000" when x"B862",
			x"0000" when x"B863",
			x"0000" when x"B864",
			x"0000" when x"B865",
			x"0000" when x"B866",
			x"0000" when x"B867",
			x"0000" when x"B868",
			x"0000" when x"B869",
			x"0000" when x"B86A",
			x"0000" when x"B86B",
			x"0000" when x"B86C",
			x"0000" when x"B86D",
			x"0000" when x"B86E",
			x"0000" when x"B86F",
			x"0000" when x"B870",
			x"0000" when x"B871",
			x"0000" when x"B872",
			x"0000" when x"B873",
			x"0000" when x"B874",
			x"0000" when x"B875",
			x"0000" when x"B876",
			x"0000" when x"B877",
			x"0000" when x"B878",
			x"0000" when x"B879",
			x"0000" when x"B87A",
			x"0000" when x"B87B",
			x"0000" when x"B87C",
			x"0000" when x"B87D",
			x"0000" when x"B87E",
			x"0000" when x"B87F",
			x"0000" when x"B880",
			x"0000" when x"B881",
			x"0000" when x"B882",
			x"0000" when x"B883",
			x"0000" when x"B884",
			x"0000" when x"B885",
			x"0000" when x"B886",
			x"0000" when x"B887",
			x"0000" when x"B888",
			x"0000" when x"B889",
			x"0000" when x"B88A",
			x"0000" when x"B88B",
			x"0000" when x"B88C",
			x"0000" when x"B88D",
			x"0000" when x"B88E",
			x"0000" when x"B88F",
			x"0000" when x"B890",
			x"0000" when x"B891",
			x"0000" when x"B892",
			x"0000" when x"B893",
			x"0000" when x"B894",
			x"0000" when x"B895",
			x"0000" when x"B896",
			x"0000" when x"B897",
			x"0000" when x"B898",
			x"0000" when x"B899",
			x"0000" when x"B89A",
			x"0000" when x"B89B",
			x"0000" when x"B89C",
			x"0000" when x"B89D",
			x"0000" when x"B89E",
			x"0000" when x"B89F",
			x"0000" when x"B8A0",
			x"0000" when x"B8A1",
			x"0000" when x"B8A2",
			x"0000" when x"B8A3",
			x"0000" when x"B8A4",
			x"0000" when x"B8A5",
			x"0000" when x"B8A6",
			x"0000" when x"B8A7",
			x"0000" when x"B8A8",
			x"0000" when x"B8A9",
			x"0000" when x"B8AA",
			x"0000" when x"B8AB",
			x"0000" when x"B8AC",
			x"0000" when x"B8AD",
			x"0000" when x"B8AE",
			x"0000" when x"B8AF",
			x"0000" when x"B8B0",
			x"0000" when x"B8B1",
			x"0000" when x"B8B2",
			x"0000" when x"B8B3",
			x"0000" when x"B8B4",
			x"0000" when x"B8B5",
			x"0000" when x"B8B6",
			x"0000" when x"B8B7",
			x"0000" when x"B8B8",
			x"0000" when x"B8B9",
			x"0000" when x"B8BA",
			x"0000" when x"B8BB",
			x"0000" when x"B8BC",
			x"0000" when x"B8BD",
			x"0000" when x"B8BE",
			x"0000" when x"B8BF",
			x"0000" when x"B8C0",
			x"0000" when x"B8C1",
			x"0000" when x"B8C2",
			x"0000" when x"B8C3",
			x"0000" when x"B8C4",
			x"0000" when x"B8C5",
			x"0000" when x"B8C6",
			x"0000" when x"B8C7",
			x"0000" when x"B8C8",
			x"0000" when x"B8C9",
			x"0000" when x"B8CA",
			x"0000" when x"B8CB",
			x"0000" when x"B8CC",
			x"0000" when x"B8CD",
			x"0000" when x"B8CE",
			x"0000" when x"B8CF",
			x"0000" when x"B8D0",
			x"0000" when x"B8D1",
			x"0000" when x"B8D2",
			x"0000" when x"B8D3",
			x"0000" when x"B8D4",
			x"0000" when x"B8D5",
			x"0000" when x"B8D6",
			x"0000" when x"B8D7",
			x"0000" when x"B8D8",
			x"0000" when x"B8D9",
			x"0000" when x"B8DA",
			x"0000" when x"B8DB",
			x"0000" when x"B8DC",
			x"0000" when x"B8DD",
			x"0000" when x"B8DE",
			x"0000" when x"B8DF",
			x"0000" when x"B8E0",
			x"0000" when x"B8E1",
			x"0000" when x"B8E2",
			x"0000" when x"B8E3",
			x"0000" when x"B8E4",
			x"0000" when x"B8E5",
			x"0000" when x"B8E6",
			x"0000" when x"B8E7",
			x"0000" when x"B8E8",
			x"0000" when x"B8E9",
			x"0000" when x"B8EA",
			x"0000" when x"B8EB",
			x"0000" when x"B8EC",
			x"0000" when x"B8ED",
			x"0000" when x"B8EE",
			x"0000" when x"B8EF",
			x"0000" when x"B8F0",
			x"0000" when x"B8F1",
			x"0000" when x"B8F2",
			x"0000" when x"B8F3",
			x"0000" when x"B8F4",
			x"0000" when x"B8F5",
			x"0000" when x"B8F6",
			x"0000" when x"B8F7",
			x"0000" when x"B8F8",
			x"0000" when x"B8F9",
			x"0000" when x"B8FA",
			x"0000" when x"B8FB",
			x"0000" when x"B8FC",
			x"0000" when x"B8FD",
			x"0000" when x"B8FE",
			x"0000" when x"B8FF",
			x"0000" when x"B900",
			x"0000" when x"B901",
			x"0000" when x"B902",
			x"0000" when x"B903",
			x"0000" when x"B904",
			x"0000" when x"B905",
			x"0000" when x"B906",
			x"0000" when x"B907",
			x"0000" when x"B908",
			x"0000" when x"B909",
			x"0000" when x"B90A",
			x"0000" when x"B90B",
			x"0000" when x"B90C",
			x"0000" when x"B90D",
			x"0000" when x"B90E",
			x"0000" when x"B90F",
			x"0000" when x"B910",
			x"0000" when x"B911",
			x"0000" when x"B912",
			x"0000" when x"B913",
			x"0000" when x"B914",
			x"0000" when x"B915",
			x"0000" when x"B916",
			x"0000" when x"B917",
			x"0000" when x"B918",
			x"0000" when x"B919",
			x"0000" when x"B91A",
			x"0000" when x"B91B",
			x"0000" when x"B91C",
			x"0000" when x"B91D",
			x"0000" when x"B91E",
			x"0000" when x"B91F",
			x"0000" when x"B920",
			x"0000" when x"B921",
			x"0000" when x"B922",
			x"0000" when x"B923",
			x"0000" when x"B924",
			x"0000" when x"B925",
			x"0000" when x"B926",
			x"0000" when x"B927",
			x"0000" when x"B928",
			x"0000" when x"B929",
			x"0000" when x"B92A",
			x"0000" when x"B92B",
			x"0000" when x"B92C",
			x"0000" when x"B92D",
			x"0000" when x"B92E",
			x"0000" when x"B92F",
			x"0000" when x"B930",
			x"0000" when x"B931",
			x"0000" when x"B932",
			x"0000" when x"B933",
			x"0000" when x"B934",
			x"0000" when x"B935",
			x"0000" when x"B936",
			x"0000" when x"B937",
			x"0000" when x"B938",
			x"0000" when x"B939",
			x"0000" when x"B93A",
			x"0000" when x"B93B",
			x"0000" when x"B93C",
			x"0000" when x"B93D",
			x"0000" when x"B93E",
			x"0000" when x"B93F",
			x"0000" when x"B940",
			x"0000" when x"B941",
			x"0000" when x"B942",
			x"0000" when x"B943",
			x"0000" when x"B944",
			x"0000" when x"B945",
			x"0000" when x"B946",
			x"0000" when x"B947",
			x"0000" when x"B948",
			x"0000" when x"B949",
			x"0000" when x"B94A",
			x"0000" when x"B94B",
			x"0000" when x"B94C",
			x"0000" when x"B94D",
			x"0000" when x"B94E",
			x"0000" when x"B94F",
			x"0000" when x"B950",
			x"0000" when x"B951",
			x"0000" when x"B952",
			x"0000" when x"B953",
			x"0000" when x"B954",
			x"0000" when x"B955",
			x"0000" when x"B956",
			x"0000" when x"B957",
			x"0000" when x"B958",
			x"0000" when x"B959",
			x"0000" when x"B95A",
			x"0000" when x"B95B",
			x"0000" when x"B95C",
			x"0000" when x"B95D",
			x"0000" when x"B95E",
			x"0000" when x"B95F",
			x"0000" when x"B960",
			x"0000" when x"B961",
			x"0000" when x"B962",
			x"0000" when x"B963",
			x"0000" when x"B964",
			x"0000" when x"B965",
			x"0000" when x"B966",
			x"0000" when x"B967",
			x"0000" when x"B968",
			x"0000" when x"B969",
			x"0000" when x"B96A",
			x"0000" when x"B96B",
			x"0000" when x"B96C",
			x"0000" when x"B96D",
			x"0000" when x"B96E",
			x"0000" when x"B96F",
			x"0000" when x"B970",
			x"0000" when x"B971",
			x"0000" when x"B972",
			x"0000" when x"B973",
			x"0000" when x"B974",
			x"0000" when x"B975",
			x"0000" when x"B976",
			x"0000" when x"B977",
			x"0000" when x"B978",
			x"0000" when x"B979",
			x"0000" when x"B97A",
			x"0000" when x"B97B",
			x"0000" when x"B97C",
			x"0000" when x"B97D",
			x"0000" when x"B97E",
			x"0000" when x"B97F",
			x"0000" when x"B980",
			x"0000" when x"B981",
			x"0000" when x"B982",
			x"0000" when x"B983",
			x"0000" when x"B984",
			x"0000" when x"B985",
			x"0000" when x"B986",
			x"0000" when x"B987",
			x"0000" when x"B988",
			x"0000" when x"B989",
			x"0000" when x"B98A",
			x"0000" when x"B98B",
			x"0000" when x"B98C",
			x"0000" when x"B98D",
			x"0000" when x"B98E",
			x"0000" when x"B98F",
			x"0000" when x"B990",
			x"0000" when x"B991",
			x"0000" when x"B992",
			x"0000" when x"B993",
			x"0000" when x"B994",
			x"0000" when x"B995",
			x"0000" when x"B996",
			x"0000" when x"B997",
			x"0000" when x"B998",
			x"0000" when x"B999",
			x"0000" when x"B99A",
			x"0000" when x"B99B",
			x"0000" when x"B99C",
			x"0000" when x"B99D",
			x"0000" when x"B99E",
			x"0000" when x"B99F",
			x"0000" when x"B9A0",
			x"0000" when x"B9A1",
			x"0000" when x"B9A2",
			x"0000" when x"B9A3",
			x"0000" when x"B9A4",
			x"0000" when x"B9A5",
			x"0000" when x"B9A6",
			x"0000" when x"B9A7",
			x"0000" when x"B9A8",
			x"0000" when x"B9A9",
			x"0000" when x"B9AA",
			x"0000" when x"B9AB",
			x"0000" when x"B9AC",
			x"0000" when x"B9AD",
			x"0000" when x"B9AE",
			x"0000" when x"B9AF",
			x"0000" when x"B9B0",
			x"0000" when x"B9B1",
			x"0000" when x"B9B2",
			x"0000" when x"B9B3",
			x"0000" when x"B9B4",
			x"0000" when x"B9B5",
			x"0000" when x"B9B6",
			x"0000" when x"B9B7",
			x"0000" when x"B9B8",
			x"0000" when x"B9B9",
			x"0000" when x"B9BA",
			x"0000" when x"B9BB",
			x"0000" when x"B9BC",
			x"0000" when x"B9BD",
			x"0000" when x"B9BE",
			x"0000" when x"B9BF",
			x"0000" when x"B9C0",
			x"0000" when x"B9C1",
			x"0000" when x"B9C2",
			x"0000" when x"B9C3",
			x"0000" when x"B9C4",
			x"0000" when x"B9C5",
			x"0000" when x"B9C6",
			x"0000" when x"B9C7",
			x"0000" when x"B9C8",
			x"0000" when x"B9C9",
			x"0000" when x"B9CA",
			x"0000" when x"B9CB",
			x"0000" when x"B9CC",
			x"0000" when x"B9CD",
			x"0000" when x"B9CE",
			x"0000" when x"B9CF",
			x"0000" when x"B9D0",
			x"0000" when x"B9D1",
			x"0000" when x"B9D2",
			x"0000" when x"B9D3",
			x"0000" when x"B9D4",
			x"0000" when x"B9D5",
			x"0000" when x"B9D6",
			x"0000" when x"B9D7",
			x"0000" when x"B9D8",
			x"0000" when x"B9D9",
			x"0000" when x"B9DA",
			x"0000" when x"B9DB",
			x"0000" when x"B9DC",
			x"0000" when x"B9DD",
			x"0000" when x"B9DE",
			x"0000" when x"B9DF",
			x"0000" when x"B9E0",
			x"0000" when x"B9E1",
			x"0000" when x"B9E2",
			x"0000" when x"B9E3",
			x"0000" when x"B9E4",
			x"0000" when x"B9E5",
			x"0000" when x"B9E6",
			x"0000" when x"B9E7",
			x"0000" when x"B9E8",
			x"0000" when x"B9E9",
			x"0000" when x"B9EA",
			x"0000" when x"B9EB",
			x"0000" when x"B9EC",
			x"0000" when x"B9ED",
			x"0000" when x"B9EE",
			x"0000" when x"B9EF",
			x"0000" when x"B9F0",
			x"0000" when x"B9F1",
			x"0000" when x"B9F2",
			x"0000" when x"B9F3",
			x"0000" when x"B9F4",
			x"0000" when x"B9F5",
			x"0000" when x"B9F6",
			x"0000" when x"B9F7",
			x"0000" when x"B9F8",
			x"0000" when x"B9F9",
			x"0000" when x"B9FA",
			x"0000" when x"B9FB",
			x"0000" when x"B9FC",
			x"0000" when x"B9FD",
			x"0000" when x"B9FE",
			x"0000" when x"B9FF",
			x"0000" when x"BA00",
			x"0000" when x"BA01",
			x"0000" when x"BA02",
			x"0000" when x"BA03",
			x"0000" when x"BA04",
			x"0000" when x"BA05",
			x"0000" when x"BA06",
			x"0000" when x"BA07",
			x"0000" when x"BA08",
			x"0000" when x"BA09",
			x"0000" when x"BA0A",
			x"0000" when x"BA0B",
			x"0000" when x"BA0C",
			x"0000" when x"BA0D",
			x"0000" when x"BA0E",
			x"0000" when x"BA0F",
			x"0000" when x"BA10",
			x"0000" when x"BA11",
			x"0000" when x"BA12",
			x"0000" when x"BA13",
			x"0000" when x"BA14",
			x"0000" when x"BA15",
			x"0000" when x"BA16",
			x"0000" when x"BA17",
			x"0000" when x"BA18",
			x"0000" when x"BA19",
			x"0000" when x"BA1A",
			x"0000" when x"BA1B",
			x"0000" when x"BA1C",
			x"0000" when x"BA1D",
			x"0000" when x"BA1E",
			x"0000" when x"BA1F",
			x"0000" when x"BA20",
			x"0000" when x"BA21",
			x"0000" when x"BA22",
			x"0000" when x"BA23",
			x"0000" when x"BA24",
			x"0000" when x"BA25",
			x"0000" when x"BA26",
			x"0000" when x"BA27",
			x"0000" when x"BA28",
			x"0000" when x"BA29",
			x"0000" when x"BA2A",
			x"0000" when x"BA2B",
			x"0000" when x"BA2C",
			x"0000" when x"BA2D",
			x"0000" when x"BA2E",
			x"0000" when x"BA2F",
			x"0000" when x"BA30",
			x"0000" when x"BA31",
			x"0000" when x"BA32",
			x"0000" when x"BA33",
			x"0000" when x"BA34",
			x"0000" when x"BA35",
			x"0000" when x"BA36",
			x"0000" when x"BA37",
			x"0000" when x"BA38",
			x"0000" when x"BA39",
			x"0000" when x"BA3A",
			x"0000" when x"BA3B",
			x"0000" when x"BA3C",
			x"0000" when x"BA3D",
			x"0000" when x"BA3E",
			x"0000" when x"BA3F",
			x"0000" when x"BA40",
			x"0000" when x"BA41",
			x"0000" when x"BA42",
			x"0000" when x"BA43",
			x"0000" when x"BA44",
			x"0000" when x"BA45",
			x"0000" when x"BA46",
			x"0000" when x"BA47",
			x"0000" when x"BA48",
			x"0000" when x"BA49",
			x"0000" when x"BA4A",
			x"0000" when x"BA4B",
			x"0000" when x"BA4C",
			x"0000" when x"BA4D",
			x"0000" when x"BA4E",
			x"0000" when x"BA4F",
			x"0000" when x"BA50",
			x"0000" when x"BA51",
			x"0000" when x"BA52",
			x"0000" when x"BA53",
			x"0000" when x"BA54",
			x"0000" when x"BA55",
			x"0000" when x"BA56",
			x"0000" when x"BA57",
			x"0000" when x"BA58",
			x"0000" when x"BA59",
			x"0000" when x"BA5A",
			x"0000" when x"BA5B",
			x"0000" when x"BA5C",
			x"0000" when x"BA5D",
			x"0000" when x"BA5E",
			x"0000" when x"BA5F",
			x"0000" when x"BA60",
			x"0000" when x"BA61",
			x"0000" when x"BA62",
			x"0000" when x"BA63",
			x"0000" when x"BA64",
			x"0000" when x"BA65",
			x"0000" when x"BA66",
			x"0000" when x"BA67",
			x"0000" when x"BA68",
			x"0000" when x"BA69",
			x"0000" when x"BA6A",
			x"0000" when x"BA6B",
			x"0000" when x"BA6C",
			x"0000" when x"BA6D",
			x"0000" when x"BA6E",
			x"0000" when x"BA6F",
			x"0000" when x"BA70",
			x"0000" when x"BA71",
			x"0000" when x"BA72",
			x"0000" when x"BA73",
			x"0000" when x"BA74",
			x"0000" when x"BA75",
			x"0000" when x"BA76",
			x"0000" when x"BA77",
			x"0000" when x"BA78",
			x"0000" when x"BA79",
			x"0000" when x"BA7A",
			x"0000" when x"BA7B",
			x"0000" when x"BA7C",
			x"0000" when x"BA7D",
			x"0000" when x"BA7E",
			x"0000" when x"BA7F",
			x"0000" when x"BA80",
			x"0000" when x"BA81",
			x"0000" when x"BA82",
			x"0000" when x"BA83",
			x"0000" when x"BA84",
			x"0000" when x"BA85",
			x"0000" when x"BA86",
			x"0000" when x"BA87",
			x"0000" when x"BA88",
			x"0000" when x"BA89",
			x"0000" when x"BA8A",
			x"0000" when x"BA8B",
			x"0000" when x"BA8C",
			x"0000" when x"BA8D",
			x"0000" when x"BA8E",
			x"0000" when x"BA8F",
			x"0000" when x"BA90",
			x"0000" when x"BA91",
			x"0000" when x"BA92",
			x"0000" when x"BA93",
			x"0000" when x"BA94",
			x"0000" when x"BA95",
			x"0000" when x"BA96",
			x"0000" when x"BA97",
			x"0000" when x"BA98",
			x"0000" when x"BA99",
			x"0000" when x"BA9A",
			x"0000" when x"BA9B",
			x"0000" when x"BA9C",
			x"0000" when x"BA9D",
			x"0000" when x"BA9E",
			x"0000" when x"BA9F",
			x"0000" when x"BAA0",
			x"0000" when x"BAA1",
			x"0000" when x"BAA2",
			x"0000" when x"BAA3",
			x"0000" when x"BAA4",
			x"0000" when x"BAA5",
			x"0000" when x"BAA6",
			x"0000" when x"BAA7",
			x"0000" when x"BAA8",
			x"0000" when x"BAA9",
			x"0000" when x"BAAA",
			x"0000" when x"BAAB",
			x"0000" when x"BAAC",
			x"0000" when x"BAAD",
			x"0000" when x"BAAE",
			x"0000" when x"BAAF",
			x"0000" when x"BAB0",
			x"0000" when x"BAB1",
			x"0000" when x"BAB2",
			x"0000" when x"BAB3",
			x"0000" when x"BAB4",
			x"0000" when x"BAB5",
			x"0000" when x"BAB6",
			x"0000" when x"BAB7",
			x"0000" when x"BAB8",
			x"0000" when x"BAB9",
			x"0000" when x"BABA",
			x"0000" when x"BABB",
			x"0000" when x"BABC",
			x"0000" when x"BABD",
			x"0000" when x"BABE",
			x"0000" when x"BABF",
			x"0000" when x"BAC0",
			x"0000" when x"BAC1",
			x"0000" when x"BAC2",
			x"0000" when x"BAC3",
			x"0000" when x"BAC4",
			x"0000" when x"BAC5",
			x"0000" when x"BAC6",
			x"0000" when x"BAC7",
			x"0000" when x"BAC8",
			x"0000" when x"BAC9",
			x"0000" when x"BACA",
			x"0000" when x"BACB",
			x"0000" when x"BACC",
			x"0000" when x"BACD",
			x"0000" when x"BACE",
			x"0000" when x"BACF",
			x"0000" when x"BAD0",
			x"0000" when x"BAD1",
			x"0000" when x"BAD2",
			x"0000" when x"BAD3",
			x"0000" when x"BAD4",
			x"0000" when x"BAD5",
			x"0000" when x"BAD6",
			x"0000" when x"BAD7",
			x"0000" when x"BAD8",
			x"0000" when x"BAD9",
			x"0000" when x"BADA",
			x"0000" when x"BADB",
			x"0000" when x"BADC",
			x"0000" when x"BADD",
			x"0000" when x"BADE",
			x"0000" when x"BADF",
			x"0000" when x"BAE0",
			x"0000" when x"BAE1",
			x"0000" when x"BAE2",
			x"0000" when x"BAE3",
			x"0000" when x"BAE4",
			x"0000" when x"BAE5",
			x"0000" when x"BAE6",
			x"0000" when x"BAE7",
			x"0000" when x"BAE8",
			x"0000" when x"BAE9",
			x"0000" when x"BAEA",
			x"0000" when x"BAEB",
			x"0000" when x"BAEC",
			x"0000" when x"BAED",
			x"0000" when x"BAEE",
			x"0000" when x"BAEF",
			x"0000" when x"BAF0",
			x"0000" when x"BAF1",
			x"0000" when x"BAF2",
			x"0000" when x"BAF3",
			x"0000" when x"BAF4",
			x"0000" when x"BAF5",
			x"0000" when x"BAF6",
			x"0000" when x"BAF7",
			x"0000" when x"BAF8",
			x"0000" when x"BAF9",
			x"0000" when x"BAFA",
			x"0000" when x"BAFB",
			x"0000" when x"BAFC",
			x"0000" when x"BAFD",
			x"0000" when x"BAFE",
			x"0000" when x"BAFF",
			x"0000" when x"BB00",
			x"0000" when x"BB01",
			x"0000" when x"BB02",
			x"0000" when x"BB03",
			x"0000" when x"BB04",
			x"0000" when x"BB05",
			x"0000" when x"BB06",
			x"0000" when x"BB07",
			x"0000" when x"BB08",
			x"0000" when x"BB09",
			x"0000" when x"BB0A",
			x"0000" when x"BB0B",
			x"0000" when x"BB0C",
			x"0000" when x"BB0D",
			x"0000" when x"BB0E",
			x"0000" when x"BB0F",
			x"0000" when x"BB10",
			x"0000" when x"BB11",
			x"0000" when x"BB12",
			x"0000" when x"BB13",
			x"0000" when x"BB14",
			x"0000" when x"BB15",
			x"0000" when x"BB16",
			x"0000" when x"BB17",
			x"0000" when x"BB18",
			x"0000" when x"BB19",
			x"0000" when x"BB1A",
			x"0000" when x"BB1B",
			x"0000" when x"BB1C",
			x"0000" when x"BB1D",
			x"0000" when x"BB1E",
			x"0000" when x"BB1F",
			x"0000" when x"BB20",
			x"0000" when x"BB21",
			x"0000" when x"BB22",
			x"0000" when x"BB23",
			x"0000" when x"BB24",
			x"0000" when x"BB25",
			x"0000" when x"BB26",
			x"0000" when x"BB27",
			x"0000" when x"BB28",
			x"0000" when x"BB29",
			x"0000" when x"BB2A",
			x"0000" when x"BB2B",
			x"0000" when x"BB2C",
			x"0000" when x"BB2D",
			x"0000" when x"BB2E",
			x"0000" when x"BB2F",
			x"0000" when x"BB30",
			x"0000" when x"BB31",
			x"0000" when x"BB32",
			x"0000" when x"BB33",
			x"0000" when x"BB34",
			x"0000" when x"BB35",
			x"0000" when x"BB36",
			x"0000" when x"BB37",
			x"0000" when x"BB38",
			x"0000" when x"BB39",
			x"0000" when x"BB3A",
			x"0000" when x"BB3B",
			x"0000" when x"BB3C",
			x"0000" when x"BB3D",
			x"0000" when x"BB3E",
			x"0000" when x"BB3F",
			x"0000" when x"BB40",
			x"0000" when x"BB41",
			x"0000" when x"BB42",
			x"0000" when x"BB43",
			x"0000" when x"BB44",
			x"0000" when x"BB45",
			x"0000" when x"BB46",
			x"0000" when x"BB47",
			x"0000" when x"BB48",
			x"0000" when x"BB49",
			x"0000" when x"BB4A",
			x"0000" when x"BB4B",
			x"0000" when x"BB4C",
			x"0000" when x"BB4D",
			x"0000" when x"BB4E",
			x"0000" when x"BB4F",
			x"0000" when x"BB50",
			x"0000" when x"BB51",
			x"0000" when x"BB52",
			x"0000" when x"BB53",
			x"0000" when x"BB54",
			x"0000" when x"BB55",
			x"0000" when x"BB56",
			x"0000" when x"BB57",
			x"0000" when x"BB58",
			x"0000" when x"BB59",
			x"0000" when x"BB5A",
			x"0000" when x"BB5B",
			x"0000" when x"BB5C",
			x"0000" when x"BB5D",
			x"0000" when x"BB5E",
			x"0000" when x"BB5F",
			x"0000" when x"BB60",
			x"0000" when x"BB61",
			x"0000" when x"BB62",
			x"0000" when x"BB63",
			x"0000" when x"BB64",
			x"0000" when x"BB65",
			x"0000" when x"BB66",
			x"0000" when x"BB67",
			x"0000" when x"BB68",
			x"0000" when x"BB69",
			x"0000" when x"BB6A",
			x"0000" when x"BB6B",
			x"0000" when x"BB6C",
			x"0000" when x"BB6D",
			x"0000" when x"BB6E",
			x"0000" when x"BB6F",
			x"0000" when x"BB70",
			x"0000" when x"BB71",
			x"0000" when x"BB72",
			x"0000" when x"BB73",
			x"0000" when x"BB74",
			x"0000" when x"BB75",
			x"0000" when x"BB76",
			x"0000" when x"BB77",
			x"0000" when x"BB78",
			x"0000" when x"BB79",
			x"0000" when x"BB7A",
			x"0000" when x"BB7B",
			x"0000" when x"BB7C",
			x"0000" when x"BB7D",
			x"0000" when x"BB7E",
			x"0000" when x"BB7F",
			x"0000" when x"BB80",
			x"0000" when x"BB81",
			x"0000" when x"BB82",
			x"0000" when x"BB83",
			x"0000" when x"BB84",
			x"0000" when x"BB85",
			x"0000" when x"BB86",
			x"0000" when x"BB87",
			x"0000" when x"BB88",
			x"0000" when x"BB89",
			x"0000" when x"BB8A",
			x"0000" when x"BB8B",
			x"0000" when x"BB8C",
			x"0000" when x"BB8D",
			x"0000" when x"BB8E",
			x"0000" when x"BB8F",
			x"0000" when x"BB90",
			x"0000" when x"BB91",
			x"0000" when x"BB92",
			x"0000" when x"BB93",
			x"0000" when x"BB94",
			x"0000" when x"BB95",
			x"0000" when x"BB96",
			x"0000" when x"BB97",
			x"0000" when x"BB98",
			x"0000" when x"BB99",
			x"0000" when x"BB9A",
			x"0000" when x"BB9B",
			x"0000" when x"BB9C",
			x"0000" when x"BB9D",
			x"0000" when x"BB9E",
			x"0000" when x"BB9F",
			x"0000" when x"BBA0",
			x"0000" when x"BBA1",
			x"0000" when x"BBA2",
			x"0000" when x"BBA3",
			x"0000" when x"BBA4",
			x"0000" when x"BBA5",
			x"0000" when x"BBA6",
			x"0000" when x"BBA7",
			x"0000" when x"BBA8",
			x"0000" when x"BBA9",
			x"0000" when x"BBAA",
			x"0000" when x"BBAB",
			x"0000" when x"BBAC",
			x"0000" when x"BBAD",
			x"0000" when x"BBAE",
			x"0000" when x"BBAF",
			x"0000" when x"BBB0",
			x"0000" when x"BBB1",
			x"0000" when x"BBB2",
			x"0000" when x"BBB3",
			x"0000" when x"BBB4",
			x"0000" when x"BBB5",
			x"0000" when x"BBB6",
			x"0000" when x"BBB7",
			x"0000" when x"BBB8",
			x"0000" when x"BBB9",
			x"0000" when x"BBBA",
			x"0000" when x"BBBB",
			x"0000" when x"BBBC",
			x"0000" when x"BBBD",
			x"0000" when x"BBBE",
			x"0000" when x"BBBF",
			x"0000" when x"BBC0",
			x"0000" when x"BBC1",
			x"0000" when x"BBC2",
			x"0000" when x"BBC3",
			x"0000" when x"BBC4",
			x"0000" when x"BBC5",
			x"0000" when x"BBC6",
			x"0000" when x"BBC7",
			x"0000" when x"BBC8",
			x"0000" when x"BBC9",
			x"0000" when x"BBCA",
			x"0000" when x"BBCB",
			x"0000" when x"BBCC",
			x"0000" when x"BBCD",
			x"0000" when x"BBCE",
			x"0000" when x"BBCF",
			x"0000" when x"BBD0",
			x"0000" when x"BBD1",
			x"0000" when x"BBD2",
			x"0000" when x"BBD3",
			x"0000" when x"BBD4",
			x"0000" when x"BBD5",
			x"0000" when x"BBD6",
			x"0000" when x"BBD7",
			x"0000" when x"BBD8",
			x"0000" when x"BBD9",
			x"0000" when x"BBDA",
			x"0000" when x"BBDB",
			x"0000" when x"BBDC",
			x"0000" when x"BBDD",
			x"0000" when x"BBDE",
			x"0000" when x"BBDF",
			x"0000" when x"BBE0",
			x"0000" when x"BBE1",
			x"0000" when x"BBE2",
			x"0000" when x"BBE3",
			x"0000" when x"BBE4",
			x"0000" when x"BBE5",
			x"0000" when x"BBE6",
			x"0000" when x"BBE7",
			x"0000" when x"BBE8",
			x"0000" when x"BBE9",
			x"0000" when x"BBEA",
			x"0000" when x"BBEB",
			x"0000" when x"BBEC",
			x"0000" when x"BBED",
			x"0000" when x"BBEE",
			x"0000" when x"BBEF",
			x"0000" when x"BBF0",
			x"0000" when x"BBF1",
			x"0000" when x"BBF2",
			x"0000" when x"BBF3",
			x"0000" when x"BBF4",
			x"0000" when x"BBF5",
			x"0000" when x"BBF6",
			x"0000" when x"BBF7",
			x"0000" when x"BBF8",
			x"0000" when x"BBF9",
			x"0000" when x"BBFA",
			x"0000" when x"BBFB",
			x"0000" when x"BBFC",
			x"0000" when x"BBFD",
			x"0000" when x"BBFE",
			x"0000" when x"BBFF",
			x"0000" when x"BC00",
			x"0000" when x"BC01",
			x"0000" when x"BC02",
			x"0000" when x"BC03",
			x"0000" when x"BC04",
			x"0000" when x"BC05",
			x"0000" when x"BC06",
			x"0000" when x"BC07",
			x"0000" when x"BC08",
			x"0000" when x"BC09",
			x"0000" when x"BC0A",
			x"0000" when x"BC0B",
			x"0000" when x"BC0C",
			x"0000" when x"BC0D",
			x"0000" when x"BC0E",
			x"0000" when x"BC0F",
			x"0000" when x"BC10",
			x"0000" when x"BC11",
			x"0000" when x"BC12",
			x"0000" when x"BC13",
			x"0000" when x"BC14",
			x"0000" when x"BC15",
			x"0000" when x"BC16",
			x"0000" when x"BC17",
			x"0000" when x"BC18",
			x"0000" when x"BC19",
			x"0000" when x"BC1A",
			x"0000" when x"BC1B",
			x"0000" when x"BC1C",
			x"0000" when x"BC1D",
			x"0000" when x"BC1E",
			x"0000" when x"BC1F",
			x"0000" when x"BC20",
			x"0000" when x"BC21",
			x"0000" when x"BC22",
			x"0000" when x"BC23",
			x"0000" when x"BC24",
			x"0000" when x"BC25",
			x"0000" when x"BC26",
			x"0000" when x"BC27",
			x"0000" when x"BC28",
			x"0000" when x"BC29",
			x"0000" when x"BC2A",
			x"0000" when x"BC2B",
			x"0000" when x"BC2C",
			x"0000" when x"BC2D",
			x"0000" when x"BC2E",
			x"0000" when x"BC2F",
			x"0000" when x"BC30",
			x"0000" when x"BC31",
			x"0000" when x"BC32",
			x"0000" when x"BC33",
			x"0000" when x"BC34",
			x"0000" when x"BC35",
			x"0000" when x"BC36",
			x"0000" when x"BC37",
			x"0000" when x"BC38",
			x"0000" when x"BC39",
			x"0000" when x"BC3A",
			x"0000" when x"BC3B",
			x"0000" when x"BC3C",
			x"0000" when x"BC3D",
			x"0000" when x"BC3E",
			x"0000" when x"BC3F",
			x"0000" when x"BC40",
			x"0000" when x"BC41",
			x"0000" when x"BC42",
			x"0000" when x"BC43",
			x"0000" when x"BC44",
			x"0000" when x"BC45",
			x"0000" when x"BC46",
			x"0000" when x"BC47",
			x"0000" when x"BC48",
			x"0000" when x"BC49",
			x"0000" when x"BC4A",
			x"0000" when x"BC4B",
			x"0000" when x"BC4C",
			x"0000" when x"BC4D",
			x"0000" when x"BC4E",
			x"0000" when x"BC4F",
			x"0000" when x"BC50",
			x"0000" when x"BC51",
			x"0000" when x"BC52",
			x"0000" when x"BC53",
			x"0000" when x"BC54",
			x"0000" when x"BC55",
			x"0000" when x"BC56",
			x"0000" when x"BC57",
			x"0000" when x"BC58",
			x"0000" when x"BC59",
			x"0000" when x"BC5A",
			x"0000" when x"BC5B",
			x"0000" when x"BC5C",
			x"0000" when x"BC5D",
			x"0000" when x"BC5E",
			x"0000" when x"BC5F",
			x"0000" when x"BC60",
			x"0000" when x"BC61",
			x"0000" when x"BC62",
			x"0000" when x"BC63",
			x"0000" when x"BC64",
			x"0000" when x"BC65",
			x"0000" when x"BC66",
			x"0000" when x"BC67",
			x"0000" when x"BC68",
			x"0000" when x"BC69",
			x"0000" when x"BC6A",
			x"0000" when x"BC6B",
			x"0000" when x"BC6C",
			x"0000" when x"BC6D",
			x"0000" when x"BC6E",
			x"0000" when x"BC6F",
			x"0000" when x"BC70",
			x"0000" when x"BC71",
			x"0000" when x"BC72",
			x"0000" when x"BC73",
			x"0000" when x"BC74",
			x"0000" when x"BC75",
			x"0000" when x"BC76",
			x"0000" when x"BC77",
			x"0000" when x"BC78",
			x"0000" when x"BC79",
			x"0000" when x"BC7A",
			x"0000" when x"BC7B",
			x"0000" when x"BC7C",
			x"0000" when x"BC7D",
			x"0000" when x"BC7E",
			x"0000" when x"BC7F",
			x"0000" when x"BC80",
			x"0000" when x"BC81",
			x"0000" when x"BC82",
			x"0000" when x"BC83",
			x"0000" when x"BC84",
			x"0000" when x"BC85",
			x"0000" when x"BC86",
			x"0000" when x"BC87",
			x"0000" when x"BC88",
			x"0000" when x"BC89",
			x"0000" when x"BC8A",
			x"0000" when x"BC8B",
			x"0000" when x"BC8C",
			x"0000" when x"BC8D",
			x"0000" when x"BC8E",
			x"0000" when x"BC8F",
			x"0000" when x"BC90",
			x"0000" when x"BC91",
			x"0000" when x"BC92",
			x"0000" when x"BC93",
			x"0000" when x"BC94",
			x"0000" when x"BC95",
			x"0000" when x"BC96",
			x"0000" when x"BC97",
			x"0000" when x"BC98",
			x"0000" when x"BC99",
			x"0000" when x"BC9A",
			x"0000" when x"BC9B",
			x"0000" when x"BC9C",
			x"0000" when x"BC9D",
			x"0000" when x"BC9E",
			x"0000" when x"BC9F",
			x"0000" when x"BCA0",
			x"0000" when x"BCA1",
			x"0000" when x"BCA2",
			x"0000" when x"BCA3",
			x"0000" when x"BCA4",
			x"0000" when x"BCA5",
			x"0000" when x"BCA6",
			x"0000" when x"BCA7",
			x"0000" when x"BCA8",
			x"0000" when x"BCA9",
			x"0000" when x"BCAA",
			x"0000" when x"BCAB",
			x"0000" when x"BCAC",
			x"0000" when x"BCAD",
			x"0000" when x"BCAE",
			x"0000" when x"BCAF",
			x"0000" when x"BCB0",
			x"0000" when x"BCB1",
			x"0000" when x"BCB2",
			x"0000" when x"BCB3",
			x"0000" when x"BCB4",
			x"0000" when x"BCB5",
			x"0000" when x"BCB6",
			x"0000" when x"BCB7",
			x"0000" when x"BCB8",
			x"0000" when x"BCB9",
			x"0000" when x"BCBA",
			x"0000" when x"BCBB",
			x"0000" when x"BCBC",
			x"0000" when x"BCBD",
			x"0000" when x"BCBE",
			x"0000" when x"BCBF",
			x"0000" when x"BCC0",
			x"0000" when x"BCC1",
			x"0000" when x"BCC2",
			x"0000" when x"BCC3",
			x"0000" when x"BCC4",
			x"0000" when x"BCC5",
			x"0000" when x"BCC6",
			x"0000" when x"BCC7",
			x"0000" when x"BCC8",
			x"0000" when x"BCC9",
			x"0000" when x"BCCA",
			x"0000" when x"BCCB",
			x"0000" when x"BCCC",
			x"0000" when x"BCCD",
			x"0000" when x"BCCE",
			x"0000" when x"BCCF",
			x"0000" when x"BCD0",
			x"0000" when x"BCD1",
			x"0000" when x"BCD2",
			x"0000" when x"BCD3",
			x"0000" when x"BCD4",
			x"0000" when x"BCD5",
			x"0000" when x"BCD6",
			x"0000" when x"BCD7",
			x"0000" when x"BCD8",
			x"0000" when x"BCD9",
			x"0000" when x"BCDA",
			x"0000" when x"BCDB",
			x"0000" when x"BCDC",
			x"0000" when x"BCDD",
			x"0000" when x"BCDE",
			x"0000" when x"BCDF",
			x"0000" when x"BCE0",
			x"0000" when x"BCE1",
			x"0000" when x"BCE2",
			x"0000" when x"BCE3",
			x"0000" when x"BCE4",
			x"0000" when x"BCE5",
			x"0000" when x"BCE6",
			x"0000" when x"BCE7",
			x"0000" when x"BCE8",
			x"0000" when x"BCE9",
			x"0000" when x"BCEA",
			x"0000" when x"BCEB",
			x"0000" when x"BCEC",
			x"0000" when x"BCED",
			x"0000" when x"BCEE",
			x"0000" when x"BCEF",
			x"0000" when x"BCF0",
			x"0000" when x"BCF1",
			x"0000" when x"BCF2",
			x"0000" when x"BCF3",
			x"0000" when x"BCF4",
			x"0000" when x"BCF5",
			x"0000" when x"BCF6",
			x"0000" when x"BCF7",
			x"0000" when x"BCF8",
			x"0000" when x"BCF9",
			x"0000" when x"BCFA",
			x"0000" when x"BCFB",
			x"0000" when x"BCFC",
			x"0000" when x"BCFD",
			x"0000" when x"BCFE",
			x"0000" when x"BCFF",
			x"0000" when x"BD00",
			x"0000" when x"BD01",
			x"0000" when x"BD02",
			x"0000" when x"BD03",
			x"0000" when x"BD04",
			x"0000" when x"BD05",
			x"0000" when x"BD06",
			x"0000" when x"BD07",
			x"0000" when x"BD08",
			x"0000" when x"BD09",
			x"0000" when x"BD0A",
			x"0000" when x"BD0B",
			x"0000" when x"BD0C",
			x"0000" when x"BD0D",
			x"0000" when x"BD0E",
			x"0000" when x"BD0F",
			x"0000" when x"BD10",
			x"0000" when x"BD11",
			x"0000" when x"BD12",
			x"0000" when x"BD13",
			x"0000" when x"BD14",
			x"0000" when x"BD15",
			x"0000" when x"BD16",
			x"0000" when x"BD17",
			x"0000" when x"BD18",
			x"0000" when x"BD19",
			x"0000" when x"BD1A",
			x"0000" when x"BD1B",
			x"0000" when x"BD1C",
			x"0000" when x"BD1D",
			x"0000" when x"BD1E",
			x"0000" when x"BD1F",
			x"0000" when x"BD20",
			x"0000" when x"BD21",
			x"0000" when x"BD22",
			x"0000" when x"BD23",
			x"0000" when x"BD24",
			x"0000" when x"BD25",
			x"0000" when x"BD26",
			x"0000" when x"BD27",
			x"0000" when x"BD28",
			x"0000" when x"BD29",
			x"0000" when x"BD2A",
			x"0000" when x"BD2B",
			x"0000" when x"BD2C",
			x"0000" when x"BD2D",
			x"0000" when x"BD2E",
			x"0000" when x"BD2F",
			x"0000" when x"BD30",
			x"0000" when x"BD31",
			x"0000" when x"BD32",
			x"0000" when x"BD33",
			x"0000" when x"BD34",
			x"0000" when x"BD35",
			x"0000" when x"BD36",
			x"0000" when x"BD37",
			x"0000" when x"BD38",
			x"0000" when x"BD39",
			x"0000" when x"BD3A",
			x"0000" when x"BD3B",
			x"0000" when x"BD3C",
			x"0000" when x"BD3D",
			x"0000" when x"BD3E",
			x"0000" when x"BD3F",
			x"0000" when x"BD40",
			x"0000" when x"BD41",
			x"0000" when x"BD42",
			x"0000" when x"BD43",
			x"0000" when x"BD44",
			x"0000" when x"BD45",
			x"0000" when x"BD46",
			x"0000" when x"BD47",
			x"0000" when x"BD48",
			x"0000" when x"BD49",
			x"0000" when x"BD4A",
			x"0000" when x"BD4B",
			x"0000" when x"BD4C",
			x"0000" when x"BD4D",
			x"0000" when x"BD4E",
			x"0000" when x"BD4F",
			x"0000" when x"BD50",
			x"0000" when x"BD51",
			x"0000" when x"BD52",
			x"0000" when x"BD53",
			x"0000" when x"BD54",
			x"0000" when x"BD55",
			x"0000" when x"BD56",
			x"0000" when x"BD57",
			x"0000" when x"BD58",
			x"0000" when x"BD59",
			x"0000" when x"BD5A",
			x"0000" when x"BD5B",
			x"0000" when x"BD5C",
			x"0000" when x"BD5D",
			x"0000" when x"BD5E",
			x"0000" when x"BD5F",
			x"0000" when x"BD60",
			x"0000" when x"BD61",
			x"0000" when x"BD62",
			x"0000" when x"BD63",
			x"0000" when x"BD64",
			x"0000" when x"BD65",
			x"0000" when x"BD66",
			x"0000" when x"BD67",
			x"0000" when x"BD68",
			x"0000" when x"BD69",
			x"0000" when x"BD6A",
			x"0000" when x"BD6B",
			x"0000" when x"BD6C",
			x"0000" when x"BD6D",
			x"0000" when x"BD6E",
			x"0000" when x"BD6F",
			x"0000" when x"BD70",
			x"0000" when x"BD71",
			x"0000" when x"BD72",
			x"0000" when x"BD73",
			x"0000" when x"BD74",
			x"0000" when x"BD75",
			x"0000" when x"BD76",
			x"0000" when x"BD77",
			x"0000" when x"BD78",
			x"0000" when x"BD79",
			x"0000" when x"BD7A",
			x"0000" when x"BD7B",
			x"0000" when x"BD7C",
			x"0000" when x"BD7D",
			x"0000" when x"BD7E",
			x"0000" when x"BD7F",
			x"0000" when x"BD80",
			x"0000" when x"BD81",
			x"0000" when x"BD82",
			x"0000" when x"BD83",
			x"0000" when x"BD84",
			x"0000" when x"BD85",
			x"0000" when x"BD86",
			x"0000" when x"BD87",
			x"0000" when x"BD88",
			x"0000" when x"BD89",
			x"0000" when x"BD8A",
			x"0000" when x"BD8B",
			x"0000" when x"BD8C",
			x"0000" when x"BD8D",
			x"0000" when x"BD8E",
			x"0000" when x"BD8F",
			x"0000" when x"BD90",
			x"0000" when x"BD91",
			x"0000" when x"BD92",
			x"0000" when x"BD93",
			x"0000" when x"BD94",
			x"0000" when x"BD95",
			x"0000" when x"BD96",
			x"0000" when x"BD97",
			x"0000" when x"BD98",
			x"0000" when x"BD99",
			x"0000" when x"BD9A",
			x"0000" when x"BD9B",
			x"0000" when x"BD9C",
			x"0000" when x"BD9D",
			x"0000" when x"BD9E",
			x"0000" when x"BD9F",
			x"0000" when x"BDA0",
			x"0000" when x"BDA1",
			x"0000" when x"BDA2",
			x"0000" when x"BDA3",
			x"0000" when x"BDA4",
			x"0000" when x"BDA5",
			x"0000" when x"BDA6",
			x"0000" when x"BDA7",
			x"0000" when x"BDA8",
			x"0000" when x"BDA9",
			x"0000" when x"BDAA",
			x"0000" when x"BDAB",
			x"0000" when x"BDAC",
			x"0000" when x"BDAD",
			x"0000" when x"BDAE",
			x"0000" when x"BDAF",
			x"0000" when x"BDB0",
			x"0000" when x"BDB1",
			x"0000" when x"BDB2",
			x"0000" when x"BDB3",
			x"0000" when x"BDB4",
			x"0000" when x"BDB5",
			x"0000" when x"BDB6",
			x"0000" when x"BDB7",
			x"0000" when x"BDB8",
			x"0000" when x"BDB9",
			x"0000" when x"BDBA",
			x"0000" when x"BDBB",
			x"0000" when x"BDBC",
			x"0000" when x"BDBD",
			x"0000" when x"BDBE",
			x"0000" when x"BDBF",
			x"0000" when x"BDC0",
			x"0000" when x"BDC1",
			x"0000" when x"BDC2",
			x"0000" when x"BDC3",
			x"0000" when x"BDC4",
			x"0000" when x"BDC5",
			x"0000" when x"BDC6",
			x"0000" when x"BDC7",
			x"0000" when x"BDC8",
			x"0000" when x"BDC9",
			x"0000" when x"BDCA",
			x"0000" when x"BDCB",
			x"0000" when x"BDCC",
			x"0000" when x"BDCD",
			x"0000" when x"BDCE",
			x"0000" when x"BDCF",
			x"0000" when x"BDD0",
			x"0000" when x"BDD1",
			x"0000" when x"BDD2",
			x"0000" when x"BDD3",
			x"0000" when x"BDD4",
			x"0000" when x"BDD5",
			x"0000" when x"BDD6",
			x"0000" when x"BDD7",
			x"0000" when x"BDD8",
			x"0000" when x"BDD9",
			x"0000" when x"BDDA",
			x"0000" when x"BDDB",
			x"0000" when x"BDDC",
			x"0000" when x"BDDD",
			x"0000" when x"BDDE",
			x"0000" when x"BDDF",
			x"0000" when x"BDE0",
			x"0000" when x"BDE1",
			x"0000" when x"BDE2",
			x"0000" when x"BDE3",
			x"0000" when x"BDE4",
			x"0000" when x"BDE5",
			x"0000" when x"BDE6",
			x"0000" when x"BDE7",
			x"0000" when x"BDE8",
			x"0000" when x"BDE9",
			x"0000" when x"BDEA",
			x"0000" when x"BDEB",
			x"0000" when x"BDEC",
			x"0000" when x"BDED",
			x"0000" when x"BDEE",
			x"0000" when x"BDEF",
			x"0000" when x"BDF0",
			x"0000" when x"BDF1",
			x"0000" when x"BDF2",
			x"0000" when x"BDF3",
			x"0000" when x"BDF4",
			x"0000" when x"BDF5",
			x"0000" when x"BDF6",
			x"0000" when x"BDF7",
			x"0000" when x"BDF8",
			x"0000" when x"BDF9",
			x"0000" when x"BDFA",
			x"0000" when x"BDFB",
			x"0000" when x"BDFC",
			x"0000" when x"BDFD",
			x"0000" when x"BDFE",
			x"0000" when x"BDFF",
			x"0000" when x"BE00",
			x"0000" when x"BE01",
			x"0000" when x"BE02",
			x"0000" when x"BE03",
			x"0000" when x"BE04",
			x"0000" when x"BE05",
			x"0000" when x"BE06",
			x"0000" when x"BE07",
			x"0000" when x"BE08",
			x"0000" when x"BE09",
			x"0000" when x"BE0A",
			x"0000" when x"BE0B",
			x"0000" when x"BE0C",
			x"0000" when x"BE0D",
			x"0000" when x"BE0E",
			x"0000" when x"BE0F",
			x"0000" when x"BE10",
			x"0000" when x"BE11",
			x"0000" when x"BE12",
			x"0000" when x"BE13",
			x"0000" when x"BE14",
			x"0000" when x"BE15",
			x"0000" when x"BE16",
			x"0000" when x"BE17",
			x"0000" when x"BE18",
			x"0000" when x"BE19",
			x"0000" when x"BE1A",
			x"0000" when x"BE1B",
			x"0000" when x"BE1C",
			x"0000" when x"BE1D",
			x"0000" when x"BE1E",
			x"0000" when x"BE1F",
			x"0000" when x"BE20",
			x"0000" when x"BE21",
			x"0000" when x"BE22",
			x"0000" when x"BE23",
			x"0000" when x"BE24",
			x"0000" when x"BE25",
			x"0000" when x"BE26",
			x"0000" when x"BE27",
			x"0000" when x"BE28",
			x"0000" when x"BE29",
			x"0000" when x"BE2A",
			x"0000" when x"BE2B",
			x"0000" when x"BE2C",
			x"0000" when x"BE2D",
			x"0000" when x"BE2E",
			x"0000" when x"BE2F",
			x"0000" when x"BE30",
			x"0000" when x"BE31",
			x"0000" when x"BE32",
			x"0000" when x"BE33",
			x"0000" when x"BE34",
			x"0000" when x"BE35",
			x"0000" when x"BE36",
			x"0000" when x"BE37",
			x"0000" when x"BE38",
			x"0000" when x"BE39",
			x"0000" when x"BE3A",
			x"0000" when x"BE3B",
			x"0000" when x"BE3C",
			x"0000" when x"BE3D",
			x"0000" when x"BE3E",
			x"0000" when x"BE3F",
			x"0000" when x"BE40",
			x"0000" when x"BE41",
			x"0000" when x"BE42",
			x"0000" when x"BE43",
			x"0000" when x"BE44",
			x"0000" when x"BE45",
			x"0000" when x"BE46",
			x"0000" when x"BE47",
			x"0000" when x"BE48",
			x"0000" when x"BE49",
			x"0000" when x"BE4A",
			x"0000" when x"BE4B",
			x"0000" when x"BE4C",
			x"0000" when x"BE4D",
			x"0000" when x"BE4E",
			x"0000" when x"BE4F",
			x"0000" when x"BE50",
			x"0000" when x"BE51",
			x"0000" when x"BE52",
			x"0000" when x"BE53",
			x"0000" when x"BE54",
			x"0000" when x"BE55",
			x"0000" when x"BE56",
			x"0000" when x"BE57",
			x"0000" when x"BE58",
			x"0000" when x"BE59",
			x"0000" when x"BE5A",
			x"0000" when x"BE5B",
			x"0000" when x"BE5C",
			x"0000" when x"BE5D",
			x"0000" when x"BE5E",
			x"0000" when x"BE5F",
			x"0000" when x"BE60",
			x"0000" when x"BE61",
			x"0000" when x"BE62",
			x"0000" when x"BE63",
			x"0000" when x"BE64",
			x"0000" when x"BE65",
			x"0000" when x"BE66",
			x"0000" when x"BE67",
			x"0000" when x"BE68",
			x"0000" when x"BE69",
			x"0000" when x"BE6A",
			x"0000" when x"BE6B",
			x"0000" when x"BE6C",
			x"0000" when x"BE6D",
			x"0000" when x"BE6E",
			x"0000" when x"BE6F",
			x"0000" when x"BE70",
			x"0000" when x"BE71",
			x"0000" when x"BE72",
			x"0000" when x"BE73",
			x"0000" when x"BE74",
			x"0000" when x"BE75",
			x"0000" when x"BE76",
			x"0000" when x"BE77",
			x"0000" when x"BE78",
			x"0000" when x"BE79",
			x"0000" when x"BE7A",
			x"0000" when x"BE7B",
			x"0000" when x"BE7C",
			x"0000" when x"BE7D",
			x"0000" when x"BE7E",
			x"0000" when x"BE7F",
			x"0000" when x"BE80",
			x"0000" when x"BE81",
			x"0000" when x"BE82",
			x"0000" when x"BE83",
			x"0000" when x"BE84",
			x"0000" when x"BE85",
			x"0000" when x"BE86",
			x"0000" when x"BE87",
			x"0000" when x"BE88",
			x"0000" when x"BE89",
			x"0000" when x"BE8A",
			x"0000" when x"BE8B",
			x"0000" when x"BE8C",
			x"0000" when x"BE8D",
			x"0000" when x"BE8E",
			x"0000" when x"BE8F",
			x"0000" when x"BE90",
			x"0000" when x"BE91",
			x"0000" when x"BE92",
			x"0000" when x"BE93",
			x"0000" when x"BE94",
			x"0000" when x"BE95",
			x"0000" when x"BE96",
			x"0000" when x"BE97",
			x"0000" when x"BE98",
			x"0000" when x"BE99",
			x"0000" when x"BE9A",
			x"0000" when x"BE9B",
			x"0000" when x"BE9C",
			x"0000" when x"BE9D",
			x"0000" when x"BE9E",
			x"0000" when x"BE9F",
			x"0000" when x"BEA0",
			x"0000" when x"BEA1",
			x"0000" when x"BEA2",
			x"0000" when x"BEA3",
			x"0000" when x"BEA4",
			x"0000" when x"BEA5",
			x"0000" when x"BEA6",
			x"0000" when x"BEA7",
			x"0000" when x"BEA8",
			x"0000" when x"BEA9",
			x"0000" when x"BEAA",
			x"0000" when x"BEAB",
			x"0000" when x"BEAC",
			x"0000" when x"BEAD",
			x"0000" when x"BEAE",
			x"0000" when x"BEAF",
			x"0000" when x"BEB0",
			x"0000" when x"BEB1",
			x"0000" when x"BEB2",
			x"0000" when x"BEB3",
			x"0000" when x"BEB4",
			x"0000" when x"BEB5",
			x"0000" when x"BEB6",
			x"0000" when x"BEB7",
			x"0000" when x"BEB8",
			x"0000" when x"BEB9",
			x"0000" when x"BEBA",
			x"0000" when x"BEBB",
			x"0000" when x"BEBC",
			x"0000" when x"BEBD",
			x"0000" when x"BEBE",
			x"0000" when x"BEBF",
			x"0000" when x"BEC0",
			x"0000" when x"BEC1",
			x"0000" when x"BEC2",
			x"0000" when x"BEC3",
			x"0000" when x"BEC4",
			x"0000" when x"BEC5",
			x"0000" when x"BEC6",
			x"0000" when x"BEC7",
			x"0000" when x"BEC8",
			x"0000" when x"BEC9",
			x"0000" when x"BECA",
			x"0000" when x"BECB",
			x"0000" when x"BECC",
			x"0000" when x"BECD",
			x"0000" when x"BECE",
			x"0000" when x"BECF",
			x"0000" when x"BED0",
			x"0000" when x"BED1",
			x"0000" when x"BED2",
			x"0000" when x"BED3",
			x"0000" when x"BED4",
			x"0000" when x"BED5",
			x"0000" when x"BED6",
			x"0000" when x"BED7",
			x"0000" when x"BED8",
			x"0000" when x"BED9",
			x"0000" when x"BEDA",
			x"0000" when x"BEDB",
			x"0000" when x"BEDC",
			x"0000" when x"BEDD",
			x"0000" when x"BEDE",
			x"0000" when x"BEDF",
			x"0000" when x"BEE0",
			x"0000" when x"BEE1",
			x"0000" when x"BEE2",
			x"0000" when x"BEE3",
			x"0000" when x"BEE4",
			x"0000" when x"BEE5",
			x"0000" when x"BEE6",
			x"0000" when x"BEE7",
			x"0000" when x"BEE8",
			x"0000" when x"BEE9",
			x"0000" when x"BEEA",
			x"0000" when x"BEEB",
			x"0000" when x"BEEC",
			x"0000" when x"BEED",
			x"0000" when x"BEEE",
			x"0000" when x"BEEF",
			x"0000" when x"BEF0",
			x"0000" when x"BEF1",
			x"0000" when x"BEF2",
			x"0000" when x"BEF3",
			x"0000" when x"BEF4",
			x"0000" when x"BEF5",
			x"0000" when x"BEF6",
			x"0000" when x"BEF7",
			x"0000" when x"BEF8",
			x"0000" when x"BEF9",
			x"0000" when x"BEFA",
			x"0000" when x"BEFB",
			x"0000" when x"BEFC",
			x"0000" when x"BEFD",
			x"0000" when x"BEFE",
			x"0000" when x"BEFF",
			x"0000" when x"BF00",
			x"0000" when x"BF01",
			x"0000" when x"BF02",
			x"0000" when x"BF03",
			x"0000" when x"BF04",
			x"0000" when x"BF05",
			x"0000" when x"BF06",
			x"0000" when x"BF07",
			x"0000" when x"BF08",
			x"0000" when x"BF09",
			x"0000" when x"BF0A",
			x"0000" when x"BF0B",
			x"0000" when x"BF0C",
			x"0000" when x"BF0D",
			x"0000" when x"BF0E",
			x"0000" when x"BF0F",
			x"0000" when x"BF10",
			x"0000" when x"BF11",
			x"0000" when x"BF12",
			x"0000" when x"BF13",
			x"0000" when x"BF14",
			x"0000" when x"BF15",
			x"0000" when x"BF16",
			x"0000" when x"BF17",
			x"0000" when x"BF18",
			x"0000" when x"BF19",
			x"0000" when x"BF1A",
			x"0000" when x"BF1B",
			x"0000" when x"BF1C",
			x"0000" when x"BF1D",
			x"0000" when x"BF1E",
			x"0000" when x"BF1F",
			x"0000" when x"BF20",
			x"0000" when x"BF21",
			x"0000" when x"BF22",
			x"0000" when x"BF23",
			x"0000" when x"BF24",
			x"0000" when x"BF25",
			x"0000" when x"BF26",
			x"0000" when x"BF27",
			x"0000" when x"BF28",
			x"0000" when x"BF29",
			x"0000" when x"BF2A",
			x"0000" when x"BF2B",
			x"0000" when x"BF2C",
			x"0000" when x"BF2D",
			x"0000" when x"BF2E",
			x"0000" when x"BF2F",
			x"0000" when x"BF30",
			x"0000" when x"BF31",
			x"0000" when x"BF32",
			x"0000" when x"BF33",
			x"0000" when x"BF34",
			x"0000" when x"BF35",
			x"0000" when x"BF36",
			x"0000" when x"BF37",
			x"0000" when x"BF38",
			x"0000" when x"BF39",
			x"0000" when x"BF3A",
			x"0000" when x"BF3B",
			x"0000" when x"BF3C",
			x"0000" when x"BF3D",
			x"0000" when x"BF3E",
			x"0000" when x"BF3F",
			x"0000" when x"BF40",
			x"0000" when x"BF41",
			x"0000" when x"BF42",
			x"0000" when x"BF43",
			x"0000" when x"BF44",
			x"0000" when x"BF45",
			x"0000" when x"BF46",
			x"0000" when x"BF47",
			x"0000" when x"BF48",
			x"0000" when x"BF49",
			x"0000" when x"BF4A",
			x"0000" when x"BF4B",
			x"0000" when x"BF4C",
			x"0000" when x"BF4D",
			x"0000" when x"BF4E",
			x"0000" when x"BF4F",
			x"0000" when x"BF50",
			x"0000" when x"BF51",
			x"0000" when x"BF52",
			x"0000" when x"BF53",
			x"0000" when x"BF54",
			x"0000" when x"BF55",
			x"0000" when x"BF56",
			x"0000" when x"BF57",
			x"0000" when x"BF58",
			x"0000" when x"BF59",
			x"0000" when x"BF5A",
			x"0000" when x"BF5B",
			x"0000" when x"BF5C",
			x"0000" when x"BF5D",
			x"0000" when x"BF5E",
			x"0000" when x"BF5F",
			x"0000" when x"BF60",
			x"0000" when x"BF61",
			x"0000" when x"BF62",
			x"0000" when x"BF63",
			x"0000" when x"BF64",
			x"0000" when x"BF65",
			x"0000" when x"BF66",
			x"0000" when x"BF67",
			x"0000" when x"BF68",
			x"0000" when x"BF69",
			x"0000" when x"BF6A",
			x"0000" when x"BF6B",
			x"0000" when x"BF6C",
			x"0000" when x"BF6D",
			x"0000" when x"BF6E",
			x"0000" when x"BF6F",
			x"0000" when x"BF70",
			x"0000" when x"BF71",
			x"0000" when x"BF72",
			x"0000" when x"BF73",
			x"0000" when x"BF74",
			x"0000" when x"BF75",
			x"0000" when x"BF76",
			x"0000" when x"BF77",
			x"0000" when x"BF78",
			x"0000" when x"BF79",
			x"0000" when x"BF7A",
			x"0000" when x"BF7B",
			x"0000" when x"BF7C",
			x"0000" when x"BF7D",
			x"0000" when x"BF7E",
			x"0000" when x"BF7F",
			x"0000" when x"BF80",
			x"0000" when x"BF81",
			x"0000" when x"BF82",
			x"0000" when x"BF83",
			x"0000" when x"BF84",
			x"0000" when x"BF85",
			x"0000" when x"BF86",
			x"0000" when x"BF87",
			x"0000" when x"BF88",
			x"0000" when x"BF89",
			x"0000" when x"BF8A",
			x"0000" when x"BF8B",
			x"0000" when x"BF8C",
			x"0000" when x"BF8D",
			x"0000" when x"BF8E",
			x"0000" when x"BF8F",
			x"0000" when x"BF90",
			x"0000" when x"BF91",
			x"0000" when x"BF92",
			x"0000" when x"BF93",
			x"0000" when x"BF94",
			x"0000" when x"BF95",
			x"0000" when x"BF96",
			x"0000" when x"BF97",
			x"0000" when x"BF98",
			x"0000" when x"BF99",
			x"0000" when x"BF9A",
			x"0000" when x"BF9B",
			x"0000" when x"BF9C",
			x"0000" when x"BF9D",
			x"0000" when x"BF9E",
			x"0000" when x"BF9F",
			x"0000" when x"BFA0",
			x"0000" when x"BFA1",
			x"0000" when x"BFA2",
			x"0000" when x"BFA3",
			x"0000" when x"BFA4",
			x"0000" when x"BFA5",
			x"0000" when x"BFA6",
			x"0000" when x"BFA7",
			x"0000" when x"BFA8",
			x"0000" when x"BFA9",
			x"0000" when x"BFAA",
			x"0000" when x"BFAB",
			x"0000" when x"BFAC",
			x"0000" when x"BFAD",
			x"0000" when x"BFAE",
			x"0000" when x"BFAF",
			x"0000" when x"BFB0",
			x"0000" when x"BFB1",
			x"0000" when x"BFB2",
			x"0000" when x"BFB3",
			x"0000" when x"BFB4",
			x"0000" when x"BFB5",
			x"0000" when x"BFB6",
			x"0000" when x"BFB7",
			x"0000" when x"BFB8",
			x"0000" when x"BFB9",
			x"0000" when x"BFBA",
			x"0000" when x"BFBB",
			x"0000" when x"BFBC",
			x"0000" when x"BFBD",
			x"0000" when x"BFBE",
			x"0000" when x"BFBF",
			x"0000" when x"BFC0",
			x"0000" when x"BFC1",
			x"0000" when x"BFC2",
			x"0000" when x"BFC3",
			x"0000" when x"BFC4",
			x"0000" when x"BFC5",
			x"0000" when x"BFC6",
			x"0000" when x"BFC7",
			x"0000" when x"BFC8",
			x"0000" when x"BFC9",
			x"0000" when x"BFCA",
			x"0000" when x"BFCB",
			x"0000" when x"BFCC",
			x"0000" when x"BFCD",
			x"0000" when x"BFCE",
			x"0000" when x"BFCF",
			x"0000" when x"BFD0",
			x"0000" when x"BFD1",
			x"0000" when x"BFD2",
			x"0000" when x"BFD3",
			x"0000" when x"BFD4",
			x"0000" when x"BFD5",
			x"0000" when x"BFD6",
			x"0000" when x"BFD7",
			x"0000" when x"BFD8",
			x"0000" when x"BFD9",
			x"0000" when x"BFDA",
			x"0000" when x"BFDB",
			x"0000" when x"BFDC",
			x"0000" when x"BFDD",
			x"0000" when x"BFDE",
			x"0000" when x"BFDF",
			x"0000" when x"BFE0",
			x"0000" when x"BFE1",
			x"0000" when x"BFE2",
			x"0000" when x"BFE3",
			x"0000" when x"BFE4",
			x"0000" when x"BFE5",
			x"0000" when x"BFE6",
			x"0000" when x"BFE7",
			x"0000" when x"BFE8",
			x"0000" when x"BFE9",
			x"0000" when x"BFEA",
			x"0000" when x"BFEB",
			x"0000" when x"BFEC",
			x"0000" when x"BFED",
			x"0000" when x"BFEE",
			x"0000" when x"BFEF",
			x"0000" when x"BFF0",
			x"0000" when x"BFF1",
			x"0000" when x"BFF2",
			x"0000" when x"BFF3",
			x"0000" when x"BFF4",
			x"0000" when x"BFF5",
			x"0000" when x"BFF6",
			x"0000" when x"BFF7",
			x"0000" when x"BFF8",
			x"0000" when x"BFF9",
			x"0000" when x"BFFA",
			x"0000" when x"BFFB",
			x"0000" when x"BFFC",
			x"0000" when x"BFFD",
			x"0000" when x"BFFE",
			x"0000" when x"BFFF",
			x"0000" when x"C000",
			x"0000" when x"C001",
			x"0000" when x"C002",
			x"0000" when x"C003",
			x"0000" when x"C004",
			x"0000" when x"C005",
			x"0000" when x"C006",
			x"0000" when x"C007",
			x"0000" when x"C008",
			x"0000" when x"C009",
			x"0000" when x"C00A",
			x"0000" when x"C00B",
			x"0000" when x"C00C",
			x"0000" when x"C00D",
			x"0000" when x"C00E",
			x"0000" when x"C00F",
			x"0000" when x"C010",
			x"0000" when x"C011",
			x"0000" when x"C012",
			x"0000" when x"C013",
			x"0000" when x"C014",
			x"0000" when x"C015",
			x"0000" when x"C016",
			x"0000" when x"C017",
			x"0000" when x"C018",
			x"0000" when x"C019",
			x"0000" when x"C01A",
			x"0000" when x"C01B",
			x"0000" when x"C01C",
			x"0000" when x"C01D",
			x"0000" when x"C01E",
			x"0000" when x"C01F",
			x"0000" when x"C020",
			x"0000" when x"C021",
			x"0000" when x"C022",
			x"0000" when x"C023",
			x"0000" when x"C024",
			x"0000" when x"C025",
			x"0000" when x"C026",
			x"0000" when x"C027",
			x"0000" when x"C028",
			x"0000" when x"C029",
			x"0000" when x"C02A",
			x"0000" when x"C02B",
			x"0000" when x"C02C",
			x"0000" when x"C02D",
			x"0000" when x"C02E",
			x"0000" when x"C02F",
			x"0000" when x"C030",
			x"0000" when x"C031",
			x"0000" when x"C032",
			x"0000" when x"C033",
			x"0000" when x"C034",
			x"0000" when x"C035",
			x"0000" when x"C036",
			x"0000" when x"C037",
			x"0000" when x"C038",
			x"0000" when x"C039",
			x"0000" when x"C03A",
			x"0000" when x"C03B",
			x"0000" when x"C03C",
			x"0000" when x"C03D",
			x"0000" when x"C03E",
			x"0000" when x"C03F",
			x"0000" when x"C040",
			x"0000" when x"C041",
			x"0000" when x"C042",
			x"0000" when x"C043",
			x"0000" when x"C044",
			x"0000" when x"C045",
			x"0000" when x"C046",
			x"0000" when x"C047",
			x"0000" when x"C048",
			x"0000" when x"C049",
			x"0000" when x"C04A",
			x"0000" when x"C04B",
			x"0000" when x"C04C",
			x"0000" when x"C04D",
			x"0000" when x"C04E",
			x"0000" when x"C04F",
			x"0000" when x"C050",
			x"0000" when x"C051",
			x"0000" when x"C052",
			x"0000" when x"C053",
			x"0000" when x"C054",
			x"0000" when x"C055",
			x"0000" when x"C056",
			x"0000" when x"C057",
			x"0000" when x"C058",
			x"0000" when x"C059",
			x"0000" when x"C05A",
			x"0000" when x"C05B",
			x"0000" when x"C05C",
			x"0000" when x"C05D",
			x"0000" when x"C05E",
			x"0000" when x"C05F",
			x"0000" when x"C060",
			x"0000" when x"C061",
			x"0000" when x"C062",
			x"0000" when x"C063",
			x"0000" when x"C064",
			x"0000" when x"C065",
			x"0000" when x"C066",
			x"0000" when x"C067",
			x"0000" when x"C068",
			x"0000" when x"C069",
			x"0000" when x"C06A",
			x"0000" when x"C06B",
			x"0000" when x"C06C",
			x"0000" when x"C06D",
			x"0000" when x"C06E",
			x"0000" when x"C06F",
			x"0000" when x"C070",
			x"0000" when x"C071",
			x"0000" when x"C072",
			x"0000" when x"C073",
			x"0000" when x"C074",
			x"0000" when x"C075",
			x"0000" when x"C076",
			x"0000" when x"C077",
			x"0000" when x"C078",
			x"0000" when x"C079",
			x"0000" when x"C07A",
			x"0000" when x"C07B",
			x"0000" when x"C07C",
			x"0000" when x"C07D",
			x"0000" when x"C07E",
			x"0000" when x"C07F",
			x"0000" when x"C080",
			x"0000" when x"C081",
			x"0000" when x"C082",
			x"0000" when x"C083",
			x"0000" when x"C084",
			x"0000" when x"C085",
			x"0000" when x"C086",
			x"0000" when x"C087",
			x"0000" when x"C088",
			x"0000" when x"C089",
			x"0000" when x"C08A",
			x"0000" when x"C08B",
			x"0000" when x"C08C",
			x"0000" when x"C08D",
			x"0000" when x"C08E",
			x"0000" when x"C08F",
			x"0000" when x"C090",
			x"0000" when x"C091",
			x"0000" when x"C092",
			x"0000" when x"C093",
			x"0000" when x"C094",
			x"0000" when x"C095",
			x"0000" when x"C096",
			x"0000" when x"C097",
			x"0000" when x"C098",
			x"0000" when x"C099",
			x"0000" when x"C09A",
			x"0000" when x"C09B",
			x"0000" when x"C09C",
			x"0000" when x"C09D",
			x"0000" when x"C09E",
			x"0000" when x"C09F",
			x"0000" when x"C0A0",
			x"0000" when x"C0A1",
			x"0000" when x"C0A2",
			x"0000" when x"C0A3",
			x"0000" when x"C0A4",
			x"0000" when x"C0A5",
			x"0000" when x"C0A6",
			x"0000" when x"C0A7",
			x"0000" when x"C0A8",
			x"0000" when x"C0A9",
			x"0000" when x"C0AA",
			x"0000" when x"C0AB",
			x"0000" when x"C0AC",
			x"0000" when x"C0AD",
			x"0000" when x"C0AE",
			x"0000" when x"C0AF",
			x"0000" when x"C0B0",
			x"0000" when x"C0B1",
			x"0000" when x"C0B2",
			x"0000" when x"C0B3",
			x"0000" when x"C0B4",
			x"0000" when x"C0B5",
			x"0000" when x"C0B6",
			x"0000" when x"C0B7",
			x"0000" when x"C0B8",
			x"0000" when x"C0B9",
			x"0000" when x"C0BA",
			x"0000" when x"C0BB",
			x"0000" when x"C0BC",
			x"0000" when x"C0BD",
			x"0000" when x"C0BE",
			x"0000" when x"C0BF",
			x"0000" when x"C0C0",
			x"0000" when x"C0C1",
			x"0000" when x"C0C2",
			x"0000" when x"C0C3",
			x"0000" when x"C0C4",
			x"0000" when x"C0C5",
			x"0000" when x"C0C6",
			x"0000" when x"C0C7",
			x"0000" when x"C0C8",
			x"0000" when x"C0C9",
			x"0000" when x"C0CA",
			x"0000" when x"C0CB",
			x"0000" when x"C0CC",
			x"0000" when x"C0CD",
			x"0000" when x"C0CE",
			x"0000" when x"C0CF",
			x"0000" when x"C0D0",
			x"0000" when x"C0D1",
			x"0000" when x"C0D2",
			x"0000" when x"C0D3",
			x"0000" when x"C0D4",
			x"0000" when x"C0D5",
			x"0000" when x"C0D6",
			x"0000" when x"C0D7",
			x"0000" when x"C0D8",
			x"0000" when x"C0D9",
			x"0000" when x"C0DA",
			x"0000" when x"C0DB",
			x"0000" when x"C0DC",
			x"0000" when x"C0DD",
			x"0000" when x"C0DE",
			x"0000" when x"C0DF",
			x"0000" when x"C0E0",
			x"0000" when x"C0E1",
			x"0000" when x"C0E2",
			x"0000" when x"C0E3",
			x"0000" when x"C0E4",
			x"0000" when x"C0E5",
			x"0000" when x"C0E6",
			x"0000" when x"C0E7",
			x"0000" when x"C0E8",
			x"0000" when x"C0E9",
			x"0000" when x"C0EA",
			x"0000" when x"C0EB",
			x"0000" when x"C0EC",
			x"0000" when x"C0ED",
			x"0000" when x"C0EE",
			x"0000" when x"C0EF",
			x"0000" when x"C0F0",
			x"0000" when x"C0F1",
			x"0000" when x"C0F2",
			x"0000" when x"C0F3",
			x"0000" when x"C0F4",
			x"0000" when x"C0F5",
			x"0000" when x"C0F6",
			x"0000" when x"C0F7",
			x"0000" when x"C0F8",
			x"0000" when x"C0F9",
			x"0000" when x"C0FA",
			x"0000" when x"C0FB",
			x"0000" when x"C0FC",
			x"0000" when x"C0FD",
			x"0000" when x"C0FE",
			x"0000" when x"C0FF",
			x"0000" when x"C100",
			x"0000" when x"C101",
			x"0000" when x"C102",
			x"0000" when x"C103",
			x"0000" when x"C104",
			x"0000" when x"C105",
			x"0000" when x"C106",
			x"0000" when x"C107",
			x"0000" when x"C108",
			x"0000" when x"C109",
			x"0000" when x"C10A",
			x"0000" when x"C10B",
			x"0000" when x"C10C",
			x"0000" when x"C10D",
			x"0000" when x"C10E",
			x"0000" when x"C10F",
			x"0000" when x"C110",
			x"0000" when x"C111",
			x"0000" when x"C112",
			x"0000" when x"C113",
			x"0000" when x"C114",
			x"0000" when x"C115",
			x"0000" when x"C116",
			x"0000" when x"C117",
			x"0000" when x"C118",
			x"0000" when x"C119",
			x"0000" when x"C11A",
			x"0000" when x"C11B",
			x"0000" when x"C11C",
			x"0000" when x"C11D",
			x"0000" when x"C11E",
			x"0000" when x"C11F",
			x"0000" when x"C120",
			x"0000" when x"C121",
			x"0000" when x"C122",
			x"0000" when x"C123",
			x"0000" when x"C124",
			x"0000" when x"C125",
			x"0000" when x"C126",
			x"0000" when x"C127",
			x"0000" when x"C128",
			x"0000" when x"C129",
			x"0000" when x"C12A",
			x"0000" when x"C12B",
			x"0000" when x"C12C",
			x"0000" when x"C12D",
			x"0000" when x"C12E",
			x"0000" when x"C12F",
			x"0000" when x"C130",
			x"0000" when x"C131",
			x"0000" when x"C132",
			x"0000" when x"C133",
			x"0000" when x"C134",
			x"0000" when x"C135",
			x"0000" when x"C136",
			x"0000" when x"C137",
			x"0000" when x"C138",
			x"0000" when x"C139",
			x"0000" when x"C13A",
			x"0000" when x"C13B",
			x"0000" when x"C13C",
			x"0000" when x"C13D",
			x"0000" when x"C13E",
			x"0000" when x"C13F",
			x"0000" when x"C140",
			x"0000" when x"C141",
			x"0000" when x"C142",
			x"0000" when x"C143",
			x"0000" when x"C144",
			x"0000" when x"C145",
			x"0000" when x"C146",
			x"0000" when x"C147",
			x"0000" when x"C148",
			x"0000" when x"C149",
			x"0000" when x"C14A",
			x"0000" when x"C14B",
			x"0000" when x"C14C",
			x"0000" when x"C14D",
			x"0000" when x"C14E",
			x"0000" when x"C14F",
			x"0000" when x"C150",
			x"0000" when x"C151",
			x"0000" when x"C152",
			x"0000" when x"C153",
			x"0000" when x"C154",
			x"0000" when x"C155",
			x"0000" when x"C156",
			x"0000" when x"C157",
			x"0000" when x"C158",
			x"0000" when x"C159",
			x"0000" when x"C15A",
			x"0000" when x"C15B",
			x"0000" when x"C15C",
			x"0000" when x"C15D",
			x"0000" when x"C15E",
			x"0000" when x"C15F",
			x"0000" when x"C160",
			x"0000" when x"C161",
			x"0000" when x"C162",
			x"0000" when x"C163",
			x"0000" when x"C164",
			x"0000" when x"C165",
			x"0000" when x"C166",
			x"0000" when x"C167",
			x"0000" when x"C168",
			x"0000" when x"C169",
			x"0000" when x"C16A",
			x"0000" when x"C16B",
			x"0000" when x"C16C",
			x"0000" when x"C16D",
			x"0000" when x"C16E",
			x"0000" when x"C16F",
			x"0000" when x"C170",
			x"0000" when x"C171",
			x"0000" when x"C172",
			x"0000" when x"C173",
			x"0000" when x"C174",
			x"0000" when x"C175",
			x"0000" when x"C176",
			x"0000" when x"C177",
			x"0000" when x"C178",
			x"0000" when x"C179",
			x"0000" when x"C17A",
			x"0000" when x"C17B",
			x"0000" when x"C17C",
			x"0000" when x"C17D",
			x"0000" when x"C17E",
			x"0000" when x"C17F",
			x"0000" when x"C180",
			x"0000" when x"C181",
			x"0000" when x"C182",
			x"0000" when x"C183",
			x"0000" when x"C184",
			x"0000" when x"C185",
			x"0000" when x"C186",
			x"0000" when x"C187",
			x"0000" when x"C188",
			x"0000" when x"C189",
			x"0000" when x"C18A",
			x"0000" when x"C18B",
			x"0000" when x"C18C",
			x"0000" when x"C18D",
			x"0000" when x"C18E",
			x"0000" when x"C18F",
			x"0000" when x"C190",
			x"0000" when x"C191",
			x"0000" when x"C192",
			x"0000" when x"C193",
			x"0000" when x"C194",
			x"0000" when x"C195",
			x"0000" when x"C196",
			x"0000" when x"C197",
			x"0000" when x"C198",
			x"0000" when x"C199",
			x"0000" when x"C19A",
			x"0000" when x"C19B",
			x"0000" when x"C19C",
			x"0000" when x"C19D",
			x"0000" when x"C19E",
			x"0000" when x"C19F",
			x"0000" when x"C1A0",
			x"0000" when x"C1A1",
			x"0000" when x"C1A2",
			x"0000" when x"C1A3",
			x"0000" when x"C1A4",
			x"0000" when x"C1A5",
			x"0000" when x"C1A6",
			x"0000" when x"C1A7",
			x"0000" when x"C1A8",
			x"0000" when x"C1A9",
			x"0000" when x"C1AA",
			x"0000" when x"C1AB",
			x"0000" when x"C1AC",
			x"0000" when x"C1AD",
			x"0000" when x"C1AE",
			x"0000" when x"C1AF",
			x"0000" when x"C1B0",
			x"0000" when x"C1B1",
			x"0000" when x"C1B2",
			x"0000" when x"C1B3",
			x"0000" when x"C1B4",
			x"0000" when x"C1B5",
			x"0000" when x"C1B6",
			x"0000" when x"C1B7",
			x"0000" when x"C1B8",
			x"0000" when x"C1B9",
			x"0000" when x"C1BA",
			x"0000" when x"C1BB",
			x"0000" when x"C1BC",
			x"0000" when x"C1BD",
			x"0000" when x"C1BE",
			x"0000" when x"C1BF",
			x"0000" when x"C1C0",
			x"0000" when x"C1C1",
			x"0000" when x"C1C2",
			x"0000" when x"C1C3",
			x"0000" when x"C1C4",
			x"0000" when x"C1C5",
			x"0000" when x"C1C6",
			x"0000" when x"C1C7",
			x"0000" when x"C1C8",
			x"0000" when x"C1C9",
			x"0000" when x"C1CA",
			x"0000" when x"C1CB",
			x"0000" when x"C1CC",
			x"0000" when x"C1CD",
			x"0000" when x"C1CE",
			x"0000" when x"C1CF",
			x"0000" when x"C1D0",
			x"0000" when x"C1D1",
			x"0000" when x"C1D2",
			x"0000" when x"C1D3",
			x"0000" when x"C1D4",
			x"0000" when x"C1D5",
			x"0000" when x"C1D6",
			x"0000" when x"C1D7",
			x"0000" when x"C1D8",
			x"0000" when x"C1D9",
			x"0000" when x"C1DA",
			x"0000" when x"C1DB",
			x"0000" when x"C1DC",
			x"0000" when x"C1DD",
			x"0000" when x"C1DE",
			x"0000" when x"C1DF",
			x"0000" when x"C1E0",
			x"0000" when x"C1E1",
			x"0000" when x"C1E2",
			x"0000" when x"C1E3",
			x"0000" when x"C1E4",
			x"0000" when x"C1E5",
			x"0000" when x"C1E6",
			x"0000" when x"C1E7",
			x"0000" when x"C1E8",
			x"0000" when x"C1E9",
			x"0000" when x"C1EA",
			x"0000" when x"C1EB",
			x"0000" when x"C1EC",
			x"0000" when x"C1ED",
			x"0000" when x"C1EE",
			x"0000" when x"C1EF",
			x"0000" when x"C1F0",
			x"0000" when x"C1F1",
			x"0000" when x"C1F2",
			x"0000" when x"C1F3",
			x"0000" when x"C1F4",
			x"0000" when x"C1F5",
			x"0000" when x"C1F6",
			x"0000" when x"C1F7",
			x"0000" when x"C1F8",
			x"0000" when x"C1F9",
			x"0000" when x"C1FA",
			x"0000" when x"C1FB",
			x"0000" when x"C1FC",
			x"0000" when x"C1FD",
			x"0000" when x"C1FE",
			x"0000" when x"C1FF",
			x"0000" when x"C200",
			x"0000" when x"C201",
			x"0000" when x"C202",
			x"0000" when x"C203",
			x"0000" when x"C204",
			x"0000" when x"C205",
			x"0000" when x"C206",
			x"0000" when x"C207",
			x"0000" when x"C208",
			x"0000" when x"C209",
			x"0000" when x"C20A",
			x"0000" when x"C20B",
			x"0000" when x"C20C",
			x"0000" when x"C20D",
			x"0000" when x"C20E",
			x"0000" when x"C20F",
			x"0000" when x"C210",
			x"0000" when x"C211",
			x"0000" when x"C212",
			x"0000" when x"C213",
			x"0000" when x"C214",
			x"0000" when x"C215",
			x"0000" when x"C216",
			x"0000" when x"C217",
			x"0000" when x"C218",
			x"0000" when x"C219",
			x"0000" when x"C21A",
			x"0000" when x"C21B",
			x"0000" when x"C21C",
			x"0000" when x"C21D",
			x"0000" when x"C21E",
			x"0000" when x"C21F",
			x"0000" when x"C220",
			x"0000" when x"C221",
			x"0000" when x"C222",
			x"0000" when x"C223",
			x"0000" when x"C224",
			x"0000" when x"C225",
			x"0000" when x"C226",
			x"0000" when x"C227",
			x"0000" when x"C228",
			x"0000" when x"C229",
			x"0000" when x"C22A",
			x"0000" when x"C22B",
			x"0000" when x"C22C",
			x"0000" when x"C22D",
			x"0000" when x"C22E",
			x"0000" when x"C22F",
			x"0000" when x"C230",
			x"0000" when x"C231",
			x"0000" when x"C232",
			x"0000" when x"C233",
			x"0000" when x"C234",
			x"0000" when x"C235",
			x"0000" when x"C236",
			x"0000" when x"C237",
			x"0000" when x"C238",
			x"0000" when x"C239",
			x"0000" when x"C23A",
			x"0000" when x"C23B",
			x"0000" when x"C23C",
			x"0000" when x"C23D",
			x"0000" when x"C23E",
			x"0000" when x"C23F",
			x"0000" when x"C240",
			x"0000" when x"C241",
			x"0000" when x"C242",
			x"0000" when x"C243",
			x"0000" when x"C244",
			x"0000" when x"C245",
			x"0000" when x"C246",
			x"0000" when x"C247",
			x"0000" when x"C248",
			x"0000" when x"C249",
			x"0000" when x"C24A",
			x"0000" when x"C24B",
			x"0000" when x"C24C",
			x"0000" when x"C24D",
			x"0000" when x"C24E",
			x"0000" when x"C24F",
			x"0000" when x"C250",
			x"0000" when x"C251",
			x"0000" when x"C252",
			x"0000" when x"C253",
			x"0000" when x"C254",
			x"0000" when x"C255",
			x"0000" when x"C256",
			x"0000" when x"C257",
			x"0000" when x"C258",
			x"0000" when x"C259",
			x"0000" when x"C25A",
			x"0000" when x"C25B",
			x"0000" when x"C25C",
			x"0000" when x"C25D",
			x"0000" when x"C25E",
			x"0000" when x"C25F",
			x"0000" when x"C260",
			x"0000" when x"C261",
			x"0000" when x"C262",
			x"0000" when x"C263",
			x"0000" when x"C264",
			x"0000" when x"C265",
			x"0000" when x"C266",
			x"0000" when x"C267",
			x"0000" when x"C268",
			x"0000" when x"C269",
			x"0000" when x"C26A",
			x"0000" when x"C26B",
			x"0000" when x"C26C",
			x"0000" when x"C26D",
			x"0000" when x"C26E",
			x"0000" when x"C26F",
			x"0000" when x"C270",
			x"0000" when x"C271",
			x"0000" when x"C272",
			x"0000" when x"C273",
			x"0000" when x"C274",
			x"0000" when x"C275",
			x"0000" when x"C276",
			x"0000" when x"C277",
			x"0000" when x"C278",
			x"0000" when x"C279",
			x"0000" when x"C27A",
			x"0000" when x"C27B",
			x"0000" when x"C27C",
			x"0000" when x"C27D",
			x"0000" when x"C27E",
			x"0000" when x"C27F",
			x"0000" when x"C280",
			x"0000" when x"C281",
			x"0000" when x"C282",
			x"0000" when x"C283",
			x"0000" when x"C284",
			x"0000" when x"C285",
			x"0000" when x"C286",
			x"0000" when x"C287",
			x"0000" when x"C288",
			x"0000" when x"C289",
			x"0000" when x"C28A",
			x"0000" when x"C28B",
			x"0000" when x"C28C",
			x"0000" when x"C28D",
			x"0000" when x"C28E",
			x"0000" when x"C28F",
			x"0000" when x"C290",
			x"0000" when x"C291",
			x"0000" when x"C292",
			x"0000" when x"C293",
			x"0000" when x"C294",
			x"0000" when x"C295",
			x"0000" when x"C296",
			x"0000" when x"C297",
			x"0000" when x"C298",
			x"0000" when x"C299",
			x"0000" when x"C29A",
			x"0000" when x"C29B",
			x"0000" when x"C29C",
			x"0000" when x"C29D",
			x"0000" when x"C29E",
			x"0000" when x"C29F",
			x"0000" when x"C2A0",
			x"0000" when x"C2A1",
			x"0000" when x"C2A2",
			x"0000" when x"C2A3",
			x"0000" when x"C2A4",
			x"0000" when x"C2A5",
			x"0000" when x"C2A6",
			x"0000" when x"C2A7",
			x"0000" when x"C2A8",
			x"0000" when x"C2A9",
			x"0000" when x"C2AA",
			x"0000" when x"C2AB",
			x"0000" when x"C2AC",
			x"0000" when x"C2AD",
			x"0000" when x"C2AE",
			x"0000" when x"C2AF",
			x"0000" when x"C2B0",
			x"0000" when x"C2B1",
			x"0000" when x"C2B2",
			x"0000" when x"C2B3",
			x"0000" when x"C2B4",
			x"0000" when x"C2B5",
			x"0000" when x"C2B6",
			x"0000" when x"C2B7",
			x"0000" when x"C2B8",
			x"0000" when x"C2B9",
			x"0000" when x"C2BA",
			x"0000" when x"C2BB",
			x"0000" when x"C2BC",
			x"0000" when x"C2BD",
			x"0000" when x"C2BE",
			x"0000" when x"C2BF",
			x"0000" when x"C2C0",
			x"0000" when x"C2C1",
			x"0000" when x"C2C2",
			x"0000" when x"C2C3",
			x"0000" when x"C2C4",
			x"0000" when x"C2C5",
			x"0000" when x"C2C6",
			x"0000" when x"C2C7",
			x"0000" when x"C2C8",
			x"0000" when x"C2C9",
			x"0000" when x"C2CA",
			x"0000" when x"C2CB",
			x"0000" when x"C2CC",
			x"0000" when x"C2CD",
			x"0000" when x"C2CE",
			x"0000" when x"C2CF",
			x"0000" when x"C2D0",
			x"0000" when x"C2D1",
			x"0000" when x"C2D2",
			x"0000" when x"C2D3",
			x"0000" when x"C2D4",
			x"0000" when x"C2D5",
			x"0000" when x"C2D6",
			x"0000" when x"C2D7",
			x"0000" when x"C2D8",
			x"0000" when x"C2D9",
			x"0000" when x"C2DA",
			x"0000" when x"C2DB",
			x"0000" when x"C2DC",
			x"0000" when x"C2DD",
			x"0000" when x"C2DE",
			x"0000" when x"C2DF",
			x"0000" when x"C2E0",
			x"0000" when x"C2E1",
			x"0000" when x"C2E2",
			x"0000" when x"C2E3",
			x"0000" when x"C2E4",
			x"0000" when x"C2E5",
			x"0000" when x"C2E6",
			x"0000" when x"C2E7",
			x"0000" when x"C2E8",
			x"0000" when x"C2E9",
			x"0000" when x"C2EA",
			x"0000" when x"C2EB",
			x"0000" when x"C2EC",
			x"0000" when x"C2ED",
			x"0000" when x"C2EE",
			x"0000" when x"C2EF",
			x"0000" when x"C2F0",
			x"0000" when x"C2F1",
			x"0000" when x"C2F2",
			x"0000" when x"C2F3",
			x"0000" when x"C2F4",
			x"0000" when x"C2F5",
			x"0000" when x"C2F6",
			x"0000" when x"C2F7",
			x"0000" when x"C2F8",
			x"0000" when x"C2F9",
			x"0000" when x"C2FA",
			x"0000" when x"C2FB",
			x"0000" when x"C2FC",
			x"0000" when x"C2FD",
			x"0000" when x"C2FE",
			x"0000" when x"C2FF",
			x"0000" when x"C300",
			x"0000" when x"C301",
			x"0000" when x"C302",
			x"0000" when x"C303",
			x"0000" when x"C304",
			x"0000" when x"C305",
			x"0000" when x"C306",
			x"0000" when x"C307",
			x"0000" when x"C308",
			x"0000" when x"C309",
			x"0000" when x"C30A",
			x"0000" when x"C30B",
			x"0000" when x"C30C",
			x"0000" when x"C30D",
			x"0000" when x"C30E",
			x"0000" when x"C30F",
			x"0000" when x"C310",
			x"0000" when x"C311",
			x"0000" when x"C312",
			x"0000" when x"C313",
			x"0000" when x"C314",
			x"0000" when x"C315",
			x"0000" when x"C316",
			x"0000" when x"C317",
			x"0000" when x"C318",
			x"0000" when x"C319",
			x"0000" when x"C31A",
			x"0000" when x"C31B",
			x"0000" when x"C31C",
			x"0000" when x"C31D",
			x"0000" when x"C31E",
			x"0000" when x"C31F",
			x"0000" when x"C320",
			x"0000" when x"C321",
			x"0000" when x"C322",
			x"0000" when x"C323",
			x"0000" when x"C324",
			x"0000" when x"C325",
			x"0000" when x"C326",
			x"0000" when x"C327",
			x"0000" when x"C328",
			x"0000" when x"C329",
			x"0000" when x"C32A",
			x"0000" when x"C32B",
			x"0000" when x"C32C",
			x"0000" when x"C32D",
			x"0000" when x"C32E",
			x"0000" when x"C32F",
			x"0000" when x"C330",
			x"0000" when x"C331",
			x"0000" when x"C332",
			x"0000" when x"C333",
			x"0000" when x"C334",
			x"0000" when x"C335",
			x"0000" when x"C336",
			x"0000" when x"C337",
			x"0000" when x"C338",
			x"0000" when x"C339",
			x"0000" when x"C33A",
			x"0000" when x"C33B",
			x"0000" when x"C33C",
			x"0000" when x"C33D",
			x"0000" when x"C33E",
			x"0000" when x"C33F",
			x"0000" when x"C340",
			x"0000" when x"C341",
			x"0000" when x"C342",
			x"0000" when x"C343",
			x"0000" when x"C344",
			x"0000" when x"C345",
			x"0000" when x"C346",
			x"0000" when x"C347",
			x"0000" when x"C348",
			x"0000" when x"C349",
			x"0000" when x"C34A",
			x"0000" when x"C34B",
			x"0000" when x"C34C",
			x"0000" when x"C34D",
			x"0000" when x"C34E",
			x"0000" when x"C34F",
			x"0000" when x"C350",
			x"0000" when x"C351",
			x"0000" when x"C352",
			x"0000" when x"C353",
			x"0000" when x"C354",
			x"0000" when x"C355",
			x"0000" when x"C356",
			x"0000" when x"C357",
			x"0000" when x"C358",
			x"0000" when x"C359",
			x"0000" when x"C35A",
			x"0000" when x"C35B",
			x"0000" when x"C35C",
			x"0000" when x"C35D",
			x"0000" when x"C35E",
			x"0000" when x"C35F",
			x"0000" when x"C360",
			x"0000" when x"C361",
			x"0000" when x"C362",
			x"0000" when x"C363",
			x"0000" when x"C364",
			x"0000" when x"C365",
			x"0000" when x"C366",
			x"0000" when x"C367",
			x"0000" when x"C368",
			x"0000" when x"C369",
			x"0000" when x"C36A",
			x"0000" when x"C36B",
			x"0000" when x"C36C",
			x"0000" when x"C36D",
			x"0000" when x"C36E",
			x"0000" when x"C36F",
			x"0000" when x"C370",
			x"0000" when x"C371",
			x"0000" when x"C372",
			x"0000" when x"C373",
			x"0000" when x"C374",
			x"0000" when x"C375",
			x"0000" when x"C376",
			x"0000" when x"C377",
			x"0000" when x"C378",
			x"0000" when x"C379",
			x"0000" when x"C37A",
			x"0000" when x"C37B",
			x"0000" when x"C37C",
			x"0000" when x"C37D",
			x"0000" when x"C37E",
			x"0000" when x"C37F",
			x"0000" when x"C380",
			x"0000" when x"C381",
			x"0000" when x"C382",
			x"0000" when x"C383",
			x"0000" when x"C384",
			x"0000" when x"C385",
			x"0000" when x"C386",
			x"0000" when x"C387",
			x"0000" when x"C388",
			x"0000" when x"C389",
			x"0000" when x"C38A",
			x"0000" when x"C38B",
			x"0000" when x"C38C",
			x"0000" when x"C38D",
			x"0000" when x"C38E",
			x"0000" when x"C38F",
			x"0000" when x"C390",
			x"0000" when x"C391",
			x"0000" when x"C392",
			x"0000" when x"C393",
			x"0000" when x"C394",
			x"0000" when x"C395",
			x"0000" when x"C396",
			x"0000" when x"C397",
			x"0000" when x"C398",
			x"0000" when x"C399",
			x"0000" when x"C39A",
			x"0000" when x"C39B",
			x"0000" when x"C39C",
			x"0000" when x"C39D",
			x"0000" when x"C39E",
			x"0000" when x"C39F",
			x"0000" when x"C3A0",
			x"0000" when x"C3A1",
			x"0000" when x"C3A2",
			x"0000" when x"C3A3",
			x"0000" when x"C3A4",
			x"0000" when x"C3A5",
			x"0000" when x"C3A6",
			x"0000" when x"C3A7",
			x"0000" when x"C3A8",
			x"0000" when x"C3A9",
			x"0000" when x"C3AA",
			x"0000" when x"C3AB",
			x"0000" when x"C3AC",
			x"0000" when x"C3AD",
			x"0000" when x"C3AE",
			x"0000" when x"C3AF",
			x"0000" when x"C3B0",
			x"0000" when x"C3B1",
			x"0000" when x"C3B2",
			x"0000" when x"C3B3",
			x"0000" when x"C3B4",
			x"0000" when x"C3B5",
			x"0000" when x"C3B6",
			x"0000" when x"C3B7",
			x"0000" when x"C3B8",
			x"0000" when x"C3B9",
			x"0000" when x"C3BA",
			x"0000" when x"C3BB",
			x"0000" when x"C3BC",
			x"0000" when x"C3BD",
			x"0000" when x"C3BE",
			x"0000" when x"C3BF",
			x"0000" when x"C3C0",
			x"0000" when x"C3C1",
			x"0000" when x"C3C2",
			x"0000" when x"C3C3",
			x"0000" when x"C3C4",
			x"0000" when x"C3C5",
			x"0000" when x"C3C6",
			x"0000" when x"C3C7",
			x"0000" when x"C3C8",
			x"0000" when x"C3C9",
			x"0000" when x"C3CA",
			x"0000" when x"C3CB",
			x"0000" when x"C3CC",
			x"0000" when x"C3CD",
			x"0000" when x"C3CE",
			x"0000" when x"C3CF",
			x"0000" when x"C3D0",
			x"0000" when x"C3D1",
			x"0000" when x"C3D2",
			x"0000" when x"C3D3",
			x"0000" when x"C3D4",
			x"0000" when x"C3D5",
			x"0000" when x"C3D6",
			x"0000" when x"C3D7",
			x"0000" when x"C3D8",
			x"0000" when x"C3D9",
			x"0000" when x"C3DA",
			x"0000" when x"C3DB",
			x"0000" when x"C3DC",
			x"0000" when x"C3DD",
			x"0000" when x"C3DE",
			x"0000" when x"C3DF",
			x"0000" when x"C3E0",
			x"0000" when x"C3E1",
			x"0000" when x"C3E2",
			x"0000" when x"C3E3",
			x"0000" when x"C3E4",
			x"0000" when x"C3E5",
			x"0000" when x"C3E6",
			x"0000" when x"C3E7",
			x"0000" when x"C3E8",
			x"0000" when x"C3E9",
			x"0000" when x"C3EA",
			x"0000" when x"C3EB",
			x"0000" when x"C3EC",
			x"0000" when x"C3ED",
			x"0000" when x"C3EE",
			x"0000" when x"C3EF",
			x"0000" when x"C3F0",
			x"0000" when x"C3F1",
			x"0000" when x"C3F2",
			x"0000" when x"C3F3",
			x"0000" when x"C3F4",
			x"0000" when x"C3F5",
			x"0000" when x"C3F6",
			x"0000" when x"C3F7",
			x"0000" when x"C3F8",
			x"0000" when x"C3F9",
			x"0000" when x"C3FA",
			x"0000" when x"C3FB",
			x"0000" when x"C3FC",
			x"0000" when x"C3FD",
			x"0000" when x"C3FE",
			x"0000" when x"C3FF",
			x"0000" when x"C400",
			x"0000" when x"C401",
			x"0000" when x"C402",
			x"0000" when x"C403",
			x"0000" when x"C404",
			x"0000" when x"C405",
			x"0000" when x"C406",
			x"0000" when x"C407",
			x"0000" when x"C408",
			x"0000" when x"C409",
			x"0000" when x"C40A",
			x"0000" when x"C40B",
			x"0000" when x"C40C",
			x"0000" when x"C40D",
			x"0000" when x"C40E",
			x"0000" when x"C40F",
			x"0000" when x"C410",
			x"0000" when x"C411",
			x"0000" when x"C412",
			x"0000" when x"C413",
			x"0000" when x"C414",
			x"0000" when x"C415",
			x"0000" when x"C416",
			x"0000" when x"C417",
			x"0000" when x"C418",
			x"0000" when x"C419",
			x"0000" when x"C41A",
			x"0000" when x"C41B",
			x"0000" when x"C41C",
			x"0000" when x"C41D",
			x"0000" when x"C41E",
			x"0000" when x"C41F",
			x"0000" when x"C420",
			x"0000" when x"C421",
			x"0000" when x"C422",
			x"0000" when x"C423",
			x"0000" when x"C424",
			x"0000" when x"C425",
			x"0000" when x"C426",
			x"0000" when x"C427",
			x"0000" when x"C428",
			x"0000" when x"C429",
			x"0000" when x"C42A",
			x"0000" when x"C42B",
			x"0000" when x"C42C",
			x"0000" when x"C42D",
			x"0000" when x"C42E",
			x"0000" when x"C42F",
			x"0000" when x"C430",
			x"0000" when x"C431",
			x"0000" when x"C432",
			x"0000" when x"C433",
			x"0000" when x"C434",
			x"0000" when x"C435",
			x"0000" when x"C436",
			x"0000" when x"C437",
			x"0000" when x"C438",
			x"0000" when x"C439",
			x"0000" when x"C43A",
			x"0000" when x"C43B",
			x"0000" when x"C43C",
			x"0000" when x"C43D",
			x"0000" when x"C43E",
			x"0000" when x"C43F",
			x"0000" when x"C440",
			x"0000" when x"C441",
			x"0000" when x"C442",
			x"0000" when x"C443",
			x"0000" when x"C444",
			x"0000" when x"C445",
			x"0000" when x"C446",
			x"0000" when x"C447",
			x"0000" when x"C448",
			x"0000" when x"C449",
			x"0000" when x"C44A",
			x"0000" when x"C44B",
			x"0000" when x"C44C",
			x"0000" when x"C44D",
			x"0000" when x"C44E",
			x"0000" when x"C44F",
			x"0000" when x"C450",
			x"0000" when x"C451",
			x"0000" when x"C452",
			x"0000" when x"C453",
			x"0000" when x"C454",
			x"0000" when x"C455",
			x"0000" when x"C456",
			x"0000" when x"C457",
			x"0000" when x"C458",
			x"0000" when x"C459",
			x"0000" when x"C45A",
			x"0000" when x"C45B",
			x"0000" when x"C45C",
			x"0000" when x"C45D",
			x"0000" when x"C45E",
			x"0000" when x"C45F",
			x"0000" when x"C460",
			x"0000" when x"C461",
			x"0000" when x"C462",
			x"0000" when x"C463",
			x"0000" when x"C464",
			x"0000" when x"C465",
			x"0000" when x"C466",
			x"0000" when x"C467",
			x"0000" when x"C468",
			x"0000" when x"C469",
			x"0000" when x"C46A",
			x"0000" when x"C46B",
			x"0000" when x"C46C",
			x"0000" when x"C46D",
			x"0000" when x"C46E",
			x"0000" when x"C46F",
			x"0000" when x"C470",
			x"0000" when x"C471",
			x"0000" when x"C472",
			x"0000" when x"C473",
			x"0000" when x"C474",
			x"0000" when x"C475",
			x"0000" when x"C476",
			x"0000" when x"C477",
			x"0000" when x"C478",
			x"0000" when x"C479",
			x"0000" when x"C47A",
			x"0000" when x"C47B",
			x"0000" when x"C47C",
			x"0000" when x"C47D",
			x"0000" when x"C47E",
			x"0000" when x"C47F",
			x"0000" when x"C480",
			x"0000" when x"C481",
			x"0000" when x"C482",
			x"0000" when x"C483",
			x"0000" when x"C484",
			x"0000" when x"C485",
			x"0000" when x"C486",
			x"0000" when x"C487",
			x"0000" when x"C488",
			x"0000" when x"C489",
			x"0000" when x"C48A",
			x"0000" when x"C48B",
			x"0000" when x"C48C",
			x"0000" when x"C48D",
			x"0000" when x"C48E",
			x"0000" when x"C48F",
			x"0000" when x"C490",
			x"0000" when x"C491",
			x"0000" when x"C492",
			x"0000" when x"C493",
			x"0000" when x"C494",
			x"0000" when x"C495",
			x"0000" when x"C496",
			x"0000" when x"C497",
			x"0000" when x"C498",
			x"0000" when x"C499",
			x"0000" when x"C49A",
			x"0000" when x"C49B",
			x"0000" when x"C49C",
			x"0000" when x"C49D",
			x"0000" when x"C49E",
			x"0000" when x"C49F",
			x"0000" when x"C4A0",
			x"0000" when x"C4A1",
			x"0000" when x"C4A2",
			x"0000" when x"C4A3",
			x"0000" when x"C4A4",
			x"0000" when x"C4A5",
			x"0000" when x"C4A6",
			x"0000" when x"C4A7",
			x"0000" when x"C4A8",
			x"0000" when x"C4A9",
			x"0000" when x"C4AA",
			x"0000" when x"C4AB",
			x"0000" when x"C4AC",
			x"0000" when x"C4AD",
			x"0000" when x"C4AE",
			x"0000" when x"C4AF",
			x"0000" when x"C4B0",
			x"0000" when x"C4B1",
			x"0000" when x"C4B2",
			x"0000" when x"C4B3",
			x"0000" when x"C4B4",
			x"0000" when x"C4B5",
			x"0000" when x"C4B6",
			x"0000" when x"C4B7",
			x"0000" when x"C4B8",
			x"0000" when x"C4B9",
			x"0000" when x"C4BA",
			x"0000" when x"C4BB",
			x"0000" when x"C4BC",
			x"0000" when x"C4BD",
			x"0000" when x"C4BE",
			x"0000" when x"C4BF",
			x"0000" when x"C4C0",
			x"0000" when x"C4C1",
			x"0000" when x"C4C2",
			x"0000" when x"C4C3",
			x"0000" when x"C4C4",
			x"0000" when x"C4C5",
			x"0000" when x"C4C6",
			x"0000" when x"C4C7",
			x"0000" when x"C4C8",
			x"0000" when x"C4C9",
			x"0000" when x"C4CA",
			x"0000" when x"C4CB",
			x"0000" when x"C4CC",
			x"0000" when x"C4CD",
			x"0000" when x"C4CE",
			x"0000" when x"C4CF",
			x"0000" when x"C4D0",
			x"0000" when x"C4D1",
			x"0000" when x"C4D2",
			x"0000" when x"C4D3",
			x"0000" when x"C4D4",
			x"0000" when x"C4D5",
			x"0000" when x"C4D6",
			x"0000" when x"C4D7",
			x"0000" when x"C4D8",
			x"0000" when x"C4D9",
			x"0000" when x"C4DA",
			x"0000" when x"C4DB",
			x"0000" when x"C4DC",
			x"0000" when x"C4DD",
			x"0000" when x"C4DE",
			x"0000" when x"C4DF",
			x"0000" when x"C4E0",
			x"0000" when x"C4E1",
			x"0000" when x"C4E2",
			x"0000" when x"C4E3",
			x"0000" when x"C4E4",
			x"0000" when x"C4E5",
			x"0000" when x"C4E6",
			x"0000" when x"C4E7",
			x"0000" when x"C4E8",
			x"0000" when x"C4E9",
			x"0000" when x"C4EA",
			x"0000" when x"C4EB",
			x"0000" when x"C4EC",
			x"0000" when x"C4ED",
			x"0000" when x"C4EE",
			x"0000" when x"C4EF",
			x"0000" when x"C4F0",
			x"0000" when x"C4F1",
			x"0000" when x"C4F2",
			x"0000" when x"C4F3",
			x"0000" when x"C4F4",
			x"0000" when x"C4F5",
			x"0000" when x"C4F6",
			x"0000" when x"C4F7",
			x"0000" when x"C4F8",
			x"0000" when x"C4F9",
			x"0000" when x"C4FA",
			x"0000" when x"C4FB",
			x"0000" when x"C4FC",
			x"0000" when x"C4FD",
			x"0000" when x"C4FE",
			x"0000" when x"C4FF",
			x"0000" when x"C500",
			x"0000" when x"C501",
			x"0000" when x"C502",
			x"0000" when x"C503",
			x"0000" when x"C504",
			x"0000" when x"C505",
			x"0000" when x"C506",
			x"0000" when x"C507",
			x"0000" when x"C508",
			x"0000" when x"C509",
			x"0000" when x"C50A",
			x"0000" when x"C50B",
			x"0000" when x"C50C",
			x"0000" when x"C50D",
			x"0000" when x"C50E",
			x"0000" when x"C50F",
			x"0000" when x"C510",
			x"0000" when x"C511",
			x"0000" when x"C512",
			x"0000" when x"C513",
			x"0000" when x"C514",
			x"0000" when x"C515",
			x"0000" when x"C516",
			x"0000" when x"C517",
			x"0000" when x"C518",
			x"0000" when x"C519",
			x"0000" when x"C51A",
			x"0000" when x"C51B",
			x"0000" when x"C51C",
			x"0000" when x"C51D",
			x"0000" when x"C51E",
			x"0000" when x"C51F",
			x"0000" when x"C520",
			x"0000" when x"C521",
			x"0000" when x"C522",
			x"0000" when x"C523",
			x"0000" when x"C524",
			x"0000" when x"C525",
			x"0000" when x"C526",
			x"0000" when x"C527",
			x"0000" when x"C528",
			x"0000" when x"C529",
			x"0000" when x"C52A",
			x"0000" when x"C52B",
			x"0000" when x"C52C",
			x"0000" when x"C52D",
			x"0000" when x"C52E",
			x"0000" when x"C52F",
			x"0000" when x"C530",
			x"0000" when x"C531",
			x"0000" when x"C532",
			x"0000" when x"C533",
			x"0000" when x"C534",
			x"0000" when x"C535",
			x"0000" when x"C536",
			x"0000" when x"C537",
			x"0000" when x"C538",
			x"0000" when x"C539",
			x"0000" when x"C53A",
			x"0000" when x"C53B",
			x"0000" when x"C53C",
			x"0000" when x"C53D",
			x"0000" when x"C53E",
			x"0000" when x"C53F",
			x"0000" when x"C540",
			x"0000" when x"C541",
			x"0000" when x"C542",
			x"0000" when x"C543",
			x"0000" when x"C544",
			x"0000" when x"C545",
			x"0000" when x"C546",
			x"0000" when x"C547",
			x"0000" when x"C548",
			x"0000" when x"C549",
			x"0000" when x"C54A",
			x"0000" when x"C54B",
			x"0000" when x"C54C",
			x"0000" when x"C54D",
			x"0000" when x"C54E",
			x"0000" when x"C54F",
			x"0000" when x"C550",
			x"0000" when x"C551",
			x"0000" when x"C552",
			x"0000" when x"C553",
			x"0000" when x"C554",
			x"0000" when x"C555",
			x"0000" when x"C556",
			x"0000" when x"C557",
			x"0000" when x"C558",
			x"0000" when x"C559",
			x"0000" when x"C55A",
			x"0000" when x"C55B",
			x"0000" when x"C55C",
			x"0000" when x"C55D",
			x"0000" when x"C55E",
			x"0000" when x"C55F",
			x"0000" when x"C560",
			x"0000" when x"C561",
			x"0000" when x"C562",
			x"0000" when x"C563",
			x"0000" when x"C564",
			x"0000" when x"C565",
			x"0000" when x"C566",
			x"0000" when x"C567",
			x"0000" when x"C568",
			x"0000" when x"C569",
			x"0000" when x"C56A",
			x"0000" when x"C56B",
			x"0000" when x"C56C",
			x"0000" when x"C56D",
			x"0000" when x"C56E",
			x"0000" when x"C56F",
			x"0000" when x"C570",
			x"0000" when x"C571",
			x"0000" when x"C572",
			x"0000" when x"C573",
			x"0000" when x"C574",
			x"0000" when x"C575",
			x"0000" when x"C576",
			x"0000" when x"C577",
			x"0000" when x"C578",
			x"0000" when x"C579",
			x"0000" when x"C57A",
			x"0000" when x"C57B",
			x"0000" when x"C57C",
			x"0000" when x"C57D",
			x"0000" when x"C57E",
			x"0000" when x"C57F",
			x"0000" when x"C580",
			x"0000" when x"C581",
			x"0000" when x"C582",
			x"0000" when x"C583",
			x"0000" when x"C584",
			x"0000" when x"C585",
			x"0000" when x"C586",
			x"0000" when x"C587",
			x"0000" when x"C588",
			x"0000" when x"C589",
			x"0000" when x"C58A",
			x"0000" when x"C58B",
			x"0000" when x"C58C",
			x"0000" when x"C58D",
			x"0000" when x"C58E",
			x"0000" when x"C58F",
			x"0000" when x"C590",
			x"0000" when x"C591",
			x"0000" when x"C592",
			x"0000" when x"C593",
			x"0000" when x"C594",
			x"0000" when x"C595",
			x"0000" when x"C596",
			x"0000" when x"C597",
			x"0000" when x"C598",
			x"0000" when x"C599",
			x"0000" when x"C59A",
			x"0000" when x"C59B",
			x"0000" when x"C59C",
			x"0000" when x"C59D",
			x"0000" when x"C59E",
			x"0000" when x"C59F",
			x"0000" when x"C5A0",
			x"0000" when x"C5A1",
			x"0000" when x"C5A2",
			x"0000" when x"C5A3",
			x"0000" when x"C5A4",
			x"0000" when x"C5A5",
			x"0000" when x"C5A6",
			x"0000" when x"C5A7",
			x"0000" when x"C5A8",
			x"0000" when x"C5A9",
			x"0000" when x"C5AA",
			x"0000" when x"C5AB",
			x"0000" when x"C5AC",
			x"0000" when x"C5AD",
			x"0000" when x"C5AE",
			x"0000" when x"C5AF",
			x"0000" when x"C5B0",
			x"0000" when x"C5B1",
			x"0000" when x"C5B2",
			x"0000" when x"C5B3",
			x"0000" when x"C5B4",
			x"0000" when x"C5B5",
			x"0000" when x"C5B6",
			x"0000" when x"C5B7",
			x"0000" when x"C5B8",
			x"0000" when x"C5B9",
			x"0000" when x"C5BA",
			x"0000" when x"C5BB",
			x"0000" when x"C5BC",
			x"0000" when x"C5BD",
			x"0000" when x"C5BE",
			x"0000" when x"C5BF",
			x"0000" when x"C5C0",
			x"0000" when x"C5C1",
			x"0000" when x"C5C2",
			x"0000" when x"C5C3",
			x"0000" when x"C5C4",
			x"0000" when x"C5C5",
			x"0000" when x"C5C6",
			x"0000" when x"C5C7",
			x"0000" when x"C5C8",
			x"0000" when x"C5C9",
			x"0000" when x"C5CA",
			x"0000" when x"C5CB",
			x"0000" when x"C5CC",
			x"0000" when x"C5CD",
			x"0000" when x"C5CE",
			x"0000" when x"C5CF",
			x"0000" when x"C5D0",
			x"0000" when x"C5D1",
			x"0000" when x"C5D2",
			x"0000" when x"C5D3",
			x"0000" when x"C5D4",
			x"0000" when x"C5D5",
			x"0000" when x"C5D6",
			x"0000" when x"C5D7",
			x"0000" when x"C5D8",
			x"0000" when x"C5D9",
			x"0000" when x"C5DA",
			x"0000" when x"C5DB",
			x"0000" when x"C5DC",
			x"0000" when x"C5DD",
			x"0000" when x"C5DE",
			x"0000" when x"C5DF",
			x"0000" when x"C5E0",
			x"0000" when x"C5E1",
			x"0000" when x"C5E2",
			x"0000" when x"C5E3",
			x"0000" when x"C5E4",
			x"0000" when x"C5E5",
			x"0000" when x"C5E6",
			x"0000" when x"C5E7",
			x"0000" when x"C5E8",
			x"0000" when x"C5E9",
			x"0000" when x"C5EA",
			x"0000" when x"C5EB",
			x"0000" when x"C5EC",
			x"0000" when x"C5ED",
			x"0000" when x"C5EE",
			x"0000" when x"C5EF",
			x"0000" when x"C5F0",
			x"0000" when x"C5F1",
			x"0000" when x"C5F2",
			x"0000" when x"C5F3",
			x"0000" when x"C5F4",
			x"0000" when x"C5F5",
			x"0000" when x"C5F6",
			x"0000" when x"C5F7",
			x"0000" when x"C5F8",
			x"0000" when x"C5F9",
			x"0000" when x"C5FA",
			x"0000" when x"C5FB",
			x"0000" when x"C5FC",
			x"0000" when x"C5FD",
			x"0000" when x"C5FE",
			x"0000" when x"C5FF",
			x"0000" when x"C600",
			x"0000" when x"C601",
			x"0000" when x"C602",
			x"0000" when x"C603",
			x"0000" when x"C604",
			x"0000" when x"C605",
			x"0000" when x"C606",
			x"0000" when x"C607",
			x"0000" when x"C608",
			x"0000" when x"C609",
			x"0000" when x"C60A",
			x"0000" when x"C60B",
			x"0000" when x"C60C",
			x"0000" when x"C60D",
			x"0000" when x"C60E",
			x"0000" when x"C60F",
			x"0000" when x"C610",
			x"0000" when x"C611",
			x"0000" when x"C612",
			x"0000" when x"C613",
			x"0000" when x"C614",
			x"0000" when x"C615",
			x"0000" when x"C616",
			x"0000" when x"C617",
			x"0000" when x"C618",
			x"0000" when x"C619",
			x"0000" when x"C61A",
			x"0000" when x"C61B",
			x"0000" when x"C61C",
			x"0000" when x"C61D",
			x"0000" when x"C61E",
			x"0000" when x"C61F",
			x"0000" when x"C620",
			x"0000" when x"C621",
			x"0000" when x"C622",
			x"0000" when x"C623",
			x"0000" when x"C624",
			x"0000" when x"C625",
			x"0000" when x"C626",
			x"0000" when x"C627",
			x"0000" when x"C628",
			x"0000" when x"C629",
			x"0000" when x"C62A",
			x"0000" when x"C62B",
			x"0000" when x"C62C",
			x"0000" when x"C62D",
			x"0000" when x"C62E",
			x"0000" when x"C62F",
			x"0000" when x"C630",
			x"0000" when x"C631",
			x"0000" when x"C632",
			x"0000" when x"C633",
			x"0000" when x"C634",
			x"0000" when x"C635",
			x"0000" when x"C636",
			x"0000" when x"C637",
			x"0000" when x"C638",
			x"0000" when x"C639",
			x"0000" when x"C63A",
			x"0000" when x"C63B",
			x"0000" when x"C63C",
			x"0000" when x"C63D",
			x"0000" when x"C63E",
			x"0000" when x"C63F",
			x"0000" when x"C640",
			x"0000" when x"C641",
			x"0000" when x"C642",
			x"0000" when x"C643",
			x"0000" when x"C644",
			x"0000" when x"C645",
			x"0000" when x"C646",
			x"0000" when x"C647",
			x"0000" when x"C648",
			x"0000" when x"C649",
			x"0000" when x"C64A",
			x"0000" when x"C64B",
			x"0000" when x"C64C",
			x"0000" when x"C64D",
			x"0000" when x"C64E",
			x"0000" when x"C64F",
			x"0000" when x"C650",
			x"0000" when x"C651",
			x"0000" when x"C652",
			x"0000" when x"C653",
			x"0000" when x"C654",
			x"0000" when x"C655",
			x"0000" when x"C656",
			x"0000" when x"C657",
			x"0000" when x"C658",
			x"0000" when x"C659",
			x"0000" when x"C65A",
			x"0000" when x"C65B",
			x"0000" when x"C65C",
			x"0000" when x"C65D",
			x"0000" when x"C65E",
			x"0000" when x"C65F",
			x"0000" when x"C660",
			x"0000" when x"C661",
			x"0000" when x"C662",
			x"0000" when x"C663",
			x"0000" when x"C664",
			x"0000" when x"C665",
			x"0000" when x"C666",
			x"0000" when x"C667",
			x"0000" when x"C668",
			x"0000" when x"C669",
			x"0000" when x"C66A",
			x"0000" when x"C66B",
			x"0000" when x"C66C",
			x"0000" when x"C66D",
			x"0000" when x"C66E",
			x"0000" when x"C66F",
			x"0000" when x"C670",
			x"0000" when x"C671",
			x"0000" when x"C672",
			x"0000" when x"C673",
			x"0000" when x"C674",
			x"0000" when x"C675",
			x"0000" when x"C676",
			x"0000" when x"C677",
			x"0000" when x"C678",
			x"0000" when x"C679",
			x"0000" when x"C67A",
			x"0000" when x"C67B",
			x"0000" when x"C67C",
			x"0000" when x"C67D",
			x"0000" when x"C67E",
			x"0000" when x"C67F",
			x"0000" when x"C680",
			x"0000" when x"C681",
			x"0000" when x"C682",
			x"0000" when x"C683",
			x"0000" when x"C684",
			x"0000" when x"C685",
			x"0000" when x"C686",
			x"0000" when x"C687",
			x"0000" when x"C688",
			x"0000" when x"C689",
			x"0000" when x"C68A",
			x"0000" when x"C68B",
			x"0000" when x"C68C",
			x"0000" when x"C68D",
			x"0000" when x"C68E",
			x"0000" when x"C68F",
			x"0000" when x"C690",
			x"0000" when x"C691",
			x"0000" when x"C692",
			x"0000" when x"C693",
			x"0000" when x"C694",
			x"0000" when x"C695",
			x"0000" when x"C696",
			x"0000" when x"C697",
			x"0000" when x"C698",
			x"0000" when x"C699",
			x"0000" when x"C69A",
			x"0000" when x"C69B",
			x"0000" when x"C69C",
			x"0000" when x"C69D",
			x"0000" when x"C69E",
			x"0000" when x"C69F",
			x"0000" when x"C6A0",
			x"0000" when x"C6A1",
			x"0000" when x"C6A2",
			x"0000" when x"C6A3",
			x"0000" when x"C6A4",
			x"0000" when x"C6A5",
			x"0000" when x"C6A6",
			x"0000" when x"C6A7",
			x"0000" when x"C6A8",
			x"0000" when x"C6A9",
			x"0000" when x"C6AA",
			x"0000" when x"C6AB",
			x"0000" when x"C6AC",
			x"0000" when x"C6AD",
			x"0000" when x"C6AE",
			x"0000" when x"C6AF",
			x"0000" when x"C6B0",
			x"0000" when x"C6B1",
			x"0000" when x"C6B2",
			x"0000" when x"C6B3",
			x"0000" when x"C6B4",
			x"0000" when x"C6B5",
			x"0000" when x"C6B6",
			x"0000" when x"C6B7",
			x"0000" when x"C6B8",
			x"0000" when x"C6B9",
			x"0000" when x"C6BA",
			x"0000" when x"C6BB",
			x"0000" when x"C6BC",
			x"0000" when x"C6BD",
			x"0000" when x"C6BE",
			x"0000" when x"C6BF",
			x"0000" when x"C6C0",
			x"0000" when x"C6C1",
			x"0000" when x"C6C2",
			x"0000" when x"C6C3",
			x"0000" when x"C6C4",
			x"0000" when x"C6C5",
			x"0000" when x"C6C6",
			x"0000" when x"C6C7",
			x"0000" when x"C6C8",
			x"0000" when x"C6C9",
			x"0000" when x"C6CA",
			x"0000" when x"C6CB",
			x"0000" when x"C6CC",
			x"0000" when x"C6CD",
			x"0000" when x"C6CE",
			x"0000" when x"C6CF",
			x"0000" when x"C6D0",
			x"0000" when x"C6D1",
			x"0000" when x"C6D2",
			x"0000" when x"C6D3",
			x"0000" when x"C6D4",
			x"0000" when x"C6D5",
			x"0000" when x"C6D6",
			x"0000" when x"C6D7",
			x"0000" when x"C6D8",
			x"0000" when x"C6D9",
			x"0000" when x"C6DA",
			x"0000" when x"C6DB",
			x"0000" when x"C6DC",
			x"0000" when x"C6DD",
			x"0000" when x"C6DE",
			x"0000" when x"C6DF",
			x"0000" when x"C6E0",
			x"0000" when x"C6E1",
			x"0000" when x"C6E2",
			x"0000" when x"C6E3",
			x"0000" when x"C6E4",
			x"0000" when x"C6E5",
			x"0000" when x"C6E6",
			x"0000" when x"C6E7",
			x"0000" when x"C6E8",
			x"0000" when x"C6E9",
			x"0000" when x"C6EA",
			x"0000" when x"C6EB",
			x"0000" when x"C6EC",
			x"0000" when x"C6ED",
			x"0000" when x"C6EE",
			x"0000" when x"C6EF",
			x"0000" when x"C6F0",
			x"0000" when x"C6F1",
			x"0000" when x"C6F2",
			x"0000" when x"C6F3",
			x"0000" when x"C6F4",
			x"0000" when x"C6F5",
			x"0000" when x"C6F6",
			x"0000" when x"C6F7",
			x"0000" when x"C6F8",
			x"0000" when x"C6F9",
			x"0000" when x"C6FA",
			x"0000" when x"C6FB",
			x"0000" when x"C6FC",
			x"0000" when x"C6FD",
			x"0000" when x"C6FE",
			x"0000" when x"C6FF",
			x"0000" when x"C700",
			x"0000" when x"C701",
			x"0000" when x"C702",
			x"0000" when x"C703",
			x"0000" when x"C704",
			x"0000" when x"C705",
			x"0000" when x"C706",
			x"0000" when x"C707",
			x"0000" when x"C708",
			x"0000" when x"C709",
			x"0000" when x"C70A",
			x"0000" when x"C70B",
			x"0000" when x"C70C",
			x"0000" when x"C70D",
			x"0000" when x"C70E",
			x"0000" when x"C70F",
			x"0000" when x"C710",
			x"0000" when x"C711",
			x"0000" when x"C712",
			x"0000" when x"C713",
			x"0000" when x"C714",
			x"0000" when x"C715",
			x"0000" when x"C716",
			x"0000" when x"C717",
			x"0000" when x"C718",
			x"0000" when x"C719",
			x"0000" when x"C71A",
			x"0000" when x"C71B",
			x"0000" when x"C71C",
			x"0000" when x"C71D",
			x"0000" when x"C71E",
			x"0000" when x"C71F",
			x"0000" when x"C720",
			x"0000" when x"C721",
			x"0000" when x"C722",
			x"0000" when x"C723",
			x"0000" when x"C724",
			x"0000" when x"C725",
			x"0000" when x"C726",
			x"0000" when x"C727",
			x"0000" when x"C728",
			x"0000" when x"C729",
			x"0000" when x"C72A",
			x"0000" when x"C72B",
			x"0000" when x"C72C",
			x"0000" when x"C72D",
			x"0000" when x"C72E",
			x"0000" when x"C72F",
			x"0000" when x"C730",
			x"0000" when x"C731",
			x"0000" when x"C732",
			x"0000" when x"C733",
			x"0000" when x"C734",
			x"0000" when x"C735",
			x"0000" when x"C736",
			x"0000" when x"C737",
			x"0000" when x"C738",
			x"0000" when x"C739",
			x"0000" when x"C73A",
			x"0000" when x"C73B",
			x"0000" when x"C73C",
			x"0000" when x"C73D",
			x"0000" when x"C73E",
			x"0000" when x"C73F",
			x"0000" when x"C740",
			x"0000" when x"C741",
			x"0000" when x"C742",
			x"0000" when x"C743",
			x"0000" when x"C744",
			x"0000" when x"C745",
			x"0000" when x"C746",
			x"0000" when x"C747",
			x"0000" when x"C748",
			x"0000" when x"C749",
			x"0000" when x"C74A",
			x"0000" when x"C74B",
			x"0000" when x"C74C",
			x"0000" when x"C74D",
			x"0000" when x"C74E",
			x"0000" when x"C74F",
			x"0000" when x"C750",
			x"0000" when x"C751",
			x"0000" when x"C752",
			x"0000" when x"C753",
			x"0000" when x"C754",
			x"0000" when x"C755",
			x"0000" when x"C756",
			x"0000" when x"C757",
			x"0000" when x"C758",
			x"0000" when x"C759",
			x"0000" when x"C75A",
			x"0000" when x"C75B",
			x"0000" when x"C75C",
			x"0000" when x"C75D",
			x"0000" when x"C75E",
			x"0000" when x"C75F",
			x"0000" when x"C760",
			x"0000" when x"C761",
			x"0000" when x"C762",
			x"0000" when x"C763",
			x"0000" when x"C764",
			x"0000" when x"C765",
			x"0000" when x"C766",
			x"0000" when x"C767",
			x"0000" when x"C768",
			x"0000" when x"C769",
			x"0000" when x"C76A",
			x"0000" when x"C76B",
			x"0000" when x"C76C",
			x"0000" when x"C76D",
			x"0000" when x"C76E",
			x"0000" when x"C76F",
			x"0000" when x"C770",
			x"0000" when x"C771",
			x"0000" when x"C772",
			x"0000" when x"C773",
			x"0000" when x"C774",
			x"0000" when x"C775",
			x"0000" when x"C776",
			x"0000" when x"C777",
			x"0000" when x"C778",
			x"0000" when x"C779",
			x"0000" when x"C77A",
			x"0000" when x"C77B",
			x"0000" when x"C77C",
			x"0000" when x"C77D",
			x"0000" when x"C77E",
			x"0000" when x"C77F",
			x"0000" when x"C780",
			x"0000" when x"C781",
			x"0000" when x"C782",
			x"0000" when x"C783",
			x"0000" when x"C784",
			x"0000" when x"C785",
			x"0000" when x"C786",
			x"0000" when x"C787",
			x"0000" when x"C788",
			x"0000" when x"C789",
			x"0000" when x"C78A",
			x"0000" when x"C78B",
			x"0000" when x"C78C",
			x"0000" when x"C78D",
			x"0000" when x"C78E",
			x"0000" when x"C78F",
			x"0000" when x"C790",
			x"0000" when x"C791",
			x"0000" when x"C792",
			x"0000" when x"C793",
			x"0000" when x"C794",
			x"0000" when x"C795",
			x"0000" when x"C796",
			x"0000" when x"C797",
			x"0000" when x"C798",
			x"0000" when x"C799",
			x"0000" when x"C79A",
			x"0000" when x"C79B",
			x"0000" when x"C79C",
			x"0000" when x"C79D",
			x"0000" when x"C79E",
			x"0000" when x"C79F",
			x"0000" when x"C7A0",
			x"0000" when x"C7A1",
			x"0000" when x"C7A2",
			x"0000" when x"C7A3",
			x"0000" when x"C7A4",
			x"0000" when x"C7A5",
			x"0000" when x"C7A6",
			x"0000" when x"C7A7",
			x"0000" when x"C7A8",
			x"0000" when x"C7A9",
			x"0000" when x"C7AA",
			x"0000" when x"C7AB",
			x"0000" when x"C7AC",
			x"0000" when x"C7AD",
			x"0000" when x"C7AE",
			x"0000" when x"C7AF",
			x"0000" when x"C7B0",
			x"0000" when x"C7B1",
			x"0000" when x"C7B2",
			x"0000" when x"C7B3",
			x"0000" when x"C7B4",
			x"0000" when x"C7B5",
			x"0000" when x"C7B6",
			x"0000" when x"C7B7",
			x"0000" when x"C7B8",
			x"0000" when x"C7B9",
			x"0000" when x"C7BA",
			x"0000" when x"C7BB",
			x"0000" when x"C7BC",
			x"0000" when x"C7BD",
			x"0000" when x"C7BE",
			x"0000" when x"C7BF",
			x"0000" when x"C7C0",
			x"0000" when x"C7C1",
			x"0000" when x"C7C2",
			x"0000" when x"C7C3",
			x"0000" when x"C7C4",
			x"0000" when x"C7C5",
			x"0000" when x"C7C6",
			x"0000" when x"C7C7",
			x"0000" when x"C7C8",
			x"0000" when x"C7C9",
			x"0000" when x"C7CA",
			x"0000" when x"C7CB",
			x"0000" when x"C7CC",
			x"0000" when x"C7CD",
			x"0000" when x"C7CE",
			x"0000" when x"C7CF",
			x"0000" when x"C7D0",
			x"0000" when x"C7D1",
			x"0000" when x"C7D2",
			x"0000" when x"C7D3",
			x"0000" when x"C7D4",
			x"0000" when x"C7D5",
			x"0000" when x"C7D6",
			x"0000" when x"C7D7",
			x"0000" when x"C7D8",
			x"0000" when x"C7D9",
			x"0000" when x"C7DA",
			x"0000" when x"C7DB",
			x"0000" when x"C7DC",
			x"0000" when x"C7DD",
			x"0000" when x"C7DE",
			x"0000" when x"C7DF",
			x"0000" when x"C7E0",
			x"0000" when x"C7E1",
			x"0000" when x"C7E2",
			x"0000" when x"C7E3",
			x"0000" when x"C7E4",
			x"0000" when x"C7E5",
			x"0000" when x"C7E6",
			x"0000" when x"C7E7",
			x"0000" when x"C7E8",
			x"0000" when x"C7E9",
			x"0000" when x"C7EA",
			x"0000" when x"C7EB",
			x"0000" when x"C7EC",
			x"0000" when x"C7ED",
			x"0000" when x"C7EE",
			x"0000" when x"C7EF",
			x"0000" when x"C7F0",
			x"0000" when x"C7F1",
			x"0000" when x"C7F2",
			x"0000" when x"C7F3",
			x"0000" when x"C7F4",
			x"0000" when x"C7F5",
			x"0000" when x"C7F6",
			x"0000" when x"C7F7",
			x"0000" when x"C7F8",
			x"0000" when x"C7F9",
			x"0000" when x"C7FA",
			x"0000" when x"C7FB",
			x"0000" when x"C7FC",
			x"0000" when x"C7FD",
			x"0000" when x"C7FE",
			x"0000" when x"C7FF",
			x"0000" when x"C800",
			x"0000" when x"C801",
			x"0000" when x"C802",
			x"0000" when x"C803",
			x"0000" when x"C804",
			x"0000" when x"C805",
			x"0000" when x"C806",
			x"0000" when x"C807",
			x"0000" when x"C808",
			x"0000" when x"C809",
			x"0000" when x"C80A",
			x"0000" when x"C80B",
			x"0000" when x"C80C",
			x"0000" when x"C80D",
			x"0000" when x"C80E",
			x"0000" when x"C80F",
			x"0000" when x"C810",
			x"0000" when x"C811",
			x"0000" when x"C812",
			x"0000" when x"C813",
			x"0000" when x"C814",
			x"0000" when x"C815",
			x"0000" when x"C816",
			x"0000" when x"C817",
			x"0000" when x"C818",
			x"0000" when x"C819",
			x"0000" when x"C81A",
			x"0000" when x"C81B",
			x"0000" when x"C81C",
			x"0000" when x"C81D",
			x"0000" when x"C81E",
			x"0000" when x"C81F",
			x"0000" when x"C820",
			x"0000" when x"C821",
			x"0000" when x"C822",
			x"0000" when x"C823",
			x"0000" when x"C824",
			x"0000" when x"C825",
			x"0000" when x"C826",
			x"0000" when x"C827",
			x"0000" when x"C828",
			x"0000" when x"C829",
			x"0000" when x"C82A",
			x"0000" when x"C82B",
			x"0000" when x"C82C",
			x"0000" when x"C82D",
			x"0000" when x"C82E",
			x"0000" when x"C82F",
			x"0000" when x"C830",
			x"0000" when x"C831",
			x"0000" when x"C832",
			x"0000" when x"C833",
			x"0000" when x"C834",
			x"0000" when x"C835",
			x"0000" when x"C836",
			x"0000" when x"C837",
			x"0000" when x"C838",
			x"0000" when x"C839",
			x"0000" when x"C83A",
			x"0000" when x"C83B",
			x"0000" when x"C83C",
			x"0000" when x"C83D",
			x"0000" when x"C83E",
			x"0000" when x"C83F",
			x"0000" when x"C840",
			x"0000" when x"C841",
			x"0000" when x"C842",
			x"0000" when x"C843",
			x"0000" when x"C844",
			x"0000" when x"C845",
			x"0000" when x"C846",
			x"0000" when x"C847",
			x"0000" when x"C848",
			x"0000" when x"C849",
			x"0000" when x"C84A",
			x"0000" when x"C84B",
			x"0000" when x"C84C",
			x"0000" when x"C84D",
			x"0000" when x"C84E",
			x"0000" when x"C84F",
			x"0000" when x"C850",
			x"0000" when x"C851",
			x"0000" when x"C852",
			x"0000" when x"C853",
			x"0000" when x"C854",
			x"0000" when x"C855",
			x"0000" when x"C856",
			x"0000" when x"C857",
			x"0000" when x"C858",
			x"0000" when x"C859",
			x"0000" when x"C85A",
			x"0000" when x"C85B",
			x"0000" when x"C85C",
			x"0000" when x"C85D",
			x"0000" when x"C85E",
			x"0000" when x"C85F",
			x"0000" when x"C860",
			x"0000" when x"C861",
			x"0000" when x"C862",
			x"0000" when x"C863",
			x"0000" when x"C864",
			x"0000" when x"C865",
			x"0000" when x"C866",
			x"0000" when x"C867",
			x"0000" when x"C868",
			x"0000" when x"C869",
			x"0000" when x"C86A",
			x"0000" when x"C86B",
			x"0000" when x"C86C",
			x"0000" when x"C86D",
			x"0000" when x"C86E",
			x"0000" when x"C86F",
			x"0000" when x"C870",
			x"0000" when x"C871",
			x"0000" when x"C872",
			x"0000" when x"C873",
			x"0000" when x"C874",
			x"0000" when x"C875",
			x"0000" when x"C876",
			x"0000" when x"C877",
			x"0000" when x"C878",
			x"0000" when x"C879",
			x"0000" when x"C87A",
			x"0000" when x"C87B",
			x"0000" when x"C87C",
			x"0000" when x"C87D",
			x"0000" when x"C87E",
			x"0000" when x"C87F",
			x"0000" when x"C880",
			x"0000" when x"C881",
			x"0000" when x"C882",
			x"0000" when x"C883",
			x"0000" when x"C884",
			x"0000" when x"C885",
			x"0000" when x"C886",
			x"0000" when x"C887",
			x"0000" when x"C888",
			x"0000" when x"C889",
			x"0000" when x"C88A",
			x"0000" when x"C88B",
			x"0000" when x"C88C",
			x"0000" when x"C88D",
			x"0000" when x"C88E",
			x"0000" when x"C88F",
			x"0000" when x"C890",
			x"0000" when x"C891",
			x"0000" when x"C892",
			x"0000" when x"C893",
			x"0000" when x"C894",
			x"0000" when x"C895",
			x"0000" when x"C896",
			x"0000" when x"C897",
			x"0000" when x"C898",
			x"0000" when x"C899",
			x"0000" when x"C89A",
			x"0000" when x"C89B",
			x"0000" when x"C89C",
			x"0000" when x"C89D",
			x"0000" when x"C89E",
			x"0000" when x"C89F",
			x"0000" when x"C8A0",
			x"0000" when x"C8A1",
			x"0000" when x"C8A2",
			x"0000" when x"C8A3",
			x"0000" when x"C8A4",
			x"0000" when x"C8A5",
			x"0000" when x"C8A6",
			x"0000" when x"C8A7",
			x"0000" when x"C8A8",
			x"0000" when x"C8A9",
			x"0000" when x"C8AA",
			x"0000" when x"C8AB",
			x"0000" when x"C8AC",
			x"0000" when x"C8AD",
			x"0000" when x"C8AE",
			x"0000" when x"C8AF",
			x"0000" when x"C8B0",
			x"0000" when x"C8B1",
			x"0000" when x"C8B2",
			x"0000" when x"C8B3",
			x"0000" when x"C8B4",
			x"0000" when x"C8B5",
			x"0000" when x"C8B6",
			x"0000" when x"C8B7",
			x"0000" when x"C8B8",
			x"0000" when x"C8B9",
			x"0000" when x"C8BA",
			x"0000" when x"C8BB",
			x"0000" when x"C8BC",
			x"0000" when x"C8BD",
			x"0000" when x"C8BE",
			x"0000" when x"C8BF",
			x"0000" when x"C8C0",
			x"0000" when x"C8C1",
			x"0000" when x"C8C2",
			x"0000" when x"C8C3",
			x"0000" when x"C8C4",
			x"0000" when x"C8C5",
			x"0000" when x"C8C6",
			x"0000" when x"C8C7",
			x"0000" when x"C8C8",
			x"0000" when x"C8C9",
			x"0000" when x"C8CA",
			x"0000" when x"C8CB",
			x"0000" when x"C8CC",
			x"0000" when x"C8CD",
			x"0000" when x"C8CE",
			x"0000" when x"C8CF",
			x"0000" when x"C8D0",
			x"0000" when x"C8D1",
			x"0000" when x"C8D2",
			x"0000" when x"C8D3",
			x"0000" when x"C8D4",
			x"0000" when x"C8D5",
			x"0000" when x"C8D6",
			x"0000" when x"C8D7",
			x"0000" when x"C8D8",
			x"0000" when x"C8D9",
			x"0000" when x"C8DA",
			x"0000" when x"C8DB",
			x"0000" when x"C8DC",
			x"0000" when x"C8DD",
			x"0000" when x"C8DE",
			x"0000" when x"C8DF",
			x"0000" when x"C8E0",
			x"0000" when x"C8E1",
			x"0000" when x"C8E2",
			x"0000" when x"C8E3",
			x"0000" when x"C8E4",
			x"0000" when x"C8E5",
			x"0000" when x"C8E6",
			x"0000" when x"C8E7",
			x"0000" when x"C8E8",
			x"0000" when x"C8E9",
			x"0000" when x"C8EA",
			x"0000" when x"C8EB",
			x"0000" when x"C8EC",
			x"0000" when x"C8ED",
			x"0000" when x"C8EE",
			x"0000" when x"C8EF",
			x"0000" when x"C8F0",
			x"0000" when x"C8F1",
			x"0000" when x"C8F2",
			x"0000" when x"C8F3",
			x"0000" when x"C8F4",
			x"0000" when x"C8F5",
			x"0000" when x"C8F6",
			x"0000" when x"C8F7",
			x"0000" when x"C8F8",
			x"0000" when x"C8F9",
			x"0000" when x"C8FA",
			x"0000" when x"C8FB",
			x"0000" when x"C8FC",
			x"0000" when x"C8FD",
			x"0000" when x"C8FE",
			x"0000" when x"C8FF",
			x"0000" when x"C900",
			x"0000" when x"C901",
			x"0000" when x"C902",
			x"0000" when x"C903",
			x"0000" when x"C904",
			x"0000" when x"C905",
			x"0000" when x"C906",
			x"0000" when x"C907",
			x"0000" when x"C908",
			x"0000" when x"C909",
			x"0000" when x"C90A",
			x"0000" when x"C90B",
			x"0000" when x"C90C",
			x"0000" when x"C90D",
			x"0000" when x"C90E",
			x"0000" when x"C90F",
			x"0000" when x"C910",
			x"0000" when x"C911",
			x"0000" when x"C912",
			x"0000" when x"C913",
			x"0000" when x"C914",
			x"0000" when x"C915",
			x"0000" when x"C916",
			x"0000" when x"C917",
			x"0000" when x"C918",
			x"0000" when x"C919",
			x"0000" when x"C91A",
			x"0000" when x"C91B",
			x"0000" when x"C91C",
			x"0000" when x"C91D",
			x"0000" when x"C91E",
			x"0000" when x"C91F",
			x"0000" when x"C920",
			x"0000" when x"C921",
			x"0000" when x"C922",
			x"0000" when x"C923",
			x"0000" when x"C924",
			x"0000" when x"C925",
			x"0000" when x"C926",
			x"0000" when x"C927",
			x"0000" when x"C928",
			x"0000" when x"C929",
			x"0000" when x"C92A",
			x"0000" when x"C92B",
			x"0000" when x"C92C",
			x"0000" when x"C92D",
			x"0000" when x"C92E",
			x"0000" when x"C92F",
			x"0000" when x"C930",
			x"0000" when x"C931",
			x"0000" when x"C932",
			x"0000" when x"C933",
			x"0000" when x"C934",
			x"0000" when x"C935",
			x"0000" when x"C936",
			x"0000" when x"C937",
			x"0000" when x"C938",
			x"0000" when x"C939",
			x"0000" when x"C93A",
			x"0000" when x"C93B",
			x"0000" when x"C93C",
			x"0000" when x"C93D",
			x"0000" when x"C93E",
			x"0000" when x"C93F",
			x"0000" when x"C940",
			x"0000" when x"C941",
			x"0000" when x"C942",
			x"0000" when x"C943",
			x"0000" when x"C944",
			x"0000" when x"C945",
			x"0000" when x"C946",
			x"0000" when x"C947",
			x"0000" when x"C948",
			x"0000" when x"C949",
			x"0000" when x"C94A",
			x"0000" when x"C94B",
			x"0000" when x"C94C",
			x"0000" when x"C94D",
			x"0000" when x"C94E",
			x"0000" when x"C94F",
			x"0000" when x"C950",
			x"0000" when x"C951",
			x"0000" when x"C952",
			x"0000" when x"C953",
			x"0000" when x"C954",
			x"0000" when x"C955",
			x"0000" when x"C956",
			x"0000" when x"C957",
			x"0000" when x"C958",
			x"0000" when x"C959",
			x"0000" when x"C95A",
			x"0000" when x"C95B",
			x"0000" when x"C95C",
			x"0000" when x"C95D",
			x"0000" when x"C95E",
			x"0000" when x"C95F",
			x"0000" when x"C960",
			x"0000" when x"C961",
			x"0000" when x"C962",
			x"0000" when x"C963",
			x"0000" when x"C964",
			x"0000" when x"C965",
			x"0000" when x"C966",
			x"0000" when x"C967",
			x"0000" when x"C968",
			x"0000" when x"C969",
			x"0000" when x"C96A",
			x"0000" when x"C96B",
			x"0000" when x"C96C",
			x"0000" when x"C96D",
			x"0000" when x"C96E",
			x"0000" when x"C96F",
			x"0000" when x"C970",
			x"0000" when x"C971",
			x"0000" when x"C972",
			x"0000" when x"C973",
			x"0000" when x"C974",
			x"0000" when x"C975",
			x"0000" when x"C976",
			x"0000" when x"C977",
			x"0000" when x"C978",
			x"0000" when x"C979",
			x"0000" when x"C97A",
			x"0000" when x"C97B",
			x"0000" when x"C97C",
			x"0000" when x"C97D",
			x"0000" when x"C97E",
			x"0000" when x"C97F",
			x"0000" when x"C980",
			x"0000" when x"C981",
			x"0000" when x"C982",
			x"0000" when x"C983",
			x"0000" when x"C984",
			x"0000" when x"C985",
			x"0000" when x"C986",
			x"0000" when x"C987",
			x"0000" when x"C988",
			x"0000" when x"C989",
			x"0000" when x"C98A",
			x"0000" when x"C98B",
			x"0000" when x"C98C",
			x"0000" when x"C98D",
			x"0000" when x"C98E",
			x"0000" when x"C98F",
			x"0000" when x"C990",
			x"0000" when x"C991",
			x"0000" when x"C992",
			x"0000" when x"C993",
			x"0000" when x"C994",
			x"0000" when x"C995",
			x"0000" when x"C996",
			x"0000" when x"C997",
			x"0000" when x"C998",
			x"0000" when x"C999",
			x"0000" when x"C99A",
			x"0000" when x"C99B",
			x"0000" when x"C99C",
			x"0000" when x"C99D",
			x"0000" when x"C99E",
			x"0000" when x"C99F",
			x"0000" when x"C9A0",
			x"0000" when x"C9A1",
			x"0000" when x"C9A2",
			x"0000" when x"C9A3",
			x"0000" when x"C9A4",
			x"0000" when x"C9A5",
			x"0000" when x"C9A6",
			x"0000" when x"C9A7",
			x"0000" when x"C9A8",
			x"0000" when x"C9A9",
			x"0000" when x"C9AA",
			x"0000" when x"C9AB",
			x"0000" when x"C9AC",
			x"0000" when x"C9AD",
			x"0000" when x"C9AE",
			x"0000" when x"C9AF",
			x"0000" when x"C9B0",
			x"0000" when x"C9B1",
			x"0000" when x"C9B2",
			x"0000" when x"C9B3",
			x"0000" when x"C9B4",
			x"0000" when x"C9B5",
			x"0000" when x"C9B6",
			x"0000" when x"C9B7",
			x"0000" when x"C9B8",
			x"0000" when x"C9B9",
			x"0000" when x"C9BA",
			x"0000" when x"C9BB",
			x"0000" when x"C9BC",
			x"0000" when x"C9BD",
			x"0000" when x"C9BE",
			x"0000" when x"C9BF",
			x"0000" when x"C9C0",
			x"0000" when x"C9C1",
			x"0000" when x"C9C2",
			x"0000" when x"C9C3",
			x"0000" when x"C9C4",
			x"0000" when x"C9C5",
			x"0000" when x"C9C6",
			x"0000" when x"C9C7",
			x"0000" when x"C9C8",
			x"0000" when x"C9C9",
			x"0000" when x"C9CA",
			x"0000" when x"C9CB",
			x"0000" when x"C9CC",
			x"0000" when x"C9CD",
			x"0000" when x"C9CE",
			x"0000" when x"C9CF",
			x"0000" when x"C9D0",
			x"0000" when x"C9D1",
			x"0000" when x"C9D2",
			x"0000" when x"C9D3",
			x"0000" when x"C9D4",
			x"0000" when x"C9D5",
			x"0000" when x"C9D6",
			x"0000" when x"C9D7",
			x"0000" when x"C9D8",
			x"0000" when x"C9D9",
			x"0000" when x"C9DA",
			x"0000" when x"C9DB",
			x"0000" when x"C9DC",
			x"0000" when x"C9DD",
			x"0000" when x"C9DE",
			x"0000" when x"C9DF",
			x"0000" when x"C9E0",
			x"0000" when x"C9E1",
			x"0000" when x"C9E2",
			x"0000" when x"C9E3",
			x"0000" when x"C9E4",
			x"0000" when x"C9E5",
			x"0000" when x"C9E6",
			x"0000" when x"C9E7",
			x"0000" when x"C9E8",
			x"0000" when x"C9E9",
			x"0000" when x"C9EA",
			x"0000" when x"C9EB",
			x"0000" when x"C9EC",
			x"0000" when x"C9ED",
			x"0000" when x"C9EE",
			x"0000" when x"C9EF",
			x"0000" when x"C9F0",
			x"0000" when x"C9F1",
			x"0000" when x"C9F2",
			x"0000" when x"C9F3",
			x"0000" when x"C9F4",
			x"0000" when x"C9F5",
			x"0000" when x"C9F6",
			x"0000" when x"C9F7",
			x"0000" when x"C9F8",
			x"0000" when x"C9F9",
			x"0000" when x"C9FA",
			x"0000" when x"C9FB",
			x"0000" when x"C9FC",
			x"0000" when x"C9FD",
			x"0000" when x"C9FE",
			x"0000" when x"C9FF",
			x"0000" when x"CA00",
			x"0000" when x"CA01",
			x"0000" when x"CA02",
			x"0000" when x"CA03",
			x"0000" when x"CA04",
			x"0000" when x"CA05",
			x"0000" when x"CA06",
			x"0000" when x"CA07",
			x"0000" when x"CA08",
			x"0000" when x"CA09",
			x"0000" when x"CA0A",
			x"0000" when x"CA0B",
			x"0000" when x"CA0C",
			x"0000" when x"CA0D",
			x"0000" when x"CA0E",
			x"0000" when x"CA0F",
			x"0000" when x"CA10",
			x"0000" when x"CA11",
			x"0000" when x"CA12",
			x"0000" when x"CA13",
			x"0000" when x"CA14",
			x"0000" when x"CA15",
			x"0000" when x"CA16",
			x"0000" when x"CA17",
			x"0000" when x"CA18",
			x"0000" when x"CA19",
			x"0000" when x"CA1A",
			x"0000" when x"CA1B",
			x"0000" when x"CA1C",
			x"0000" when x"CA1D",
			x"0000" when x"CA1E",
			x"0000" when x"CA1F",
			x"0000" when x"CA20",
			x"0000" when x"CA21",
			x"0000" when x"CA22",
			x"0000" when x"CA23",
			x"0000" when x"CA24",
			x"0000" when x"CA25",
			x"0000" when x"CA26",
			x"0000" when x"CA27",
			x"0000" when x"CA28",
			x"0000" when x"CA29",
			x"0000" when x"CA2A",
			x"0000" when x"CA2B",
			x"0000" when x"CA2C",
			x"0000" when x"CA2D",
			x"0000" when x"CA2E",
			x"0000" when x"CA2F",
			x"0000" when x"CA30",
			x"0000" when x"CA31",
			x"0000" when x"CA32",
			x"0000" when x"CA33",
			x"0000" when x"CA34",
			x"0000" when x"CA35",
			x"0000" when x"CA36",
			x"0000" when x"CA37",
			x"0000" when x"CA38",
			x"0000" when x"CA39",
			x"0000" when x"CA3A",
			x"0000" when x"CA3B",
			x"0000" when x"CA3C",
			x"0000" when x"CA3D",
			x"0000" when x"CA3E",
			x"0000" when x"CA3F",
			x"0000" when x"CA40",
			x"0000" when x"CA41",
			x"0000" when x"CA42",
			x"0000" when x"CA43",
			x"0000" when x"CA44",
			x"0000" when x"CA45",
			x"0000" when x"CA46",
			x"0000" when x"CA47",
			x"0000" when x"CA48",
			x"0000" when x"CA49",
			x"0000" when x"CA4A",
			x"0000" when x"CA4B",
			x"0000" when x"CA4C",
			x"0000" when x"CA4D",
			x"0000" when x"CA4E",
			x"0000" when x"CA4F",
			x"0000" when x"CA50",
			x"0000" when x"CA51",
			x"0000" when x"CA52",
			x"0000" when x"CA53",
			x"0000" when x"CA54",
			x"0000" when x"CA55",
			x"0000" when x"CA56",
			x"0000" when x"CA57",
			x"0000" when x"CA58",
			x"0000" when x"CA59",
			x"0000" when x"CA5A",
			x"0000" when x"CA5B",
			x"0000" when x"CA5C",
			x"0000" when x"CA5D",
			x"0000" when x"CA5E",
			x"0000" when x"CA5F",
			x"0000" when x"CA60",
			x"0000" when x"CA61",
			x"0000" when x"CA62",
			x"0000" when x"CA63",
			x"0000" when x"CA64",
			x"0000" when x"CA65",
			x"0000" when x"CA66",
			x"0000" when x"CA67",
			x"0000" when x"CA68",
			x"0000" when x"CA69",
			x"0000" when x"CA6A",
			x"0000" when x"CA6B",
			x"0000" when x"CA6C",
			x"0000" when x"CA6D",
			x"0000" when x"CA6E",
			x"0000" when x"CA6F",
			x"0000" when x"CA70",
			x"0000" when x"CA71",
			x"0000" when x"CA72",
			x"0000" when x"CA73",
			x"0000" when x"CA74",
			x"0000" when x"CA75",
			x"0000" when x"CA76",
			x"0000" when x"CA77",
			x"0000" when x"CA78",
			x"0000" when x"CA79",
			x"0000" when x"CA7A",
			x"0000" when x"CA7B",
			x"0000" when x"CA7C",
			x"0000" when x"CA7D",
			x"0000" when x"CA7E",
			x"0000" when x"CA7F",
			x"0000" when x"CA80",
			x"0000" when x"CA81",
			x"0000" when x"CA82",
			x"0000" when x"CA83",
			x"0000" when x"CA84",
			x"0000" when x"CA85",
			x"0000" when x"CA86",
			x"0000" when x"CA87",
			x"0000" when x"CA88",
			x"0000" when x"CA89",
			x"0000" when x"CA8A",
			x"0000" when x"CA8B",
			x"0000" when x"CA8C",
			x"0000" when x"CA8D",
			x"0000" when x"CA8E",
			x"0000" when x"CA8F",
			x"0000" when x"CA90",
			x"0000" when x"CA91",
			x"0000" when x"CA92",
			x"0000" when x"CA93",
			x"0000" when x"CA94",
			x"0000" when x"CA95",
			x"0000" when x"CA96",
			x"0000" when x"CA97",
			x"0000" when x"CA98",
			x"0000" when x"CA99",
			x"0000" when x"CA9A",
			x"0000" when x"CA9B",
			x"0000" when x"CA9C",
			x"0000" when x"CA9D",
			x"0000" when x"CA9E",
			x"0000" when x"CA9F",
			x"0000" when x"CAA0",
			x"0000" when x"CAA1",
			x"0000" when x"CAA2",
			x"0000" when x"CAA3",
			x"0000" when x"CAA4",
			x"0000" when x"CAA5",
			x"0000" when x"CAA6",
			x"0000" when x"CAA7",
			x"0000" when x"CAA8",
			x"0000" when x"CAA9",
			x"0000" when x"CAAA",
			x"0000" when x"CAAB",
			x"0000" when x"CAAC",
			x"0000" when x"CAAD",
			x"0000" when x"CAAE",
			x"0000" when x"CAAF",
			x"0000" when x"CAB0",
			x"0000" when x"CAB1",
			x"0000" when x"CAB2",
			x"0000" when x"CAB3",
			x"0000" when x"CAB4",
			x"0000" when x"CAB5",
			x"0000" when x"CAB6",
			x"0000" when x"CAB7",
			x"0000" when x"CAB8",
			x"0000" when x"CAB9",
			x"0000" when x"CABA",
			x"0000" when x"CABB",
			x"0000" when x"CABC",
			x"0000" when x"CABD",
			x"0000" when x"CABE",
			x"0000" when x"CABF",
			x"0000" when x"CAC0",
			x"0000" when x"CAC1",
			x"0000" when x"CAC2",
			x"0000" when x"CAC3",
			x"0000" when x"CAC4",
			x"0000" when x"CAC5",
			x"0000" when x"CAC6",
			x"0000" when x"CAC7",
			x"0000" when x"CAC8",
			x"0000" when x"CAC9",
			x"0000" when x"CACA",
			x"0000" when x"CACB",
			x"0000" when x"CACC",
			x"0000" when x"CACD",
			x"0000" when x"CACE",
			x"0000" when x"CACF",
			x"0000" when x"CAD0",
			x"0000" when x"CAD1",
			x"0000" when x"CAD2",
			x"0000" when x"CAD3",
			x"0000" when x"CAD4",
			x"0000" when x"CAD5",
			x"0000" when x"CAD6",
			x"0000" when x"CAD7",
			x"0000" when x"CAD8",
			x"0000" when x"CAD9",
			x"0000" when x"CADA",
			x"0000" when x"CADB",
			x"0000" when x"CADC",
			x"0000" when x"CADD",
			x"0000" when x"CADE",
			x"0000" when x"CADF",
			x"0000" when x"CAE0",
			x"0000" when x"CAE1",
			x"0000" when x"CAE2",
			x"0000" when x"CAE3",
			x"0000" when x"CAE4",
			x"0000" when x"CAE5",
			x"0000" when x"CAE6",
			x"0000" when x"CAE7",
			x"0000" when x"CAE8",
			x"0000" when x"CAE9",
			x"0000" when x"CAEA",
			x"0000" when x"CAEB",
			x"0000" when x"CAEC",
			x"0000" when x"CAED",
			x"0000" when x"CAEE",
			x"0000" when x"CAEF",
			x"0000" when x"CAF0",
			x"0000" when x"CAF1",
			x"0000" when x"CAF2",
			x"0000" when x"CAF3",
			x"0000" when x"CAF4",
			x"0000" when x"CAF5",
			x"0000" when x"CAF6",
			x"0000" when x"CAF7",
			x"0000" when x"CAF8",
			x"0000" when x"CAF9",
			x"0000" when x"CAFA",
			x"0000" when x"CAFB",
			x"0000" when x"CAFC",
			x"0000" when x"CAFD",
			x"0000" when x"CAFE",
			x"0000" when x"CAFF",
			x"0000" when x"CB00",
			x"0000" when x"CB01",
			x"0000" when x"CB02",
			x"0000" when x"CB03",
			x"0000" when x"CB04",
			x"0000" when x"CB05",
			x"0000" when x"CB06",
			x"0000" when x"CB07",
			x"0000" when x"CB08",
			x"0000" when x"CB09",
			x"0000" when x"CB0A",
			x"0000" when x"CB0B",
			x"0000" when x"CB0C",
			x"0000" when x"CB0D",
			x"0000" when x"CB0E",
			x"0000" when x"CB0F",
			x"0000" when x"CB10",
			x"0000" when x"CB11",
			x"0000" when x"CB12",
			x"0000" when x"CB13",
			x"0000" when x"CB14",
			x"0000" when x"CB15",
			x"0000" when x"CB16",
			x"0000" when x"CB17",
			x"0000" when x"CB18",
			x"0000" when x"CB19",
			x"0000" when x"CB1A",
			x"0000" when x"CB1B",
			x"0000" when x"CB1C",
			x"0000" when x"CB1D",
			x"0000" when x"CB1E",
			x"0000" when x"CB1F",
			x"0000" when x"CB20",
			x"0000" when x"CB21",
			x"0000" when x"CB22",
			x"0000" when x"CB23",
			x"0000" when x"CB24",
			x"0000" when x"CB25",
			x"0000" when x"CB26",
			x"0000" when x"CB27",
			x"0000" when x"CB28",
			x"0000" when x"CB29",
			x"0000" when x"CB2A",
			x"0000" when x"CB2B",
			x"0000" when x"CB2C",
			x"0000" when x"CB2D",
			x"0000" when x"CB2E",
			x"0000" when x"CB2F",
			x"0000" when x"CB30",
			x"0000" when x"CB31",
			x"0000" when x"CB32",
			x"0000" when x"CB33",
			x"0000" when x"CB34",
			x"0000" when x"CB35",
			x"0000" when x"CB36",
			x"0000" when x"CB37",
			x"0000" when x"CB38",
			x"0000" when x"CB39",
			x"0000" when x"CB3A",
			x"0000" when x"CB3B",
			x"0000" when x"CB3C",
			x"0000" when x"CB3D",
			x"0000" when x"CB3E",
			x"0000" when x"CB3F",
			x"0000" when x"CB40",
			x"0000" when x"CB41",
			x"0000" when x"CB42",
			x"0000" when x"CB43",
			x"0000" when x"CB44",
			x"0000" when x"CB45",
			x"0000" when x"CB46",
			x"0000" when x"CB47",
			x"0000" when x"CB48",
			x"0000" when x"CB49",
			x"0000" when x"CB4A",
			x"0000" when x"CB4B",
			x"0000" when x"CB4C",
			x"0000" when x"CB4D",
			x"0000" when x"CB4E",
			x"0000" when x"CB4F",
			x"0000" when x"CB50",
			x"0000" when x"CB51",
			x"0000" when x"CB52",
			x"0000" when x"CB53",
			x"0000" when x"CB54",
			x"0000" when x"CB55",
			x"0000" when x"CB56",
			x"0000" when x"CB57",
			x"0000" when x"CB58",
			x"0000" when x"CB59",
			x"0000" when x"CB5A",
			x"0000" when x"CB5B",
			x"0000" when x"CB5C",
			x"0000" when x"CB5D",
			x"0000" when x"CB5E",
			x"0000" when x"CB5F",
			x"0000" when x"CB60",
			x"0000" when x"CB61",
			x"0000" when x"CB62",
			x"0000" when x"CB63",
			x"0000" when x"CB64",
			x"0000" when x"CB65",
			x"0000" when x"CB66",
			x"0000" when x"CB67",
			x"0000" when x"CB68",
			x"0000" when x"CB69",
			x"0000" when x"CB6A",
			x"0000" when x"CB6B",
			x"0000" when x"CB6C",
			x"0000" when x"CB6D",
			x"0000" when x"CB6E",
			x"0000" when x"CB6F",
			x"0000" when x"CB70",
			x"0000" when x"CB71",
			x"0000" when x"CB72",
			x"0000" when x"CB73",
			x"0000" when x"CB74",
			x"0000" when x"CB75",
			x"0000" when x"CB76",
			x"0000" when x"CB77",
			x"0000" when x"CB78",
			x"0000" when x"CB79",
			x"0000" when x"CB7A",
			x"0000" when x"CB7B",
			x"0000" when x"CB7C",
			x"0000" when x"CB7D",
			x"0000" when x"CB7E",
			x"0000" when x"CB7F",
			x"0000" when x"CB80",
			x"0000" when x"CB81",
			x"0000" when x"CB82",
			x"0000" when x"CB83",
			x"0000" when x"CB84",
			x"0000" when x"CB85",
			x"0000" when x"CB86",
			x"0000" when x"CB87",
			x"0000" when x"CB88",
			x"0000" when x"CB89",
			x"0000" when x"CB8A",
			x"0000" when x"CB8B",
			x"0000" when x"CB8C",
			x"0000" when x"CB8D",
			x"0000" when x"CB8E",
			x"0000" when x"CB8F",
			x"0000" when x"CB90",
			x"0000" when x"CB91",
			x"0000" when x"CB92",
			x"0000" when x"CB93",
			x"0000" when x"CB94",
			x"0000" when x"CB95",
			x"0000" when x"CB96",
			x"0000" when x"CB97",
			x"0000" when x"CB98",
			x"0000" when x"CB99",
			x"0000" when x"CB9A",
			x"0000" when x"CB9B",
			x"0000" when x"CB9C",
			x"0000" when x"CB9D",
			x"0000" when x"CB9E",
			x"0000" when x"CB9F",
			x"0000" when x"CBA0",
			x"0000" when x"CBA1",
			x"0000" when x"CBA2",
			x"0000" when x"CBA3",
			x"0000" when x"CBA4",
			x"0000" when x"CBA5",
			x"0000" when x"CBA6",
			x"0000" when x"CBA7",
			x"0000" when x"CBA8",
			x"0000" when x"CBA9",
			x"0000" when x"CBAA",
			x"0000" when x"CBAB",
			x"0000" when x"CBAC",
			x"0000" when x"CBAD",
			x"0000" when x"CBAE",
			x"0000" when x"CBAF",
			x"0000" when x"CBB0",
			x"0000" when x"CBB1",
			x"0000" when x"CBB2",
			x"0000" when x"CBB3",
			x"0000" when x"CBB4",
			x"0000" when x"CBB5",
			x"0000" when x"CBB6",
			x"0000" when x"CBB7",
			x"0000" when x"CBB8",
			x"0000" when x"CBB9",
			x"0000" when x"CBBA",
			x"0000" when x"CBBB",
			x"0000" when x"CBBC",
			x"0000" when x"CBBD",
			x"0000" when x"CBBE",
			x"0000" when x"CBBF",
			x"0000" when x"CBC0",
			x"0000" when x"CBC1",
			x"0000" when x"CBC2",
			x"0000" when x"CBC3",
			x"0000" when x"CBC4",
			x"0000" when x"CBC5",
			x"0000" when x"CBC6",
			x"0000" when x"CBC7",
			x"0000" when x"CBC8",
			x"0000" when x"CBC9",
			x"0000" when x"CBCA",
			x"0000" when x"CBCB",
			x"0000" when x"CBCC",
			x"0000" when x"CBCD",
			x"0000" when x"CBCE",
			x"0000" when x"CBCF",
			x"0000" when x"CBD0",
			x"0000" when x"CBD1",
			x"0000" when x"CBD2",
			x"0000" when x"CBD3",
			x"0000" when x"CBD4",
			x"0000" when x"CBD5",
			x"0000" when x"CBD6",
			x"0000" when x"CBD7",
			x"0000" when x"CBD8",
			x"0000" when x"CBD9",
			x"0000" when x"CBDA",
			x"0000" when x"CBDB",
			x"0000" when x"CBDC",
			x"0000" when x"CBDD",
			x"0000" when x"CBDE",
			x"0000" when x"CBDF",
			x"0000" when x"CBE0",
			x"0000" when x"CBE1",
			x"0000" when x"CBE2",
			x"0000" when x"CBE3",
			x"0000" when x"CBE4",
			x"0000" when x"CBE5",
			x"0000" when x"CBE6",
			x"0000" when x"CBE7",
			x"0000" when x"CBE8",
			x"0000" when x"CBE9",
			x"0000" when x"CBEA",
			x"0000" when x"CBEB",
			x"0000" when x"CBEC",
			x"0000" when x"CBED",
			x"0000" when x"CBEE",
			x"0000" when x"CBEF",
			x"0000" when x"CBF0",
			x"0000" when x"CBF1",
			x"0000" when x"CBF2",
			x"0000" when x"CBF3",
			x"0000" when x"CBF4",
			x"0000" when x"CBF5",
			x"0000" when x"CBF6",
			x"0000" when x"CBF7",
			x"0000" when x"CBF8",
			x"0000" when x"CBF9",
			x"0000" when x"CBFA",
			x"0000" when x"CBFB",
			x"0000" when x"CBFC",
			x"0000" when x"CBFD",
			x"0000" when x"CBFE",
			x"0000" when x"CBFF",
			x"0000" when x"CC00",
			x"0000" when x"CC01",
			x"0000" when x"CC02",
			x"0000" when x"CC03",
			x"0000" when x"CC04",
			x"0000" when x"CC05",
			x"0000" when x"CC06",
			x"0000" when x"CC07",
			x"0000" when x"CC08",
			x"0000" when x"CC09",
			x"0000" when x"CC0A",
			x"0000" when x"CC0B",
			x"0000" when x"CC0C",
			x"0000" when x"CC0D",
			x"0000" when x"CC0E",
			x"0000" when x"CC0F",
			x"0000" when x"CC10",
			x"0000" when x"CC11",
			x"0000" when x"CC12",
			x"0000" when x"CC13",
			x"0000" when x"CC14",
			x"0000" when x"CC15",
			x"0000" when x"CC16",
			x"0000" when x"CC17",
			x"0000" when x"CC18",
			x"0000" when x"CC19",
			x"0000" when x"CC1A",
			x"0000" when x"CC1B",
			x"0000" when x"CC1C",
			x"0000" when x"CC1D",
			x"0000" when x"CC1E",
			x"0000" when x"CC1F",
			x"0000" when x"CC20",
			x"0000" when x"CC21",
			x"0000" when x"CC22",
			x"0000" when x"CC23",
			x"0000" when x"CC24",
			x"0000" when x"CC25",
			x"0000" when x"CC26",
			x"0000" when x"CC27",
			x"0000" when x"CC28",
			x"0000" when x"CC29",
			x"0000" when x"CC2A",
			x"0000" when x"CC2B",
			x"0000" when x"CC2C",
			x"0000" when x"CC2D",
			x"0000" when x"CC2E",
			x"0000" when x"CC2F",
			x"0000" when x"CC30",
			x"0000" when x"CC31",
			x"0000" when x"CC32",
			x"0000" when x"CC33",
			x"0000" when x"CC34",
			x"0000" when x"CC35",
			x"0000" when x"CC36",
			x"0000" when x"CC37",
			x"0000" when x"CC38",
			x"0000" when x"CC39",
			x"0000" when x"CC3A",
			x"0000" when x"CC3B",
			x"0000" when x"CC3C",
			x"0000" when x"CC3D",
			x"0000" when x"CC3E",
			x"0000" when x"CC3F",
			x"0000" when x"CC40",
			x"0000" when x"CC41",
			x"0000" when x"CC42",
			x"0000" when x"CC43",
			x"0000" when x"CC44",
			x"0000" when x"CC45",
			x"0000" when x"CC46",
			x"0000" when x"CC47",
			x"0000" when x"CC48",
			x"0000" when x"CC49",
			x"0000" when x"CC4A",
			x"0000" when x"CC4B",
			x"0000" when x"CC4C",
			x"0000" when x"CC4D",
			x"0000" when x"CC4E",
			x"0000" when x"CC4F",
			x"0000" when x"CC50",
			x"0000" when x"CC51",
			x"0000" when x"CC52",
			x"0000" when x"CC53",
			x"0000" when x"CC54",
			x"0000" when x"CC55",
			x"0000" when x"CC56",
			x"0000" when x"CC57",
			x"0000" when x"CC58",
			x"0000" when x"CC59",
			x"0000" when x"CC5A",
			x"0000" when x"CC5B",
			x"0000" when x"CC5C",
			x"0000" when x"CC5D",
			x"0000" when x"CC5E",
			x"0000" when x"CC5F",
			x"0000" when x"CC60",
			x"0000" when x"CC61",
			x"0000" when x"CC62",
			x"0000" when x"CC63",
			x"0000" when x"CC64",
			x"0000" when x"CC65",
			x"0000" when x"CC66",
			x"0000" when x"CC67",
			x"0000" when x"CC68",
			x"0000" when x"CC69",
			x"0000" when x"CC6A",
			x"0000" when x"CC6B",
			x"0000" when x"CC6C",
			x"0000" when x"CC6D",
			x"0000" when x"CC6E",
			x"0000" when x"CC6F",
			x"0000" when x"CC70",
			x"0000" when x"CC71",
			x"0000" when x"CC72",
			x"0000" when x"CC73",
			x"0000" when x"CC74",
			x"0000" when x"CC75",
			x"0000" when x"CC76",
			x"0000" when x"CC77",
			x"0000" when x"CC78",
			x"0000" when x"CC79",
			x"0000" when x"CC7A",
			x"0000" when x"CC7B",
			x"0000" when x"CC7C",
			x"0000" when x"CC7D",
			x"0000" when x"CC7E",
			x"0000" when x"CC7F",
			x"0000" when x"CC80",
			x"0000" when x"CC81",
			x"0000" when x"CC82",
			x"0000" when x"CC83",
			x"0000" when x"CC84",
			x"0000" when x"CC85",
			x"0000" when x"CC86",
			x"0000" when x"CC87",
			x"0000" when x"CC88",
			x"0000" when x"CC89",
			x"0000" when x"CC8A",
			x"0000" when x"CC8B",
			x"0000" when x"CC8C",
			x"0000" when x"CC8D",
			x"0000" when x"CC8E",
			x"0000" when x"CC8F",
			x"0000" when x"CC90",
			x"0000" when x"CC91",
			x"0000" when x"CC92",
			x"0000" when x"CC93",
			x"0000" when x"CC94",
			x"0000" when x"CC95",
			x"0000" when x"CC96",
			x"0000" when x"CC97",
			x"0000" when x"CC98",
			x"0000" when x"CC99",
			x"0000" when x"CC9A",
			x"0000" when x"CC9B",
			x"0000" when x"CC9C",
			x"0000" when x"CC9D",
			x"0000" when x"CC9E",
			x"0000" when x"CC9F",
			x"0000" when x"CCA0",
			x"0000" when x"CCA1",
			x"0000" when x"CCA2",
			x"0000" when x"CCA3",
			x"0000" when x"CCA4",
			x"0000" when x"CCA5",
			x"0000" when x"CCA6",
			x"0000" when x"CCA7",
			x"0000" when x"CCA8",
			x"0000" when x"CCA9",
			x"0000" when x"CCAA",
			x"0000" when x"CCAB",
			x"0000" when x"CCAC",
			x"0000" when x"CCAD",
			x"0000" when x"CCAE",
			x"0000" when x"CCAF",
			x"0000" when x"CCB0",
			x"0000" when x"CCB1",
			x"0000" when x"CCB2",
			x"0000" when x"CCB3",
			x"0000" when x"CCB4",
			x"0000" when x"CCB5",
			x"0000" when x"CCB6",
			x"0000" when x"CCB7",
			x"0000" when x"CCB8",
			x"0000" when x"CCB9",
			x"0000" when x"CCBA",
			x"0000" when x"CCBB",
			x"0000" when x"CCBC",
			x"0000" when x"CCBD",
			x"0000" when x"CCBE",
			x"0000" when x"CCBF",
			x"0000" when x"CCC0",
			x"0000" when x"CCC1",
			x"0000" when x"CCC2",
			x"0000" when x"CCC3",
			x"0000" when x"CCC4",
			x"0000" when x"CCC5",
			x"0000" when x"CCC6",
			x"0000" when x"CCC7",
			x"0000" when x"CCC8",
			x"0000" when x"CCC9",
			x"0000" when x"CCCA",
			x"0000" when x"CCCB",
			x"0000" when x"CCCC",
			x"0000" when x"CCCD",
			x"0000" when x"CCCE",
			x"0000" when x"CCCF",
			x"0000" when x"CCD0",
			x"0000" when x"CCD1",
			x"0000" when x"CCD2",
			x"0000" when x"CCD3",
			x"0000" when x"CCD4",
			x"0000" when x"CCD5",
			x"0000" when x"CCD6",
			x"0000" when x"CCD7",
			x"0000" when x"CCD8",
			x"0000" when x"CCD9",
			x"0000" when x"CCDA",
			x"0000" when x"CCDB",
			x"0000" when x"CCDC",
			x"0000" when x"CCDD",
			x"0000" when x"CCDE",
			x"0000" when x"CCDF",
			x"0000" when x"CCE0",
			x"0000" when x"CCE1",
			x"0000" when x"CCE2",
			x"0000" when x"CCE3",
			x"0000" when x"CCE4",
			x"0000" when x"CCE5",
			x"0000" when x"CCE6",
			x"0000" when x"CCE7",
			x"0000" when x"CCE8",
			x"0000" when x"CCE9",
			x"0000" when x"CCEA",
			x"0000" when x"CCEB",
			x"0000" when x"CCEC",
			x"0000" when x"CCED",
			x"0000" when x"CCEE",
			x"0000" when x"CCEF",
			x"0000" when x"CCF0",
			x"0000" when x"CCF1",
			x"0000" when x"CCF2",
			x"0000" when x"CCF3",
			x"0000" when x"CCF4",
			x"0000" when x"CCF5",
			x"0000" when x"CCF6",
			x"0000" when x"CCF7",
			x"0000" when x"CCF8",
			x"0000" when x"CCF9",
			x"0000" when x"CCFA",
			x"0000" when x"CCFB",
			x"0000" when x"CCFC",
			x"0000" when x"CCFD",
			x"0000" when x"CCFE",
			x"0000" when x"CCFF",
			x"0000" when x"CD00",
			x"0000" when x"CD01",
			x"0000" when x"CD02",
			x"0000" when x"CD03",
			x"0000" when x"CD04",
			x"0000" when x"CD05",
			x"0000" when x"CD06",
			x"0000" when x"CD07",
			x"0000" when x"CD08",
			x"0000" when x"CD09",
			x"0000" when x"CD0A",
			x"0000" when x"CD0B",
			x"0000" when x"CD0C",
			x"0000" when x"CD0D",
			x"0000" when x"CD0E",
			x"0000" when x"CD0F",
			x"0000" when x"CD10",
			x"0000" when x"CD11",
			x"0000" when x"CD12",
			x"0000" when x"CD13",
			x"0000" when x"CD14",
			x"0000" when x"CD15",
			x"0000" when x"CD16",
			x"0000" when x"CD17",
			x"0000" when x"CD18",
			x"0000" when x"CD19",
			x"0000" when x"CD1A",
			x"0000" when x"CD1B",
			x"0000" when x"CD1C",
			x"0000" when x"CD1D",
			x"0000" when x"CD1E",
			x"0000" when x"CD1F",
			x"0000" when x"CD20",
			x"0000" when x"CD21",
			x"0000" when x"CD22",
			x"0000" when x"CD23",
			x"0000" when x"CD24",
			x"0000" when x"CD25",
			x"0000" when x"CD26",
			x"0000" when x"CD27",
			x"0000" when x"CD28",
			x"0000" when x"CD29",
			x"0000" when x"CD2A",
			x"0000" when x"CD2B",
			x"0000" when x"CD2C",
			x"0000" when x"CD2D",
			x"0000" when x"CD2E",
			x"0000" when x"CD2F",
			x"0000" when x"CD30",
			x"0000" when x"CD31",
			x"0000" when x"CD32",
			x"0000" when x"CD33",
			x"0000" when x"CD34",
			x"0000" when x"CD35",
			x"0000" when x"CD36",
			x"0000" when x"CD37",
			x"0000" when x"CD38",
			x"0000" when x"CD39",
			x"0000" when x"CD3A",
			x"0000" when x"CD3B",
			x"0000" when x"CD3C",
			x"0000" when x"CD3D",
			x"0000" when x"CD3E",
			x"0000" when x"CD3F",
			x"0000" when x"CD40",
			x"0000" when x"CD41",
			x"0000" when x"CD42",
			x"0000" when x"CD43",
			x"0000" when x"CD44",
			x"0000" when x"CD45",
			x"0000" when x"CD46",
			x"0000" when x"CD47",
			x"0000" when x"CD48",
			x"0000" when x"CD49",
			x"0000" when x"CD4A",
			x"0000" when x"CD4B",
			x"0000" when x"CD4C",
			x"0000" when x"CD4D",
			x"0000" when x"CD4E",
			x"0000" when x"CD4F",
			x"0000" when x"CD50",
			x"0000" when x"CD51",
			x"0000" when x"CD52",
			x"0000" when x"CD53",
			x"0000" when x"CD54",
			x"0000" when x"CD55",
			x"0000" when x"CD56",
			x"0000" when x"CD57",
			x"0000" when x"CD58",
			x"0000" when x"CD59",
			x"0000" when x"CD5A",
			x"0000" when x"CD5B",
			x"0000" when x"CD5C",
			x"0000" when x"CD5D",
			x"0000" when x"CD5E",
			x"0000" when x"CD5F",
			x"0000" when x"CD60",
			x"0000" when x"CD61",
			x"0000" when x"CD62",
			x"0000" when x"CD63",
			x"0000" when x"CD64",
			x"0000" when x"CD65",
			x"0000" when x"CD66",
			x"0000" when x"CD67",
			x"0000" when x"CD68",
			x"0000" when x"CD69",
			x"0000" when x"CD6A",
			x"0000" when x"CD6B",
			x"0000" when x"CD6C",
			x"0000" when x"CD6D",
			x"0000" when x"CD6E",
			x"0000" when x"CD6F",
			x"0000" when x"CD70",
			x"0000" when x"CD71",
			x"0000" when x"CD72",
			x"0000" when x"CD73",
			x"0000" when x"CD74",
			x"0000" when x"CD75",
			x"0000" when x"CD76",
			x"0000" when x"CD77",
			x"0000" when x"CD78",
			x"0000" when x"CD79",
			x"0000" when x"CD7A",
			x"0000" when x"CD7B",
			x"0000" when x"CD7C",
			x"0000" when x"CD7D",
			x"0000" when x"CD7E",
			x"0000" when x"CD7F",
			x"0000" when x"CD80",
			x"0000" when x"CD81",
			x"0000" when x"CD82",
			x"0000" when x"CD83",
			x"0000" when x"CD84",
			x"0000" when x"CD85",
			x"0000" when x"CD86",
			x"0000" when x"CD87",
			x"0000" when x"CD88",
			x"0000" when x"CD89",
			x"0000" when x"CD8A",
			x"0000" when x"CD8B",
			x"0000" when x"CD8C",
			x"0000" when x"CD8D",
			x"0000" when x"CD8E",
			x"0000" when x"CD8F",
			x"0000" when x"CD90",
			x"0000" when x"CD91",
			x"0000" when x"CD92",
			x"0000" when x"CD93",
			x"0000" when x"CD94",
			x"0000" when x"CD95",
			x"0000" when x"CD96",
			x"0000" when x"CD97",
			x"0000" when x"CD98",
			x"0000" when x"CD99",
			x"0000" when x"CD9A",
			x"0000" when x"CD9B",
			x"0000" when x"CD9C",
			x"0000" when x"CD9D",
			x"0000" when x"CD9E",
			x"0000" when x"CD9F",
			x"0000" when x"CDA0",
			x"0000" when x"CDA1",
			x"0000" when x"CDA2",
			x"0000" when x"CDA3",
			x"0000" when x"CDA4",
			x"0000" when x"CDA5",
			x"0000" when x"CDA6",
			x"0000" when x"CDA7",
			x"0000" when x"CDA8",
			x"0000" when x"CDA9",
			x"0000" when x"CDAA",
			x"0000" when x"CDAB",
			x"0000" when x"CDAC",
			x"0000" when x"CDAD",
			x"0000" when x"CDAE",
			x"0000" when x"CDAF",
			x"0000" when x"CDB0",
			x"0000" when x"CDB1",
			x"0000" when x"CDB2",
			x"0000" when x"CDB3",
			x"0000" when x"CDB4",
			x"0000" when x"CDB5",
			x"0000" when x"CDB6",
			x"0000" when x"CDB7",
			x"0000" when x"CDB8",
			x"0000" when x"CDB9",
			x"0000" when x"CDBA",
			x"0000" when x"CDBB",
			x"0000" when x"CDBC",
			x"0000" when x"CDBD",
			x"0000" when x"CDBE",
			x"0000" when x"CDBF",
			x"0000" when x"CDC0",
			x"0000" when x"CDC1",
			x"0000" when x"CDC2",
			x"0000" when x"CDC3",
			x"0000" when x"CDC4",
			x"0000" when x"CDC5",
			x"0000" when x"CDC6",
			x"0000" when x"CDC7",
			x"0000" when x"CDC8",
			x"0000" when x"CDC9",
			x"0000" when x"CDCA",
			x"0000" when x"CDCB",
			x"0000" when x"CDCC",
			x"0000" when x"CDCD",
			x"0000" when x"CDCE",
			x"0000" when x"CDCF",
			x"0000" when x"CDD0",
			x"0000" when x"CDD1",
			x"0000" when x"CDD2",
			x"0000" when x"CDD3",
			x"0000" when x"CDD4",
			x"0000" when x"CDD5",
			x"0000" when x"CDD6",
			x"0000" when x"CDD7",
			x"0000" when x"CDD8",
			x"0000" when x"CDD9",
			x"0000" when x"CDDA",
			x"0000" when x"CDDB",
			x"0000" when x"CDDC",
			x"0000" when x"CDDD",
			x"0000" when x"CDDE",
			x"0000" when x"CDDF",
			x"0000" when x"CDE0",
			x"0000" when x"CDE1",
			x"0000" when x"CDE2",
			x"0000" when x"CDE3",
			x"0000" when x"CDE4",
			x"0000" when x"CDE5",
			x"0000" when x"CDE6",
			x"0000" when x"CDE7",
			x"0000" when x"CDE8",
			x"0000" when x"CDE9",
			x"0000" when x"CDEA",
			x"0000" when x"CDEB",
			x"0000" when x"CDEC",
			x"0000" when x"CDED",
			x"0000" when x"CDEE",
			x"0000" when x"CDEF",
			x"0000" when x"CDF0",
			x"0000" when x"CDF1",
			x"0000" when x"CDF2",
			x"0000" when x"CDF3",
			x"0000" when x"CDF4",
			x"0000" when x"CDF5",
			x"0000" when x"CDF6",
			x"0000" when x"CDF7",
			x"0000" when x"CDF8",
			x"0000" when x"CDF9",
			x"0000" when x"CDFA",
			x"0000" when x"CDFB",
			x"0000" when x"CDFC",
			x"0000" when x"CDFD",
			x"0000" when x"CDFE",
			x"0000" when x"CDFF",
			x"0000" when x"CE00",
			x"0000" when x"CE01",
			x"0000" when x"CE02",
			x"0000" when x"CE03",
			x"0000" when x"CE04",
			x"0000" when x"CE05",
			x"0000" when x"CE06",
			x"0000" when x"CE07",
			x"0000" when x"CE08",
			x"0000" when x"CE09",
			x"0000" when x"CE0A",
			x"0000" when x"CE0B",
			x"0000" when x"CE0C",
			x"0000" when x"CE0D",
			x"0000" when x"CE0E",
			x"0000" when x"CE0F",
			x"0000" when x"CE10",
			x"0000" when x"CE11",
			x"0000" when x"CE12",
			x"0000" when x"CE13",
			x"0000" when x"CE14",
			x"0000" when x"CE15",
			x"0000" when x"CE16",
			x"0000" when x"CE17",
			x"0000" when x"CE18",
			x"0000" when x"CE19",
			x"0000" when x"CE1A",
			x"0000" when x"CE1B",
			x"0000" when x"CE1C",
			x"0000" when x"CE1D",
			x"0000" when x"CE1E",
			x"0000" when x"CE1F",
			x"0000" when x"CE20",
			x"0000" when x"CE21",
			x"0000" when x"CE22",
			x"0000" when x"CE23",
			x"0000" when x"CE24",
			x"0000" when x"CE25",
			x"0000" when x"CE26",
			x"0000" when x"CE27",
			x"0000" when x"CE28",
			x"0000" when x"CE29",
			x"0000" when x"CE2A",
			x"0000" when x"CE2B",
			x"0000" when x"CE2C",
			x"0000" when x"CE2D",
			x"0000" when x"CE2E",
			x"0000" when x"CE2F",
			x"0000" when x"CE30",
			x"0000" when x"CE31",
			x"0000" when x"CE32",
			x"0000" when x"CE33",
			x"0000" when x"CE34",
			x"0000" when x"CE35",
			x"0000" when x"CE36",
			x"0000" when x"CE37",
			x"0000" when x"CE38",
			x"0000" when x"CE39",
			x"0000" when x"CE3A",
			x"0000" when x"CE3B",
			x"0000" when x"CE3C",
			x"0000" when x"CE3D",
			x"0000" when x"CE3E",
			x"0000" when x"CE3F",
			x"0000" when x"CE40",
			x"0000" when x"CE41",
			x"0000" when x"CE42",
			x"0000" when x"CE43",
			x"0000" when x"CE44",
			x"0000" when x"CE45",
			x"0000" when x"CE46",
			x"0000" when x"CE47",
			x"0000" when x"CE48",
			x"0000" when x"CE49",
			x"0000" when x"CE4A",
			x"0000" when x"CE4B",
			x"0000" when x"CE4C",
			x"0000" when x"CE4D",
			x"0000" when x"CE4E",
			x"0000" when x"CE4F",
			x"0000" when x"CE50",
			x"0000" when x"CE51",
			x"0000" when x"CE52",
			x"0000" when x"CE53",
			x"0000" when x"CE54",
			x"0000" when x"CE55",
			x"0000" when x"CE56",
			x"0000" when x"CE57",
			x"0000" when x"CE58",
			x"0000" when x"CE59",
			x"0000" when x"CE5A",
			x"0000" when x"CE5B",
			x"0000" when x"CE5C",
			x"0000" when x"CE5D",
			x"0000" when x"CE5E",
			x"0000" when x"CE5F",
			x"0000" when x"CE60",
			x"0000" when x"CE61",
			x"0000" when x"CE62",
			x"0000" when x"CE63",
			x"0000" when x"CE64",
			x"0000" when x"CE65",
			x"0000" when x"CE66",
			x"0000" when x"CE67",
			x"0000" when x"CE68",
			x"0000" when x"CE69",
			x"0000" when x"CE6A",
			x"0000" when x"CE6B",
			x"0000" when x"CE6C",
			x"0000" when x"CE6D",
			x"0000" when x"CE6E",
			x"0000" when x"CE6F",
			x"0000" when x"CE70",
			x"0000" when x"CE71",
			x"0000" when x"CE72",
			x"0000" when x"CE73",
			x"0000" when x"CE74",
			x"0000" when x"CE75",
			x"0000" when x"CE76",
			x"0000" when x"CE77",
			x"0000" when x"CE78",
			x"0000" when x"CE79",
			x"0000" when x"CE7A",
			x"0000" when x"CE7B",
			x"0000" when x"CE7C",
			x"0000" when x"CE7D",
			x"0000" when x"CE7E",
			x"0000" when x"CE7F",
			x"0000" when x"CE80",
			x"0000" when x"CE81",
			x"0000" when x"CE82",
			x"0000" when x"CE83",
			x"0000" when x"CE84",
			x"0000" when x"CE85",
			x"0000" when x"CE86",
			x"0000" when x"CE87",
			x"0000" when x"CE88",
			x"0000" when x"CE89",
			x"0000" when x"CE8A",
			x"0000" when x"CE8B",
			x"0000" when x"CE8C",
			x"0000" when x"CE8D",
			x"0000" when x"CE8E",
			x"0000" when x"CE8F",
			x"0000" when x"CE90",
			x"0000" when x"CE91",
			x"0000" when x"CE92",
			x"0000" when x"CE93",
			x"0000" when x"CE94",
			x"0000" when x"CE95",
			x"0000" when x"CE96",
			x"0000" when x"CE97",
			x"0000" when x"CE98",
			x"0000" when x"CE99",
			x"0000" when x"CE9A",
			x"0000" when x"CE9B",
			x"0000" when x"CE9C",
			x"0000" when x"CE9D",
			x"0000" when x"CE9E",
			x"0000" when x"CE9F",
			x"0000" when x"CEA0",
			x"0000" when x"CEA1",
			x"0000" when x"CEA2",
			x"0000" when x"CEA3",
			x"0000" when x"CEA4",
			x"0000" when x"CEA5",
			x"0000" when x"CEA6",
			x"0000" when x"CEA7",
			x"0000" when x"CEA8",
			x"0000" when x"CEA9",
			x"0000" when x"CEAA",
			x"0000" when x"CEAB",
			x"0000" when x"CEAC",
			x"0000" when x"CEAD",
			x"0000" when x"CEAE",
			x"0000" when x"CEAF",
			x"0000" when x"CEB0",
			x"0000" when x"CEB1",
			x"0000" when x"CEB2",
			x"0000" when x"CEB3",
			x"0000" when x"CEB4",
			x"0000" when x"CEB5",
			x"0000" when x"CEB6",
			x"0000" when x"CEB7",
			x"0000" when x"CEB8",
			x"0000" when x"CEB9",
			x"0000" when x"CEBA",
			x"0000" when x"CEBB",
			x"0000" when x"CEBC",
			x"0000" when x"CEBD",
			x"0000" when x"CEBE",
			x"0000" when x"CEBF",
			x"0000" when x"CEC0",
			x"0000" when x"CEC1",
			x"0000" when x"CEC2",
			x"0000" when x"CEC3",
			x"0000" when x"CEC4",
			x"0000" when x"CEC5",
			x"0000" when x"CEC6",
			x"0000" when x"CEC7",
			x"0000" when x"CEC8",
			x"0000" when x"CEC9",
			x"0000" when x"CECA",
			x"0000" when x"CECB",
			x"0000" when x"CECC",
			x"0000" when x"CECD",
			x"0000" when x"CECE",
			x"0000" when x"CECF",
			x"0000" when x"CED0",
			x"0000" when x"CED1",
			x"0000" when x"CED2",
			x"0000" when x"CED3",
			x"0000" when x"CED4",
			x"0000" when x"CED5",
			x"0000" when x"CED6",
			x"0000" when x"CED7",
			x"0000" when x"CED8",
			x"0000" when x"CED9",
			x"0000" when x"CEDA",
			x"0000" when x"CEDB",
			x"0000" when x"CEDC",
			x"0000" when x"CEDD",
			x"0000" when x"CEDE",
			x"0000" when x"CEDF",
			x"0000" when x"CEE0",
			x"0000" when x"CEE1",
			x"0000" when x"CEE2",
			x"0000" when x"CEE3",
			x"0000" when x"CEE4",
			x"0000" when x"CEE5",
			x"0000" when x"CEE6",
			x"0000" when x"CEE7",
			x"0000" when x"CEE8",
			x"0000" when x"CEE9",
			x"0000" when x"CEEA",
			x"0000" when x"CEEB",
			x"0000" when x"CEEC",
			x"0000" when x"CEED",
			x"0000" when x"CEEE",
			x"0000" when x"CEEF",
			x"0000" when x"CEF0",
			x"0000" when x"CEF1",
			x"0000" when x"CEF2",
			x"0000" when x"CEF3",
			x"0000" when x"CEF4",
			x"0000" when x"CEF5",
			x"0000" when x"CEF6",
			x"0000" when x"CEF7",
			x"0000" when x"CEF8",
			x"0000" when x"CEF9",
			x"0000" when x"CEFA",
			x"0000" when x"CEFB",
			x"0000" when x"CEFC",
			x"0000" when x"CEFD",
			x"0000" when x"CEFE",
			x"0000" when x"CEFF",
			x"0000" when x"CF00",
			x"0000" when x"CF01",
			x"0000" when x"CF02",
			x"0000" when x"CF03",
			x"0000" when x"CF04",
			x"0000" when x"CF05",
			x"0000" when x"CF06",
			x"0000" when x"CF07",
			x"0000" when x"CF08",
			x"0000" when x"CF09",
			x"0000" when x"CF0A",
			x"0000" when x"CF0B",
			x"0000" when x"CF0C",
			x"0000" when x"CF0D",
			x"0000" when x"CF0E",
			x"0000" when x"CF0F",
			x"0000" when x"CF10",
			x"0000" when x"CF11",
			x"0000" when x"CF12",
			x"0000" when x"CF13",
			x"0000" when x"CF14",
			x"0000" when x"CF15",
			x"0000" when x"CF16",
			x"0000" when x"CF17",
			x"0000" when x"CF18",
			x"0000" when x"CF19",
			x"0000" when x"CF1A",
			x"0000" when x"CF1B",
			x"0000" when x"CF1C",
			x"0000" when x"CF1D",
			x"0000" when x"CF1E",
			x"0000" when x"CF1F",
			x"0000" when x"CF20",
			x"0000" when x"CF21",
			x"0000" when x"CF22",
			x"0000" when x"CF23",
			x"0000" when x"CF24",
			x"0000" when x"CF25",
			x"0000" when x"CF26",
			x"0000" when x"CF27",
			x"0000" when x"CF28",
			x"0000" when x"CF29",
			x"0000" when x"CF2A",
			x"0000" when x"CF2B",
			x"0000" when x"CF2C",
			x"0000" when x"CF2D",
			x"0000" when x"CF2E",
			x"0000" when x"CF2F",
			x"0000" when x"CF30",
			x"0000" when x"CF31",
			x"0000" when x"CF32",
			x"0000" when x"CF33",
			x"0000" when x"CF34",
			x"0000" when x"CF35",
			x"0000" when x"CF36",
			x"0000" when x"CF37",
			x"0000" when x"CF38",
			x"0000" when x"CF39",
			x"0000" when x"CF3A",
			x"0000" when x"CF3B",
			x"0000" when x"CF3C",
			x"0000" when x"CF3D",
			x"0000" when x"CF3E",
			x"0000" when x"CF3F",
			x"0000" when x"CF40",
			x"0000" when x"CF41",
			x"0000" when x"CF42",
			x"0000" when x"CF43",
			x"0000" when x"CF44",
			x"0000" when x"CF45",
			x"0000" when x"CF46",
			x"0000" when x"CF47",
			x"0000" when x"CF48",
			x"0000" when x"CF49",
			x"0000" when x"CF4A",
			x"0000" when x"CF4B",
			x"0000" when x"CF4C",
			x"0000" when x"CF4D",
			x"0000" when x"CF4E",
			x"0000" when x"CF4F",
			x"0000" when x"CF50",
			x"0000" when x"CF51",
			x"0000" when x"CF52",
			x"0000" when x"CF53",
			x"0000" when x"CF54",
			x"0000" when x"CF55",
			x"0000" when x"CF56",
			x"0000" when x"CF57",
			x"0000" when x"CF58",
			x"0000" when x"CF59",
			x"0000" when x"CF5A",
			x"0000" when x"CF5B",
			x"0000" when x"CF5C",
			x"0000" when x"CF5D",
			x"0000" when x"CF5E",
			x"0000" when x"CF5F",
			x"0000" when x"CF60",
			x"0000" when x"CF61",
			x"0000" when x"CF62",
			x"0000" when x"CF63",
			x"0000" when x"CF64",
			x"0000" when x"CF65",
			x"0000" when x"CF66",
			x"0000" when x"CF67",
			x"0000" when x"CF68",
			x"0000" when x"CF69",
			x"0000" when x"CF6A",
			x"0000" when x"CF6B",
			x"0000" when x"CF6C",
			x"0000" when x"CF6D",
			x"0000" when x"CF6E",
			x"0000" when x"CF6F",
			x"0000" when x"CF70",
			x"0000" when x"CF71",
			x"0000" when x"CF72",
			x"0000" when x"CF73",
			x"0000" when x"CF74",
			x"0000" when x"CF75",
			x"0000" when x"CF76",
			x"0000" when x"CF77",
			x"0000" when x"CF78",
			x"0000" when x"CF79",
			x"0000" when x"CF7A",
			x"0000" when x"CF7B",
			x"0000" when x"CF7C",
			x"0000" when x"CF7D",
			x"0000" when x"CF7E",
			x"0000" when x"CF7F",
			x"0000" when x"CF80",
			x"0000" when x"CF81",
			x"0000" when x"CF82",
			x"0000" when x"CF83",
			x"0000" when x"CF84",
			x"0000" when x"CF85",
			x"0000" when x"CF86",
			x"0000" when x"CF87",
			x"0000" when x"CF88",
			x"0000" when x"CF89",
			x"0000" when x"CF8A",
			x"0000" when x"CF8B",
			x"0000" when x"CF8C",
			x"0000" when x"CF8D",
			x"0000" when x"CF8E",
			x"0000" when x"CF8F",
			x"0000" when x"CF90",
			x"0000" when x"CF91",
			x"0000" when x"CF92",
			x"0000" when x"CF93",
			x"0000" when x"CF94",
			x"0000" when x"CF95",
			x"0000" when x"CF96",
			x"0000" when x"CF97",
			x"0000" when x"CF98",
			x"0000" when x"CF99",
			x"0000" when x"CF9A",
			x"0000" when x"CF9B",
			x"0000" when x"CF9C",
			x"0000" when x"CF9D",
			x"0000" when x"CF9E",
			x"0000" when x"CF9F",
			x"0000" when x"CFA0",
			x"0000" when x"CFA1",
			x"0000" when x"CFA2",
			x"0000" when x"CFA3",
			x"0000" when x"CFA4",
			x"0000" when x"CFA5",
			x"0000" when x"CFA6",
			x"0000" when x"CFA7",
			x"0000" when x"CFA8",
			x"0000" when x"CFA9",
			x"0000" when x"CFAA",
			x"0000" when x"CFAB",
			x"0000" when x"CFAC",
			x"0000" when x"CFAD",
			x"0000" when x"CFAE",
			x"0000" when x"CFAF",
			x"0000" when x"CFB0",
			x"0000" when x"CFB1",
			x"0000" when x"CFB2",
			x"0000" when x"CFB3",
			x"0000" when x"CFB4",
			x"0000" when x"CFB5",
			x"0000" when x"CFB6",
			x"0000" when x"CFB7",
			x"0000" when x"CFB8",
			x"0000" when x"CFB9",
			x"0000" when x"CFBA",
			x"0000" when x"CFBB",
			x"0000" when x"CFBC",
			x"0000" when x"CFBD",
			x"0000" when x"CFBE",
			x"0000" when x"CFBF",
			x"0000" when x"CFC0",
			x"0000" when x"CFC1",
			x"0000" when x"CFC2",
			x"0000" when x"CFC3",
			x"0000" when x"CFC4",
			x"0000" when x"CFC5",
			x"0000" when x"CFC6",
			x"0000" when x"CFC7",
			x"0000" when x"CFC8",
			x"0000" when x"CFC9",
			x"0000" when x"CFCA",
			x"0000" when x"CFCB",
			x"0000" when x"CFCC",
			x"0000" when x"CFCD",
			x"0000" when x"CFCE",
			x"0000" when x"CFCF",
			x"0000" when x"CFD0",
			x"0000" when x"CFD1",
			x"0000" when x"CFD2",
			x"0000" when x"CFD3",
			x"0000" when x"CFD4",
			x"0000" when x"CFD5",
			x"0000" when x"CFD6",
			x"0000" when x"CFD7",
			x"0000" when x"CFD8",
			x"0000" when x"CFD9",
			x"0000" when x"CFDA",
			x"0000" when x"CFDB",
			x"0000" when x"CFDC",
			x"0000" when x"CFDD",
			x"0000" when x"CFDE",
			x"0000" when x"CFDF",
			x"0000" when x"CFE0",
			x"0000" when x"CFE1",
			x"0000" when x"CFE2",
			x"0000" when x"CFE3",
			x"0000" when x"CFE4",
			x"0000" when x"CFE5",
			x"0000" when x"CFE6",
			x"0000" when x"CFE7",
			x"0000" when x"CFE8",
			x"0000" when x"CFE9",
			x"0000" when x"CFEA",
			x"0000" when x"CFEB",
			x"0000" when x"CFEC",
			x"0000" when x"CFED",
			x"0000" when x"CFEE",
			x"0000" when x"CFEF",
			x"0000" when x"CFF0",
			x"0000" when x"CFF1",
			x"0000" when x"CFF2",
			x"0000" when x"CFF3",
			x"0000" when x"CFF4",
			x"0000" when x"CFF5",
			x"0000" when x"CFF6",
			x"0000" when x"CFF7",
			x"0000" when x"CFF8",
			x"0000" when x"CFF9",
			x"0000" when x"CFFA",
			x"0000" when x"CFFB",
			x"0000" when x"CFFC",
			x"0000" when x"CFFD",
			x"0000" when x"CFFE",
			x"0000" when x"CFFF",
			x"0000" when x"D000",
			x"0000" when x"D001",
			x"0000" when x"D002",
			x"0000" when x"D003",
			x"0000" when x"D004",
			x"0000" when x"D005",
			x"0000" when x"D006",
			x"0000" when x"D007",
			x"0000" when x"D008",
			x"0000" when x"D009",
			x"0000" when x"D00A",
			x"0000" when x"D00B",
			x"0000" when x"D00C",
			x"0000" when x"D00D",
			x"0000" when x"D00E",
			x"0000" when x"D00F",
			x"0000" when x"D010",
			x"0000" when x"D011",
			x"0000" when x"D012",
			x"0000" when x"D013",
			x"0000" when x"D014",
			x"0000" when x"D015",
			x"0000" when x"D016",
			x"0000" when x"D017",
			x"0000" when x"D018",
			x"0000" when x"D019",
			x"0000" when x"D01A",
			x"0000" when x"D01B",
			x"0000" when x"D01C",
			x"0000" when x"D01D",
			x"0000" when x"D01E",
			x"0000" when x"D01F",
			x"0000" when x"D020",
			x"0000" when x"D021",
			x"0000" when x"D022",
			x"0000" when x"D023",
			x"0000" when x"D024",
			x"0000" when x"D025",
			x"0000" when x"D026",
			x"0000" when x"D027",
			x"0000" when x"D028",
			x"0000" when x"D029",
			x"0000" when x"D02A",
			x"0000" when x"D02B",
			x"0000" when x"D02C",
			x"0000" when x"D02D",
			x"0000" when x"D02E",
			x"0000" when x"D02F",
			x"0000" when x"D030",
			x"0000" when x"D031",
			x"0000" when x"D032",
			x"0000" when x"D033",
			x"0000" when x"D034",
			x"0000" when x"D035",
			x"0000" when x"D036",
			x"0000" when x"D037",
			x"0000" when x"D038",
			x"0000" when x"D039",
			x"0000" when x"D03A",
			x"0000" when x"D03B",
			x"0000" when x"D03C",
			x"0000" when x"D03D",
			x"0000" when x"D03E",
			x"0000" when x"D03F",
			x"0000" when x"D040",
			x"0000" when x"D041",
			x"0000" when x"D042",
			x"0000" when x"D043",
			x"0000" when x"D044",
			x"0000" when x"D045",
			x"0000" when x"D046",
			x"0000" when x"D047",
			x"0000" when x"D048",
			x"0000" when x"D049",
			x"0000" when x"D04A",
			x"0000" when x"D04B",
			x"0000" when x"D04C",
			x"0000" when x"D04D",
			x"0000" when x"D04E",
			x"0000" when x"D04F",
			x"0000" when x"D050",
			x"0000" when x"D051",
			x"0000" when x"D052",
			x"0000" when x"D053",
			x"0000" when x"D054",
			x"0000" when x"D055",
			x"0000" when x"D056",
			x"0000" when x"D057",
			x"0000" when x"D058",
			x"0000" when x"D059",
			x"0000" when x"D05A",
			x"0000" when x"D05B",
			x"0000" when x"D05C",
			x"0000" when x"D05D",
			x"0000" when x"D05E",
			x"0000" when x"D05F",
			x"0000" when x"D060",
			x"0000" when x"D061",
			x"0000" when x"D062",
			x"0000" when x"D063",
			x"0000" when x"D064",
			x"0000" when x"D065",
			x"0000" when x"D066",
			x"0000" when x"D067",
			x"0000" when x"D068",
			x"0000" when x"D069",
			x"0000" when x"D06A",
			x"0000" when x"D06B",
			x"0000" when x"D06C",
			x"0000" when x"D06D",
			x"0000" when x"D06E",
			x"0000" when x"D06F",
			x"0000" when x"D070",
			x"0000" when x"D071",
			x"0000" when x"D072",
			x"0000" when x"D073",
			x"0000" when x"D074",
			x"0000" when x"D075",
			x"0000" when x"D076",
			x"0000" when x"D077",
			x"0000" when x"D078",
			x"0000" when x"D079",
			x"0000" when x"D07A",
			x"0000" when x"D07B",
			x"0000" when x"D07C",
			x"0000" when x"D07D",
			x"0000" when x"D07E",
			x"0000" when x"D07F",
			x"0000" when x"D080",
			x"0000" when x"D081",
			x"0000" when x"D082",
			x"0000" when x"D083",
			x"0000" when x"D084",
			x"0000" when x"D085",
			x"0000" when x"D086",
			x"0000" when x"D087",
			x"0000" when x"D088",
			x"0000" when x"D089",
			x"0000" when x"D08A",
			x"0000" when x"D08B",
			x"0000" when x"D08C",
			x"0000" when x"D08D",
			x"0000" when x"D08E",
			x"0000" when x"D08F",
			x"0000" when x"D090",
			x"0000" when x"D091",
			x"0000" when x"D092",
			x"0000" when x"D093",
			x"0000" when x"D094",
			x"0000" when x"D095",
			x"0000" when x"D096",
			x"0000" when x"D097",
			x"0000" when x"D098",
			x"0000" when x"D099",
			x"0000" when x"D09A",
			x"0000" when x"D09B",
			x"0000" when x"D09C",
			x"0000" when x"D09D",
			x"0000" when x"D09E",
			x"0000" when x"D09F",
			x"0000" when x"D0A0",
			x"0000" when x"D0A1",
			x"0000" when x"D0A2",
			x"0000" when x"D0A3",
			x"0000" when x"D0A4",
			x"0000" when x"D0A5",
			x"0000" when x"D0A6",
			x"0000" when x"D0A7",
			x"0000" when x"D0A8",
			x"0000" when x"D0A9",
			x"0000" when x"D0AA",
			x"0000" when x"D0AB",
			x"0000" when x"D0AC",
			x"0000" when x"D0AD",
			x"0000" when x"D0AE",
			x"0000" when x"D0AF",
			x"0000" when x"D0B0",
			x"0000" when x"D0B1",
			x"0000" when x"D0B2",
			x"0000" when x"D0B3",
			x"0000" when x"D0B4",
			x"0000" when x"D0B5",
			x"0000" when x"D0B6",
			x"0000" when x"D0B7",
			x"0000" when x"D0B8",
			x"0000" when x"D0B9",
			x"0000" when x"D0BA",
			x"0000" when x"D0BB",
			x"0000" when x"D0BC",
			x"0000" when x"D0BD",
			x"0000" when x"D0BE",
			x"0000" when x"D0BF",
			x"0000" when x"D0C0",
			x"0000" when x"D0C1",
			x"0000" when x"D0C2",
			x"0000" when x"D0C3",
			x"0000" when x"D0C4",
			x"0000" when x"D0C5",
			x"0000" when x"D0C6",
			x"0000" when x"D0C7",
			x"0000" when x"D0C8",
			x"0000" when x"D0C9",
			x"0000" when x"D0CA",
			x"0000" when x"D0CB",
			x"0000" when x"D0CC",
			x"0000" when x"D0CD",
			x"0000" when x"D0CE",
			x"0000" when x"D0CF",
			x"0000" when x"D0D0",
			x"0000" when x"D0D1",
			x"0000" when x"D0D2",
			x"0000" when x"D0D3",
			x"0000" when x"D0D4",
			x"0000" when x"D0D5",
			x"0000" when x"D0D6",
			x"0000" when x"D0D7",
			x"0000" when x"D0D8",
			x"0000" when x"D0D9",
			x"0000" when x"D0DA",
			x"0000" when x"D0DB",
			x"0000" when x"D0DC",
			x"0000" when x"D0DD",
			x"0000" when x"D0DE",
			x"0000" when x"D0DF",
			x"0000" when x"D0E0",
			x"0000" when x"D0E1",
			x"0000" when x"D0E2",
			x"0000" when x"D0E3",
			x"0000" when x"D0E4",
			x"0000" when x"D0E5",
			x"0000" when x"D0E6",
			x"0000" when x"D0E7",
			x"0000" when x"D0E8",
			x"0000" when x"D0E9",
			x"0000" when x"D0EA",
			x"0000" when x"D0EB",
			x"0000" when x"D0EC",
			x"0000" when x"D0ED",
			x"0000" when x"D0EE",
			x"0000" when x"D0EF",
			x"0000" when x"D0F0",
			x"0000" when x"D0F1",
			x"0000" when x"D0F2",
			x"0000" when x"D0F3",
			x"0000" when x"D0F4",
			x"0000" when x"D0F5",
			x"0000" when x"D0F6",
			x"0000" when x"D0F7",
			x"0000" when x"D0F8",
			x"0000" when x"D0F9",
			x"0000" when x"D0FA",
			x"0000" when x"D0FB",
			x"0000" when x"D0FC",
			x"0000" when x"D0FD",
			x"0000" when x"D0FE",
			x"0000" when x"D0FF",
			x"0000" when x"D100",
			x"0000" when x"D101",
			x"0000" when x"D102",
			x"0000" when x"D103",
			x"0000" when x"D104",
			x"0000" when x"D105",
			x"0000" when x"D106",
			x"0000" when x"D107",
			x"0000" when x"D108",
			x"0000" when x"D109",
			x"0000" when x"D10A",
			x"0000" when x"D10B",
			x"0000" when x"D10C",
			x"0000" when x"D10D",
			x"0000" when x"D10E",
			x"0000" when x"D10F",
			x"0000" when x"D110",
			x"0000" when x"D111",
			x"0000" when x"D112",
			x"0000" when x"D113",
			x"0000" when x"D114",
			x"0000" when x"D115",
			x"0000" when x"D116",
			x"0000" when x"D117",
			x"0000" when x"D118",
			x"0000" when x"D119",
			x"0000" when x"D11A",
			x"0000" when x"D11B",
			x"0000" when x"D11C",
			x"0000" when x"D11D",
			x"0000" when x"D11E",
			x"0000" when x"D11F",
			x"0000" when x"D120",
			x"0000" when x"D121",
			x"0000" when x"D122",
			x"0000" when x"D123",
			x"0000" when x"D124",
			x"0000" when x"D125",
			x"0000" when x"D126",
			x"0000" when x"D127",
			x"0000" when x"D128",
			x"0000" when x"D129",
			x"0000" when x"D12A",
			x"0000" when x"D12B",
			x"0000" when x"D12C",
			x"0000" when x"D12D",
			x"0000" when x"D12E",
			x"0000" when x"D12F",
			x"0000" when x"D130",
			x"0000" when x"D131",
			x"0000" when x"D132",
			x"0000" when x"D133",
			x"0000" when x"D134",
			x"0000" when x"D135",
			x"0000" when x"D136",
			x"0000" when x"D137",
			x"0000" when x"D138",
			x"0000" when x"D139",
			x"0000" when x"D13A",
			x"0000" when x"D13B",
			x"0000" when x"D13C",
			x"0000" when x"D13D",
			x"0000" when x"D13E",
			x"0000" when x"D13F",
			x"0000" when x"D140",
			x"0000" when x"D141",
			x"0000" when x"D142",
			x"0000" when x"D143",
			x"0000" when x"D144",
			x"0000" when x"D145",
			x"0000" when x"D146",
			x"0000" when x"D147",
			x"0000" when x"D148",
			x"0000" when x"D149",
			x"0000" when x"D14A",
			x"0000" when x"D14B",
			x"0000" when x"D14C",
			x"0000" when x"D14D",
			x"0000" when x"D14E",
			x"0000" when x"D14F",
			x"0000" when x"D150",
			x"0000" when x"D151",
			x"0000" when x"D152",
			x"0000" when x"D153",
			x"0000" when x"D154",
			x"0000" when x"D155",
			x"0000" when x"D156",
			x"0000" when x"D157",
			x"0000" when x"D158",
			x"0000" when x"D159",
			x"0000" when x"D15A",
			x"0000" when x"D15B",
			x"0000" when x"D15C",
			x"0000" when x"D15D",
			x"0000" when x"D15E",
			x"0000" when x"D15F",
			x"0000" when x"D160",
			x"0000" when x"D161",
			x"0000" when x"D162",
			x"0000" when x"D163",
			x"0000" when x"D164",
			x"0000" when x"D165",
			x"0000" when x"D166",
			x"0000" when x"D167",
			x"0000" when x"D168",
			x"0000" when x"D169",
			x"0000" when x"D16A",
			x"0000" when x"D16B",
			x"0000" when x"D16C",
			x"0000" when x"D16D",
			x"0000" when x"D16E",
			x"0000" when x"D16F",
			x"0000" when x"D170",
			x"0000" when x"D171",
			x"0000" when x"D172",
			x"0000" when x"D173",
			x"0000" when x"D174",
			x"0000" when x"D175",
			x"0000" when x"D176",
			x"0000" when x"D177",
			x"0000" when x"D178",
			x"0000" when x"D179",
			x"0000" when x"D17A",
			x"0000" when x"D17B",
			x"0000" when x"D17C",
			x"0000" when x"D17D",
			x"0000" when x"D17E",
			x"0000" when x"D17F",
			x"0000" when x"D180",
			x"0000" when x"D181",
			x"0000" when x"D182",
			x"0000" when x"D183",
			x"0000" when x"D184",
			x"0000" when x"D185",
			x"0000" when x"D186",
			x"0000" when x"D187",
			x"0000" when x"D188",
			x"0000" when x"D189",
			x"0000" when x"D18A",
			x"0000" when x"D18B",
			x"0000" when x"D18C",
			x"0000" when x"D18D",
			x"0000" when x"D18E",
			x"0000" when x"D18F",
			x"0000" when x"D190",
			x"0000" when x"D191",
			x"0000" when x"D192",
			x"0000" when x"D193",
			x"0000" when x"D194",
			x"0000" when x"D195",
			x"0000" when x"D196",
			x"0000" when x"D197",
			x"0000" when x"D198",
			x"0000" when x"D199",
			x"0000" when x"D19A",
			x"0000" when x"D19B",
			x"0000" when x"D19C",
			x"0000" when x"D19D",
			x"0000" when x"D19E",
			x"0000" when x"D19F",
			x"0000" when x"D1A0",
			x"0000" when x"D1A1",
			x"0000" when x"D1A2",
			x"0000" when x"D1A3",
			x"0000" when x"D1A4",
			x"0000" when x"D1A5",
			x"0000" when x"D1A6",
			x"0000" when x"D1A7",
			x"0000" when x"D1A8",
			x"0000" when x"D1A9",
			x"0000" when x"D1AA",
			x"0000" when x"D1AB",
			x"0000" when x"D1AC",
			x"0000" when x"D1AD",
			x"0000" when x"D1AE",
			x"0000" when x"D1AF",
			x"0000" when x"D1B0",
			x"0000" when x"D1B1",
			x"0000" when x"D1B2",
			x"0000" when x"D1B3",
			x"0000" when x"D1B4",
			x"0000" when x"D1B5",
			x"0000" when x"D1B6",
			x"0000" when x"D1B7",
			x"0000" when x"D1B8",
			x"0000" when x"D1B9",
			x"0000" when x"D1BA",
			x"0000" when x"D1BB",
			x"0000" when x"D1BC",
			x"0000" when x"D1BD",
			x"0000" when x"D1BE",
			x"0000" when x"D1BF",
			x"0000" when x"D1C0",
			x"0000" when x"D1C1",
			x"0000" when x"D1C2",
			x"0000" when x"D1C3",
			x"0000" when x"D1C4",
			x"0000" when x"D1C5",
			x"0000" when x"D1C6",
			x"0000" when x"D1C7",
			x"0000" when x"D1C8",
			x"0000" when x"D1C9",
			x"0000" when x"D1CA",
			x"0000" when x"D1CB",
			x"0000" when x"D1CC",
			x"0000" when x"D1CD",
			x"0000" when x"D1CE",
			x"0000" when x"D1CF",
			x"0000" when x"D1D0",
			x"0000" when x"D1D1",
			x"0000" when x"D1D2",
			x"0000" when x"D1D3",
			x"0000" when x"D1D4",
			x"0000" when x"D1D5",
			x"0000" when x"D1D6",
			x"0000" when x"D1D7",
			x"0000" when x"D1D8",
			x"0000" when x"D1D9",
			x"0000" when x"D1DA",
			x"0000" when x"D1DB",
			x"0000" when x"D1DC",
			x"0000" when x"D1DD",
			x"0000" when x"D1DE",
			x"0000" when x"D1DF",
			x"0000" when x"D1E0",
			x"0000" when x"D1E1",
			x"0000" when x"D1E2",
			x"0000" when x"D1E3",
			x"0000" when x"D1E4",
			x"0000" when x"D1E5",
			x"0000" when x"D1E6",
			x"0000" when x"D1E7",
			x"0000" when x"D1E8",
			x"0000" when x"D1E9",
			x"0000" when x"D1EA",
			x"0000" when x"D1EB",
			x"0000" when x"D1EC",
			x"0000" when x"D1ED",
			x"0000" when x"D1EE",
			x"0000" when x"D1EF",
			x"0000" when x"D1F0",
			x"0000" when x"D1F1",
			x"0000" when x"D1F2",
			x"0000" when x"D1F3",
			x"0000" when x"D1F4",
			x"0000" when x"D1F5",
			x"0000" when x"D1F6",
			x"0000" when x"D1F7",
			x"0000" when x"D1F8",
			x"0000" when x"D1F9",
			x"0000" when x"D1FA",
			x"0000" when x"D1FB",
			x"0000" when x"D1FC",
			x"0000" when x"D1FD",
			x"0000" when x"D1FE",
			x"0000" when x"D1FF",
			x"0000" when x"D200",
			x"0000" when x"D201",
			x"0000" when x"D202",
			x"0000" when x"D203",
			x"0000" when x"D204",
			x"0000" when x"D205",
			x"0000" when x"D206",
			x"0000" when x"D207",
			x"0000" when x"D208",
			x"0000" when x"D209",
			x"0000" when x"D20A",
			x"0000" when x"D20B",
			x"0000" when x"D20C",
			x"0000" when x"D20D",
			x"0000" when x"D20E",
			x"0000" when x"D20F",
			x"0000" when x"D210",
			x"0000" when x"D211",
			x"0000" when x"D212",
			x"0000" when x"D213",
			x"0000" when x"D214",
			x"0000" when x"D215",
			x"0000" when x"D216",
			x"0000" when x"D217",
			x"0000" when x"D218",
			x"0000" when x"D219",
			x"0000" when x"D21A",
			x"0000" when x"D21B",
			x"0000" when x"D21C",
			x"0000" when x"D21D",
			x"0000" when x"D21E",
			x"0000" when x"D21F",
			x"0000" when x"D220",
			x"0000" when x"D221",
			x"0000" when x"D222",
			x"0000" when x"D223",
			x"0000" when x"D224",
			x"0000" when x"D225",
			x"0000" when x"D226",
			x"0000" when x"D227",
			x"0000" when x"D228",
			x"0000" when x"D229",
			x"0000" when x"D22A",
			x"0000" when x"D22B",
			x"0000" when x"D22C",
			x"0000" when x"D22D",
			x"0000" when x"D22E",
			x"0000" when x"D22F",
			x"0000" when x"D230",
			x"0000" when x"D231",
			x"0000" when x"D232",
			x"0000" when x"D233",
			x"0000" when x"D234",
			x"0000" when x"D235",
			x"0000" when x"D236",
			x"0000" when x"D237",
			x"0000" when x"D238",
			x"0000" when x"D239",
			x"0000" when x"D23A",
			x"0000" when x"D23B",
			x"0000" when x"D23C",
			x"0000" when x"D23D",
			x"0000" when x"D23E",
			x"0000" when x"D23F",
			x"0000" when x"D240",
			x"0000" when x"D241",
			x"0000" when x"D242",
			x"0000" when x"D243",
			x"0000" when x"D244",
			x"0000" when x"D245",
			x"0000" when x"D246",
			x"0000" when x"D247",
			x"0000" when x"D248",
			x"0000" when x"D249",
			x"0000" when x"D24A",
			x"0000" when x"D24B",
			x"0000" when x"D24C",
			x"0000" when x"D24D",
			x"0000" when x"D24E",
			x"0000" when x"D24F",
			x"0000" when x"D250",
			x"0000" when x"D251",
			x"0000" when x"D252",
			x"0000" when x"D253",
			x"0000" when x"D254",
			x"0000" when x"D255",
			x"0000" when x"D256",
			x"0000" when x"D257",
			x"0000" when x"D258",
			x"0000" when x"D259",
			x"0000" when x"D25A",
			x"0000" when x"D25B",
			x"0000" when x"D25C",
			x"0000" when x"D25D",
			x"0000" when x"D25E",
			x"0000" when x"D25F",
			x"0000" when x"D260",
			x"0000" when x"D261",
			x"0000" when x"D262",
			x"0000" when x"D263",
			x"0000" when x"D264",
			x"0000" when x"D265",
			x"0000" when x"D266",
			x"0000" when x"D267",
			x"0000" when x"D268",
			x"0000" when x"D269",
			x"0000" when x"D26A",
			x"0000" when x"D26B",
			x"0000" when x"D26C",
			x"0000" when x"D26D",
			x"0000" when x"D26E",
			x"0000" when x"D26F",
			x"0000" when x"D270",
			x"0000" when x"D271",
			x"0000" when x"D272",
			x"0000" when x"D273",
			x"0000" when x"D274",
			x"0000" when x"D275",
			x"0000" when x"D276",
			x"0000" when x"D277",
			x"0000" when x"D278",
			x"0000" when x"D279",
			x"0000" when x"D27A",
			x"0000" when x"D27B",
			x"0000" when x"D27C",
			x"0000" when x"D27D",
			x"0000" when x"D27E",
			x"0000" when x"D27F",
			x"0000" when x"D280",
			x"0000" when x"D281",
			x"0000" when x"D282",
			x"0000" when x"D283",
			x"0000" when x"D284",
			x"0000" when x"D285",
			x"0000" when x"D286",
			x"0000" when x"D287",
			x"0000" when x"D288",
			x"0000" when x"D289",
			x"0000" when x"D28A",
			x"0000" when x"D28B",
			x"0000" when x"D28C",
			x"0000" when x"D28D",
			x"0000" when x"D28E",
			x"0000" when x"D28F",
			x"0000" when x"D290",
			x"0000" when x"D291",
			x"0000" when x"D292",
			x"0000" when x"D293",
			x"0000" when x"D294",
			x"0000" when x"D295",
			x"0000" when x"D296",
			x"0000" when x"D297",
			x"0000" when x"D298",
			x"0000" when x"D299",
			x"0000" when x"D29A",
			x"0000" when x"D29B",
			x"0000" when x"D29C",
			x"0000" when x"D29D",
			x"0000" when x"D29E",
			x"0000" when x"D29F",
			x"0000" when x"D2A0",
			x"0000" when x"D2A1",
			x"0000" when x"D2A2",
			x"0000" when x"D2A3",
			x"0000" when x"D2A4",
			x"0000" when x"D2A5",
			x"0000" when x"D2A6",
			x"0000" when x"D2A7",
			x"0000" when x"D2A8",
			x"0000" when x"D2A9",
			x"0000" when x"D2AA",
			x"0000" when x"D2AB",
			x"0000" when x"D2AC",
			x"0000" when x"D2AD",
			x"0000" when x"D2AE",
			x"0000" when x"D2AF",
			x"0000" when x"D2B0",
			x"0000" when x"D2B1",
			x"0000" when x"D2B2",
			x"0000" when x"D2B3",
			x"0000" when x"D2B4",
			x"0000" when x"D2B5",
			x"0000" when x"D2B6",
			x"0000" when x"D2B7",
			x"0000" when x"D2B8",
			x"0000" when x"D2B9",
			x"0000" when x"D2BA",
			x"0000" when x"D2BB",
			x"0000" when x"D2BC",
			x"0000" when x"D2BD",
			x"0000" when x"D2BE",
			x"0000" when x"D2BF",
			x"0000" when x"D2C0",
			x"0000" when x"D2C1",
			x"0000" when x"D2C2",
			x"0000" when x"D2C3",
			x"0000" when x"D2C4",
			x"0000" when x"D2C5",
			x"0000" when x"D2C6",
			x"0000" when x"D2C7",
			x"0000" when x"D2C8",
			x"0000" when x"D2C9",
			x"0000" when x"D2CA",
			x"0000" when x"D2CB",
			x"0000" when x"D2CC",
			x"0000" when x"D2CD",
			x"0000" when x"D2CE",
			x"0000" when x"D2CF",
			x"0000" when x"D2D0",
			x"0000" when x"D2D1",
			x"0000" when x"D2D2",
			x"0000" when x"D2D3",
			x"0000" when x"D2D4",
			x"0000" when x"D2D5",
			x"0000" when x"D2D6",
			x"0000" when x"D2D7",
			x"0000" when x"D2D8",
			x"0000" when x"D2D9",
			x"0000" when x"D2DA",
			x"0000" when x"D2DB",
			x"0000" when x"D2DC",
			x"0000" when x"D2DD",
			x"0000" when x"D2DE",
			x"0000" when x"D2DF",
			x"0000" when x"D2E0",
			x"0000" when x"D2E1",
			x"0000" when x"D2E2",
			x"0000" when x"D2E3",
			x"0000" when x"D2E4",
			x"0000" when x"D2E5",
			x"0000" when x"D2E6",
			x"0000" when x"D2E7",
			x"0000" when x"D2E8",
			x"0000" when x"D2E9",
			x"0000" when x"D2EA",
			x"0000" when x"D2EB",
			x"0000" when x"D2EC",
			x"0000" when x"D2ED",
			x"0000" when x"D2EE",
			x"0000" when x"D2EF",
			x"0000" when x"D2F0",
			x"0000" when x"D2F1",
			x"0000" when x"D2F2",
			x"0000" when x"D2F3",
			x"0000" when x"D2F4",
			x"0000" when x"D2F5",
			x"0000" when x"D2F6",
			x"0000" when x"D2F7",
			x"0000" when x"D2F8",
			x"0000" when x"D2F9",
			x"0000" when x"D2FA",
			x"0000" when x"D2FB",
			x"0000" when x"D2FC",
			x"0000" when x"D2FD",
			x"0000" when x"D2FE",
			x"0000" when x"D2FF",
			x"0000" when x"D300",
			x"0000" when x"D301",
			x"0000" when x"D302",
			x"0000" when x"D303",
			x"0000" when x"D304",
			x"0000" when x"D305",
			x"0000" when x"D306",
			x"0000" when x"D307",
			x"0000" when x"D308",
			x"0000" when x"D309",
			x"0000" when x"D30A",
			x"0000" when x"D30B",
			x"0000" when x"D30C",
			x"0000" when x"D30D",
			x"0000" when x"D30E",
			x"0000" when x"D30F",
			x"0000" when x"D310",
			x"0000" when x"D311",
			x"0000" when x"D312",
			x"0000" when x"D313",
			x"0000" when x"D314",
			x"0000" when x"D315",
			x"0000" when x"D316",
			x"0000" when x"D317",
			x"0000" when x"D318",
			x"0000" when x"D319",
			x"0000" when x"D31A",
			x"0000" when x"D31B",
			x"0000" when x"D31C",
			x"0000" when x"D31D",
			x"0000" when x"D31E",
			x"0000" when x"D31F",
			x"0000" when x"D320",
			x"0000" when x"D321",
			x"0000" when x"D322",
			x"0000" when x"D323",
			x"0000" when x"D324",
			x"0000" when x"D325",
			x"0000" when x"D326",
			x"0000" when x"D327",
			x"0000" when x"D328",
			x"0000" when x"D329",
			x"0000" when x"D32A",
			x"0000" when x"D32B",
			x"0000" when x"D32C",
			x"0000" when x"D32D",
			x"0000" when x"D32E",
			x"0000" when x"D32F",
			x"0000" when x"D330",
			x"0000" when x"D331",
			x"0000" when x"D332",
			x"0000" when x"D333",
			x"0000" when x"D334",
			x"0000" when x"D335",
			x"0000" when x"D336",
			x"0000" when x"D337",
			x"0000" when x"D338",
			x"0000" when x"D339",
			x"0000" when x"D33A",
			x"0000" when x"D33B",
			x"0000" when x"D33C",
			x"0000" when x"D33D",
			x"0000" when x"D33E",
			x"0000" when x"D33F",
			x"0000" when x"D340",
			x"0000" when x"D341",
			x"0000" when x"D342",
			x"0000" when x"D343",
			x"0000" when x"D344",
			x"0000" when x"D345",
			x"0000" when x"D346",
			x"0000" when x"D347",
			x"0000" when x"D348",
			x"0000" when x"D349",
			x"0000" when x"D34A",
			x"0000" when x"D34B",
			x"0000" when x"D34C",
			x"0000" when x"D34D",
			x"0000" when x"D34E",
			x"0000" when x"D34F",
			x"0000" when x"D350",
			x"0000" when x"D351",
			x"0000" when x"D352",
			x"0000" when x"D353",
			x"0000" when x"D354",
			x"0000" when x"D355",
			x"0000" when x"D356",
			x"0000" when x"D357",
			x"0000" when x"D358",
			x"0000" when x"D359",
			x"0000" when x"D35A",
			x"0000" when x"D35B",
			x"0000" when x"D35C",
			x"0000" when x"D35D",
			x"0000" when x"D35E",
			x"0000" when x"D35F",
			x"0000" when x"D360",
			x"0000" when x"D361",
			x"0000" when x"D362",
			x"0000" when x"D363",
			x"0000" when x"D364",
			x"0000" when x"D365",
			x"0000" when x"D366",
			x"0000" when x"D367",
			x"0000" when x"D368",
			x"0000" when x"D369",
			x"0000" when x"D36A",
			x"0000" when x"D36B",
			x"0000" when x"D36C",
			x"0000" when x"D36D",
			x"0000" when x"D36E",
			x"0000" when x"D36F",
			x"0000" when x"D370",
			x"0000" when x"D371",
			x"0000" when x"D372",
			x"0000" when x"D373",
			x"0000" when x"D374",
			x"0000" when x"D375",
			x"0000" when x"D376",
			x"0000" when x"D377",
			x"0000" when x"D378",
			x"0000" when x"D379",
			x"0000" when x"D37A",
			x"0000" when x"D37B",
			x"0000" when x"D37C",
			x"0000" when x"D37D",
			x"0000" when x"D37E",
			x"0000" when x"D37F",
			x"0000" when x"D380",
			x"0000" when x"D381",
			x"0000" when x"D382",
			x"0000" when x"D383",
			x"0000" when x"D384",
			x"0000" when x"D385",
			x"0000" when x"D386",
			x"0000" when x"D387",
			x"0000" when x"D388",
			x"0000" when x"D389",
			x"0000" when x"D38A",
			x"0000" when x"D38B",
			x"0000" when x"D38C",
			x"0000" when x"D38D",
			x"0000" when x"D38E",
			x"0000" when x"D38F",
			x"0000" when x"D390",
			x"0000" when x"D391",
			x"0000" when x"D392",
			x"0000" when x"D393",
			x"0000" when x"D394",
			x"0000" when x"D395",
			x"0000" when x"D396",
			x"0000" when x"D397",
			x"0000" when x"D398",
			x"0000" when x"D399",
			x"0000" when x"D39A",
			x"0000" when x"D39B",
			x"0000" when x"D39C",
			x"0000" when x"D39D",
			x"0000" when x"D39E",
			x"0000" when x"D39F",
			x"0000" when x"D3A0",
			x"0000" when x"D3A1",
			x"0000" when x"D3A2",
			x"0000" when x"D3A3",
			x"0000" when x"D3A4",
			x"0000" when x"D3A5",
			x"0000" when x"D3A6",
			x"0000" when x"D3A7",
			x"0000" when x"D3A8",
			x"0000" when x"D3A9",
			x"0000" when x"D3AA",
			x"0000" when x"D3AB",
			x"0000" when x"D3AC",
			x"0000" when x"D3AD",
			x"0000" when x"D3AE",
			x"0000" when x"D3AF",
			x"0000" when x"D3B0",
			x"0000" when x"D3B1",
			x"0000" when x"D3B2",
			x"0000" when x"D3B3",
			x"0000" when x"D3B4",
			x"0000" when x"D3B5",
			x"0000" when x"D3B6",
			x"0000" when x"D3B7",
			x"0000" when x"D3B8",
			x"0000" when x"D3B9",
			x"0000" when x"D3BA",
			x"0000" when x"D3BB",
			x"0000" when x"D3BC",
			x"0000" when x"D3BD",
			x"0000" when x"D3BE",
			x"0000" when x"D3BF",
			x"0000" when x"D3C0",
			x"0000" when x"D3C1",
			x"0000" when x"D3C2",
			x"0000" when x"D3C3",
			x"0000" when x"D3C4",
			x"0000" when x"D3C5",
			x"0000" when x"D3C6",
			x"0000" when x"D3C7",
			x"0000" when x"D3C8",
			x"0000" when x"D3C9",
			x"0000" when x"D3CA",
			x"0000" when x"D3CB",
			x"0000" when x"D3CC",
			x"0000" when x"D3CD",
			x"0000" when x"D3CE",
			x"0000" when x"D3CF",
			x"0000" when x"D3D0",
			x"0000" when x"D3D1",
			x"0000" when x"D3D2",
			x"0000" when x"D3D3",
			x"0000" when x"D3D4",
			x"0000" when x"D3D5",
			x"0000" when x"D3D6",
			x"0000" when x"D3D7",
			x"0000" when x"D3D8",
			x"0000" when x"D3D9",
			x"0000" when x"D3DA",
			x"0000" when x"D3DB",
			x"0000" when x"D3DC",
			x"0000" when x"D3DD",
			x"0000" when x"D3DE",
			x"0000" when x"D3DF",
			x"0000" when x"D3E0",
			x"0000" when x"D3E1",
			x"0000" when x"D3E2",
			x"0000" when x"D3E3",
			x"0000" when x"D3E4",
			x"0000" when x"D3E5",
			x"0000" when x"D3E6",
			x"0000" when x"D3E7",
			x"0000" when x"D3E8",
			x"0000" when x"D3E9",
			x"0000" when x"D3EA",
			x"0000" when x"D3EB",
			x"0000" when x"D3EC",
			x"0000" when x"D3ED",
			x"0000" when x"D3EE",
			x"0000" when x"D3EF",
			x"0000" when x"D3F0",
			x"0000" when x"D3F1",
			x"0000" when x"D3F2",
			x"0000" when x"D3F3",
			x"0000" when x"D3F4",
			x"0000" when x"D3F5",
			x"0000" when x"D3F6",
			x"0000" when x"D3F7",
			x"0000" when x"D3F8",
			x"0000" when x"D3F9",
			x"0000" when x"D3FA",
			x"0000" when x"D3FB",
			x"0000" when x"D3FC",
			x"0000" when x"D3FD",
			x"0000" when x"D3FE",
			x"0000" when x"D3FF",
			x"0000" when x"D400",
			x"0000" when x"D401",
			x"0000" when x"D402",
			x"0000" when x"D403",
			x"0000" when x"D404",
			x"0000" when x"D405",
			x"0000" when x"D406",
			x"0000" when x"D407",
			x"0000" when x"D408",
			x"0000" when x"D409",
			x"0000" when x"D40A",
			x"0000" when x"D40B",
			x"0000" when x"D40C",
			x"0000" when x"D40D",
			x"0000" when x"D40E",
			x"0000" when x"D40F",
			x"0000" when x"D410",
			x"0000" when x"D411",
			x"0000" when x"D412",
			x"0000" when x"D413",
			x"0000" when x"D414",
			x"0000" when x"D415",
			x"0000" when x"D416",
			x"0000" when x"D417",
			x"0000" when x"D418",
			x"0000" when x"D419",
			x"0000" when x"D41A",
			x"0000" when x"D41B",
			x"0000" when x"D41C",
			x"0000" when x"D41D",
			x"0000" when x"D41E",
			x"0000" when x"D41F",
			x"0000" when x"D420",
			x"0000" when x"D421",
			x"0000" when x"D422",
			x"0000" when x"D423",
			x"0000" when x"D424",
			x"0000" when x"D425",
			x"0000" when x"D426",
			x"0000" when x"D427",
			x"0000" when x"D428",
			x"0000" when x"D429",
			x"0000" when x"D42A",
			x"0000" when x"D42B",
			x"0000" when x"D42C",
			x"0000" when x"D42D",
			x"0000" when x"D42E",
			x"0000" when x"D42F",
			x"0000" when x"D430",
			x"0000" when x"D431",
			x"0000" when x"D432",
			x"0000" when x"D433",
			x"0000" when x"D434",
			x"0000" when x"D435",
			x"0000" when x"D436",
			x"0000" when x"D437",
			x"0000" when x"D438",
			x"0000" when x"D439",
			x"0000" when x"D43A",
			x"0000" when x"D43B",
			x"0000" when x"D43C",
			x"0000" when x"D43D",
			x"0000" when x"D43E",
			x"0000" when x"D43F",
			x"0000" when x"D440",
			x"0000" when x"D441",
			x"0000" when x"D442",
			x"0000" when x"D443",
			x"0000" when x"D444",
			x"0000" when x"D445",
			x"0000" when x"D446",
			x"0000" when x"D447",
			x"0000" when x"D448",
			x"0000" when x"D449",
			x"0000" when x"D44A",
			x"0000" when x"D44B",
			x"0000" when x"D44C",
			x"0000" when x"D44D",
			x"0000" when x"D44E",
			x"0000" when x"D44F",
			x"0000" when x"D450",
			x"0000" when x"D451",
			x"0000" when x"D452",
			x"0000" when x"D453",
			x"0000" when x"D454",
			x"0000" when x"D455",
			x"0000" when x"D456",
			x"0000" when x"D457",
			x"0000" when x"D458",
			x"0000" when x"D459",
			x"0000" when x"D45A",
			x"0000" when x"D45B",
			x"0000" when x"D45C",
			x"0000" when x"D45D",
			x"0000" when x"D45E",
			x"0000" when x"D45F",
			x"0000" when x"D460",
			x"0000" when x"D461",
			x"0000" when x"D462",
			x"0000" when x"D463",
			x"0000" when x"D464",
			x"0000" when x"D465",
			x"0000" when x"D466",
			x"0000" when x"D467",
			x"0000" when x"D468",
			x"0000" when x"D469",
			x"0000" when x"D46A",
			x"0000" when x"D46B",
			x"0000" when x"D46C",
			x"0000" when x"D46D",
			x"0000" when x"D46E",
			x"0000" when x"D46F",
			x"0000" when x"D470",
			x"0000" when x"D471",
			x"0000" when x"D472",
			x"0000" when x"D473",
			x"0000" when x"D474",
			x"0000" when x"D475",
			x"0000" when x"D476",
			x"0000" when x"D477",
			x"0000" when x"D478",
			x"0000" when x"D479",
			x"0000" when x"D47A",
			x"0000" when x"D47B",
			x"0000" when x"D47C",
			x"0000" when x"D47D",
			x"0000" when x"D47E",
			x"0000" when x"D47F",
			x"0000" when x"D480",
			x"0000" when x"D481",
			x"0000" when x"D482",
			x"0000" when x"D483",
			x"0000" when x"D484",
			x"0000" when x"D485",
			x"0000" when x"D486",
			x"0000" when x"D487",
			x"0000" when x"D488",
			x"0000" when x"D489",
			x"0000" when x"D48A",
			x"0000" when x"D48B",
			x"0000" when x"D48C",
			x"0000" when x"D48D",
			x"0000" when x"D48E",
			x"0000" when x"D48F",
			x"0000" when x"D490",
			x"0000" when x"D491",
			x"0000" when x"D492",
			x"0000" when x"D493",
			x"0000" when x"D494",
			x"0000" when x"D495",
			x"0000" when x"D496",
			x"0000" when x"D497",
			x"0000" when x"D498",
			x"0000" when x"D499",
			x"0000" when x"D49A",
			x"0000" when x"D49B",
			x"0000" when x"D49C",
			x"0000" when x"D49D",
			x"0000" when x"D49E",
			x"0000" when x"D49F",
			x"0000" when x"D4A0",
			x"0000" when x"D4A1",
			x"0000" when x"D4A2",
			x"0000" when x"D4A3",
			x"0000" when x"D4A4",
			x"0000" when x"D4A5",
			x"0000" when x"D4A6",
			x"0000" when x"D4A7",
			x"0000" when x"D4A8",
			x"0000" when x"D4A9",
			x"0000" when x"D4AA",
			x"0000" when x"D4AB",
			x"0000" when x"D4AC",
			x"0000" when x"D4AD",
			x"0000" when x"D4AE",
			x"0000" when x"D4AF",
			x"0000" when x"D4B0",
			x"0000" when x"D4B1",
			x"0000" when x"D4B2",
			x"0000" when x"D4B3",
			x"0000" when x"D4B4",
			x"0000" when x"D4B5",
			x"0000" when x"D4B6",
			x"0000" when x"D4B7",
			x"0000" when x"D4B8",
			x"0000" when x"D4B9",
			x"0000" when x"D4BA",
			x"0000" when x"D4BB",
			x"0000" when x"D4BC",
			x"0000" when x"D4BD",
			x"0000" when x"D4BE",
			x"0000" when x"D4BF",
			x"0000" when x"D4C0",
			x"0000" when x"D4C1",
			x"0000" when x"D4C2",
			x"0000" when x"D4C3",
			x"0000" when x"D4C4",
			x"0000" when x"D4C5",
			x"0000" when x"D4C6",
			x"0000" when x"D4C7",
			x"0000" when x"D4C8",
			x"0000" when x"D4C9",
			x"0000" when x"D4CA",
			x"0000" when x"D4CB",
			x"0000" when x"D4CC",
			x"0000" when x"D4CD",
			x"0000" when x"D4CE",
			x"0000" when x"D4CF",
			x"0000" when x"D4D0",
			x"0000" when x"D4D1",
			x"0000" when x"D4D2",
			x"0000" when x"D4D3",
			x"0000" when x"D4D4",
			x"0000" when x"D4D5",
			x"0000" when x"D4D6",
			x"0000" when x"D4D7",
			x"0000" when x"D4D8",
			x"0000" when x"D4D9",
			x"0000" when x"D4DA",
			x"0000" when x"D4DB",
			x"0000" when x"D4DC",
			x"0000" when x"D4DD",
			x"0000" when x"D4DE",
			x"0000" when x"D4DF",
			x"0000" when x"D4E0",
			x"0000" when x"D4E1",
			x"0000" when x"D4E2",
			x"0000" when x"D4E3",
			x"0000" when x"D4E4",
			x"0000" when x"D4E5",
			x"0000" when x"D4E6",
			x"0000" when x"D4E7",
			x"0000" when x"D4E8",
			x"0000" when x"D4E9",
			x"0000" when x"D4EA",
			x"0000" when x"D4EB",
			x"0000" when x"D4EC",
			x"0000" when x"D4ED",
			x"0000" when x"D4EE",
			x"0000" when x"D4EF",
			x"0000" when x"D4F0",
			x"0000" when x"D4F1",
			x"0000" when x"D4F2",
			x"0000" when x"D4F3",
			x"0000" when x"D4F4",
			x"0000" when x"D4F5",
			x"0000" when x"D4F6",
			x"0000" when x"D4F7",
			x"0000" when x"D4F8",
			x"0000" when x"D4F9",
			x"0000" when x"D4FA",
			x"0000" when x"D4FB",
			x"0000" when x"D4FC",
			x"0000" when x"D4FD",
			x"0000" when x"D4FE",
			x"0000" when x"D4FF",
			x"0000" when x"D500",
			x"0000" when x"D501",
			x"0000" when x"D502",
			x"0000" when x"D503",
			x"0000" when x"D504",
			x"0000" when x"D505",
			x"0000" when x"D506",
			x"0000" when x"D507",
			x"0000" when x"D508",
			x"0000" when x"D509",
			x"0000" when x"D50A",
			x"0000" when x"D50B",
			x"0000" when x"D50C",
			x"0000" when x"D50D",
			x"0000" when x"D50E",
			x"0000" when x"D50F",
			x"0000" when x"D510",
			x"0000" when x"D511",
			x"0000" when x"D512",
			x"0000" when x"D513",
			x"0000" when x"D514",
			x"0000" when x"D515",
			x"0000" when x"D516",
			x"0000" when x"D517",
			x"0000" when x"D518",
			x"0000" when x"D519",
			x"0000" when x"D51A",
			x"0000" when x"D51B",
			x"0000" when x"D51C",
			x"0000" when x"D51D",
			x"0000" when x"D51E",
			x"0000" when x"D51F",
			x"0000" when x"D520",
			x"0000" when x"D521",
			x"0000" when x"D522",
			x"0000" when x"D523",
			x"0000" when x"D524",
			x"0000" when x"D525",
			x"0000" when x"D526",
			x"0000" when x"D527",
			x"0000" when x"D528",
			x"0000" when x"D529",
			x"0000" when x"D52A",
			x"0000" when x"D52B",
			x"0000" when x"D52C",
			x"0000" when x"D52D",
			x"0000" when x"D52E",
			x"0000" when x"D52F",
			x"0000" when x"D530",
			x"0000" when x"D531",
			x"0000" when x"D532",
			x"0000" when x"D533",
			x"0000" when x"D534",
			x"0000" when x"D535",
			x"0000" when x"D536",
			x"0000" when x"D537",
			x"0000" when x"D538",
			x"0000" when x"D539",
			x"0000" when x"D53A",
			x"0000" when x"D53B",
			x"0000" when x"D53C",
			x"0000" when x"D53D",
			x"0000" when x"D53E",
			x"0000" when x"D53F",
			x"0000" when x"D540",
			x"0000" when x"D541",
			x"0000" when x"D542",
			x"0000" when x"D543",
			x"0000" when x"D544",
			x"0000" when x"D545",
			x"0000" when x"D546",
			x"0000" when x"D547",
			x"0000" when x"D548",
			x"0000" when x"D549",
			x"0000" when x"D54A",
			x"0000" when x"D54B",
			x"0000" when x"D54C",
			x"0000" when x"D54D",
			x"0000" when x"D54E",
			x"0000" when x"D54F",
			x"0000" when x"D550",
			x"0000" when x"D551",
			x"0000" when x"D552",
			x"0000" when x"D553",
			x"0000" when x"D554",
			x"0000" when x"D555",
			x"0000" when x"D556",
			x"0000" when x"D557",
			x"0000" when x"D558",
			x"0000" when x"D559",
			x"0000" when x"D55A",
			x"0000" when x"D55B",
			x"0000" when x"D55C",
			x"0000" when x"D55D",
			x"0000" when x"D55E",
			x"0000" when x"D55F",
			x"0000" when x"D560",
			x"0000" when x"D561",
			x"0000" when x"D562",
			x"0000" when x"D563",
			x"0000" when x"D564",
			x"0000" when x"D565",
			x"0000" when x"D566",
			x"0000" when x"D567",
			x"0000" when x"D568",
			x"0000" when x"D569",
			x"0000" when x"D56A",
			x"0000" when x"D56B",
			x"0000" when x"D56C",
			x"0000" when x"D56D",
			x"0000" when x"D56E",
			x"0000" when x"D56F",
			x"0000" when x"D570",
			x"0000" when x"D571",
			x"0000" when x"D572",
			x"0000" when x"D573",
			x"0000" when x"D574",
			x"0000" when x"D575",
			x"0000" when x"D576",
			x"0000" when x"D577",
			x"0000" when x"D578",
			x"0000" when x"D579",
			x"0000" when x"D57A",
			x"0000" when x"D57B",
			x"0000" when x"D57C",
			x"0000" when x"D57D",
			x"0000" when x"D57E",
			x"0000" when x"D57F",
			x"0000" when x"D580",
			x"0000" when x"D581",
			x"0000" when x"D582",
			x"0000" when x"D583",
			x"0000" when x"D584",
			x"0000" when x"D585",
			x"0000" when x"D586",
			x"0000" when x"D587",
			x"0000" when x"D588",
			x"0000" when x"D589",
			x"0000" when x"D58A",
			x"0000" when x"D58B",
			x"0000" when x"D58C",
			x"0000" when x"D58D",
			x"0000" when x"D58E",
			x"0000" when x"D58F",
			x"0000" when x"D590",
			x"0000" when x"D591",
			x"0000" when x"D592",
			x"0000" when x"D593",
			x"0000" when x"D594",
			x"0000" when x"D595",
			x"0000" when x"D596",
			x"0000" when x"D597",
			x"0000" when x"D598",
			x"0000" when x"D599",
			x"0000" when x"D59A",
			x"0000" when x"D59B",
			x"0000" when x"D59C",
			x"0000" when x"D59D",
			x"0000" when x"D59E",
			x"0000" when x"D59F",
			x"0000" when x"D5A0",
			x"0000" when x"D5A1",
			x"0000" when x"D5A2",
			x"0000" when x"D5A3",
			x"0000" when x"D5A4",
			x"0000" when x"D5A5",
			x"0000" when x"D5A6",
			x"0000" when x"D5A7",
			x"0000" when x"D5A8",
			x"0000" when x"D5A9",
			x"0000" when x"D5AA",
			x"0000" when x"D5AB",
			x"0000" when x"D5AC",
			x"0000" when x"D5AD",
			x"0000" when x"D5AE",
			x"0000" when x"D5AF",
			x"0000" when x"D5B0",
			x"0000" when x"D5B1",
			x"0000" when x"D5B2",
			x"0000" when x"D5B3",
			x"0000" when x"D5B4",
			x"0000" when x"D5B5",
			x"0000" when x"D5B6",
			x"0000" when x"D5B7",
			x"0000" when x"D5B8",
			x"0000" when x"D5B9",
			x"0000" when x"D5BA",
			x"0000" when x"D5BB",
			x"0000" when x"D5BC",
			x"0000" when x"D5BD",
			x"0000" when x"D5BE",
			x"0000" when x"D5BF",
			x"0000" when x"D5C0",
			x"0000" when x"D5C1",
			x"0000" when x"D5C2",
			x"0000" when x"D5C3",
			x"0000" when x"D5C4",
			x"0000" when x"D5C5",
			x"0000" when x"D5C6",
			x"0000" when x"D5C7",
			x"0000" when x"D5C8",
			x"0000" when x"D5C9",
			x"0000" when x"D5CA",
			x"0000" when x"D5CB",
			x"0000" when x"D5CC",
			x"0000" when x"D5CD",
			x"0000" when x"D5CE",
			x"0000" when x"D5CF",
			x"0000" when x"D5D0",
			x"0000" when x"D5D1",
			x"0000" when x"D5D2",
			x"0000" when x"D5D3",
			x"0000" when x"D5D4",
			x"0000" when x"D5D5",
			x"0000" when x"D5D6",
			x"0000" when x"D5D7",
			x"0000" when x"D5D8",
			x"0000" when x"D5D9",
			x"0000" when x"D5DA",
			x"0000" when x"D5DB",
			x"0000" when x"D5DC",
			x"0000" when x"D5DD",
			x"0000" when x"D5DE",
			x"0000" when x"D5DF",
			x"0000" when x"D5E0",
			x"0000" when x"D5E1",
			x"0000" when x"D5E2",
			x"0000" when x"D5E3",
			x"0000" when x"D5E4",
			x"0000" when x"D5E5",
			x"0000" when x"D5E6",
			x"0000" when x"D5E7",
			x"0000" when x"D5E8",
			x"0000" when x"D5E9",
			x"0000" when x"D5EA",
			x"0000" when x"D5EB",
			x"0000" when x"D5EC",
			x"0000" when x"D5ED",
			x"0000" when x"D5EE",
			x"0000" when x"D5EF",
			x"0000" when x"D5F0",
			x"0000" when x"D5F1",
			x"0000" when x"D5F2",
			x"0000" when x"D5F3",
			x"0000" when x"D5F4",
			x"0000" when x"D5F5",
			x"0000" when x"D5F6",
			x"0000" when x"D5F7",
			x"0000" when x"D5F8",
			x"0000" when x"D5F9",
			x"0000" when x"D5FA",
			x"0000" when x"D5FB",
			x"0000" when x"D5FC",
			x"0000" when x"D5FD",
			x"0000" when x"D5FE",
			x"0000" when x"D5FF",
			x"0000" when x"D600",
			x"0000" when x"D601",
			x"0000" when x"D602",
			x"0000" when x"D603",
			x"0000" when x"D604",
			x"0000" when x"D605",
			x"0000" when x"D606",
			x"0000" when x"D607",
			x"0000" when x"D608",
			x"0000" when x"D609",
			x"0000" when x"D60A",
			x"0000" when x"D60B",
			x"0000" when x"D60C",
			x"0000" when x"D60D",
			x"0000" when x"D60E",
			x"0000" when x"D60F",
			x"0000" when x"D610",
			x"0000" when x"D611",
			x"0000" when x"D612",
			x"0000" when x"D613",
			x"0000" when x"D614",
			x"0000" when x"D615",
			x"0000" when x"D616",
			x"0000" when x"D617",
			x"0000" when x"D618",
			x"0000" when x"D619",
			x"0000" when x"D61A",
			x"0000" when x"D61B",
			x"0000" when x"D61C",
			x"0000" when x"D61D",
			x"0000" when x"D61E",
			x"0000" when x"D61F",
			x"0000" when x"D620",
			x"0000" when x"D621",
			x"0000" when x"D622",
			x"0000" when x"D623",
			x"0000" when x"D624",
			x"0000" when x"D625",
			x"0000" when x"D626",
			x"0000" when x"D627",
			x"0000" when x"D628",
			x"0000" when x"D629",
			x"0000" when x"D62A",
			x"0000" when x"D62B",
			x"0000" when x"D62C",
			x"0000" when x"D62D",
			x"0000" when x"D62E",
			x"0000" when x"D62F",
			x"0000" when x"D630",
			x"0000" when x"D631",
			x"0000" when x"D632",
			x"0000" when x"D633",
			x"0000" when x"D634",
			x"0000" when x"D635",
			x"0000" when x"D636",
			x"0000" when x"D637",
			x"0000" when x"D638",
			x"0000" when x"D639",
			x"0000" when x"D63A",
			x"0000" when x"D63B",
			x"0000" when x"D63C",
			x"0000" when x"D63D",
			x"0000" when x"D63E",
			x"0000" when x"D63F",
			x"0000" when x"D640",
			x"0000" when x"D641",
			x"0000" when x"D642",
			x"0000" when x"D643",
			x"0000" when x"D644",
			x"0000" when x"D645",
			x"0000" when x"D646",
			x"0000" when x"D647",
			x"0000" when x"D648",
			x"0000" when x"D649",
			x"0000" when x"D64A",
			x"0000" when x"D64B",
			x"0000" when x"D64C",
			x"0000" when x"D64D",
			x"0000" when x"D64E",
			x"0000" when x"D64F",
			x"0000" when x"D650",
			x"0000" when x"D651",
			x"0000" when x"D652",
			x"0000" when x"D653",
			x"0000" when x"D654",
			x"0000" when x"D655",
			x"0000" when x"D656",
			x"0000" when x"D657",
			x"0000" when x"D658",
			x"0000" when x"D659",
			x"0000" when x"D65A",
			x"0000" when x"D65B",
			x"0000" when x"D65C",
			x"0000" when x"D65D",
			x"0000" when x"D65E",
			x"0000" when x"D65F",
			x"0000" when x"D660",
			x"0000" when x"D661",
			x"0000" when x"D662",
			x"0000" when x"D663",
			x"0000" when x"D664",
			x"0000" when x"D665",
			x"0000" when x"D666",
			x"0000" when x"D667",
			x"0000" when x"D668",
			x"0000" when x"D669",
			x"0000" when x"D66A",
			x"0000" when x"D66B",
			x"0000" when x"D66C",
			x"0000" when x"D66D",
			x"0000" when x"D66E",
			x"0000" when x"D66F",
			x"0000" when x"D670",
			x"0000" when x"D671",
			x"0000" when x"D672",
			x"0000" when x"D673",
			x"0000" when x"D674",
			x"0000" when x"D675",
			x"0000" when x"D676",
			x"0000" when x"D677",
			x"0000" when x"D678",
			x"0000" when x"D679",
			x"0000" when x"D67A",
			x"0000" when x"D67B",
			x"0000" when x"D67C",
			x"0000" when x"D67D",
			x"0000" when x"D67E",
			x"0000" when x"D67F",
			x"0000" when x"D680",
			x"0000" when x"D681",
			x"0000" when x"D682",
			x"0000" when x"D683",
			x"0000" when x"D684",
			x"0000" when x"D685",
			x"0000" when x"D686",
			x"0000" when x"D687",
			x"0000" when x"D688",
			x"0000" when x"D689",
			x"0000" when x"D68A",
			x"0000" when x"D68B",
			x"0000" when x"D68C",
			x"0000" when x"D68D",
			x"0000" when x"D68E",
			x"0000" when x"D68F",
			x"0000" when x"D690",
			x"0000" when x"D691",
			x"0000" when x"D692",
			x"0000" when x"D693",
			x"0000" when x"D694",
			x"0000" when x"D695",
			x"0000" when x"D696",
			x"0000" when x"D697",
			x"0000" when x"D698",
			x"0000" when x"D699",
			x"0000" when x"D69A",
			x"0000" when x"D69B",
			x"0000" when x"D69C",
			x"0000" when x"D69D",
			x"0000" when x"D69E",
			x"0000" when x"D69F",
			x"0000" when x"D6A0",
			x"0000" when x"D6A1",
			x"0000" when x"D6A2",
			x"0000" when x"D6A3",
			x"0000" when x"D6A4",
			x"0000" when x"D6A5",
			x"0000" when x"D6A6",
			x"0000" when x"D6A7",
			x"0000" when x"D6A8",
			x"0000" when x"D6A9",
			x"0000" when x"D6AA",
			x"0000" when x"D6AB",
			x"0000" when x"D6AC",
			x"0000" when x"D6AD",
			x"0000" when x"D6AE",
			x"0000" when x"D6AF",
			x"0000" when x"D6B0",
			x"0000" when x"D6B1",
			x"0000" when x"D6B2",
			x"0000" when x"D6B3",
			x"0000" when x"D6B4",
			x"0000" when x"D6B5",
			x"0000" when x"D6B6",
			x"0000" when x"D6B7",
			x"0000" when x"D6B8",
			x"0000" when x"D6B9",
			x"0000" when x"D6BA",
			x"0000" when x"D6BB",
			x"0000" when x"D6BC",
			x"0000" when x"D6BD",
			x"0000" when x"D6BE",
			x"0000" when x"D6BF",
			x"0000" when x"D6C0",
			x"0000" when x"D6C1",
			x"0000" when x"D6C2",
			x"0000" when x"D6C3",
			x"0000" when x"D6C4",
			x"0000" when x"D6C5",
			x"0000" when x"D6C6",
			x"0000" when x"D6C7",
			x"0000" when x"D6C8",
			x"0000" when x"D6C9",
			x"0000" when x"D6CA",
			x"0000" when x"D6CB",
			x"0000" when x"D6CC",
			x"0000" when x"D6CD",
			x"0000" when x"D6CE",
			x"0000" when x"D6CF",
			x"0000" when x"D6D0",
			x"0000" when x"D6D1",
			x"0000" when x"D6D2",
			x"0000" when x"D6D3",
			x"0000" when x"D6D4",
			x"0000" when x"D6D5",
			x"0000" when x"D6D6",
			x"0000" when x"D6D7",
			x"0000" when x"D6D8",
			x"0000" when x"D6D9",
			x"0000" when x"D6DA",
			x"0000" when x"D6DB",
			x"0000" when x"D6DC",
			x"0000" when x"D6DD",
			x"0000" when x"D6DE",
			x"0000" when x"D6DF",
			x"0000" when x"D6E0",
			x"0000" when x"D6E1",
			x"0000" when x"D6E2",
			x"0000" when x"D6E3",
			x"0000" when x"D6E4",
			x"0000" when x"D6E5",
			x"0000" when x"D6E6",
			x"0000" when x"D6E7",
			x"0000" when x"D6E8",
			x"0000" when x"D6E9",
			x"0000" when x"D6EA",
			x"0000" when x"D6EB",
			x"0000" when x"D6EC",
			x"0000" when x"D6ED",
			x"0000" when x"D6EE",
			x"0000" when x"D6EF",
			x"0000" when x"D6F0",
			x"0000" when x"D6F1",
			x"0000" when x"D6F2",
			x"0000" when x"D6F3",
			x"0000" when x"D6F4",
			x"0000" when x"D6F5",
			x"0000" when x"D6F6",
			x"0000" when x"D6F7",
			x"0000" when x"D6F8",
			x"0000" when x"D6F9",
			x"0000" when x"D6FA",
			x"0000" when x"D6FB",
			x"0000" when x"D6FC",
			x"0000" when x"D6FD",
			x"0000" when x"D6FE",
			x"0000" when x"D6FF",
			x"0000" when x"D700",
			x"0000" when x"D701",
			x"0000" when x"D702",
			x"0000" when x"D703",
			x"0000" when x"D704",
			x"0000" when x"D705",
			x"0000" when x"D706",
			x"0000" when x"D707",
			x"0000" when x"D708",
			x"0000" when x"D709",
			x"0000" when x"D70A",
			x"0000" when x"D70B",
			x"0000" when x"D70C",
			x"0000" when x"D70D",
			x"0000" when x"D70E",
			x"0000" when x"D70F",
			x"0000" when x"D710",
			x"0000" when x"D711",
			x"0000" when x"D712",
			x"0000" when x"D713",
			x"0000" when x"D714",
			x"0000" when x"D715",
			x"0000" when x"D716",
			x"0000" when x"D717",
			x"0000" when x"D718",
			x"0000" when x"D719",
			x"0000" when x"D71A",
			x"0000" when x"D71B",
			x"0000" when x"D71C",
			x"0000" when x"D71D",
			x"0000" when x"D71E",
			x"0000" when x"D71F",
			x"0000" when x"D720",
			x"0000" when x"D721",
			x"0000" when x"D722",
			x"0000" when x"D723",
			x"0000" when x"D724",
			x"0000" when x"D725",
			x"0000" when x"D726",
			x"0000" when x"D727",
			x"0000" when x"D728",
			x"0000" when x"D729",
			x"0000" when x"D72A",
			x"0000" when x"D72B",
			x"0000" when x"D72C",
			x"0000" when x"D72D",
			x"0000" when x"D72E",
			x"0000" when x"D72F",
			x"0000" when x"D730",
			x"0000" when x"D731",
			x"0000" when x"D732",
			x"0000" when x"D733",
			x"0000" when x"D734",
			x"0000" when x"D735",
			x"0000" when x"D736",
			x"0000" when x"D737",
			x"0000" when x"D738",
			x"0000" when x"D739",
			x"0000" when x"D73A",
			x"0000" when x"D73B",
			x"0000" when x"D73C",
			x"0000" when x"D73D",
			x"0000" when x"D73E",
			x"0000" when x"D73F",
			x"0000" when x"D740",
			x"0000" when x"D741",
			x"0000" when x"D742",
			x"0000" when x"D743",
			x"0000" when x"D744",
			x"0000" when x"D745",
			x"0000" when x"D746",
			x"0000" when x"D747",
			x"0000" when x"D748",
			x"0000" when x"D749",
			x"0000" when x"D74A",
			x"0000" when x"D74B",
			x"0000" when x"D74C",
			x"0000" when x"D74D",
			x"0000" when x"D74E",
			x"0000" when x"D74F",
			x"0000" when x"D750",
			x"0000" when x"D751",
			x"0000" when x"D752",
			x"0000" when x"D753",
			x"0000" when x"D754",
			x"0000" when x"D755",
			x"0000" when x"D756",
			x"0000" when x"D757",
			x"0000" when x"D758",
			x"0000" when x"D759",
			x"0000" when x"D75A",
			x"0000" when x"D75B",
			x"0000" when x"D75C",
			x"0000" when x"D75D",
			x"0000" when x"D75E",
			x"0000" when x"D75F",
			x"0000" when x"D760",
			x"0000" when x"D761",
			x"0000" when x"D762",
			x"0000" when x"D763",
			x"0000" when x"D764",
			x"0000" when x"D765",
			x"0000" when x"D766",
			x"0000" when x"D767",
			x"0000" when x"D768",
			x"0000" when x"D769",
			x"0000" when x"D76A",
			x"0000" when x"D76B",
			x"0000" when x"D76C",
			x"0000" when x"D76D",
			x"0000" when x"D76E",
			x"0000" when x"D76F",
			x"0000" when x"D770",
			x"0000" when x"D771",
			x"0000" when x"D772",
			x"0000" when x"D773",
			x"0000" when x"D774",
			x"0000" when x"D775",
			x"0000" when x"D776",
			x"0000" when x"D777",
			x"0000" when x"D778",
			x"0000" when x"D779",
			x"0000" when x"D77A",
			x"0000" when x"D77B",
			x"0000" when x"D77C",
			x"0000" when x"D77D",
			x"0000" when x"D77E",
			x"0000" when x"D77F",
			x"0000" when x"D780",
			x"0000" when x"D781",
			x"0000" when x"D782",
			x"0000" when x"D783",
			x"0000" when x"D784",
			x"0000" when x"D785",
			x"0000" when x"D786",
			x"0000" when x"D787",
			x"0000" when x"D788",
			x"0000" when x"D789",
			x"0000" when x"D78A",
			x"0000" when x"D78B",
			x"0000" when x"D78C",
			x"0000" when x"D78D",
			x"0000" when x"D78E",
			x"0000" when x"D78F",
			x"0000" when x"D790",
			x"0000" when x"D791",
			x"0000" when x"D792",
			x"0000" when x"D793",
			x"0000" when x"D794",
			x"0000" when x"D795",
			x"0000" when x"D796",
			x"0000" when x"D797",
			x"0000" when x"D798",
			x"0000" when x"D799",
			x"0000" when x"D79A",
			x"0000" when x"D79B",
			x"0000" when x"D79C",
			x"0000" when x"D79D",
			x"0000" when x"D79E",
			x"0000" when x"D79F",
			x"0000" when x"D7A0",
			x"0000" when x"D7A1",
			x"0000" when x"D7A2",
			x"0000" when x"D7A3",
			x"0000" when x"D7A4",
			x"0000" when x"D7A5",
			x"0000" when x"D7A6",
			x"0000" when x"D7A7",
			x"0000" when x"D7A8",
			x"0000" when x"D7A9",
			x"0000" when x"D7AA",
			x"0000" when x"D7AB",
			x"0000" when x"D7AC",
			x"0000" when x"D7AD",
			x"0000" when x"D7AE",
			x"0000" when x"D7AF",
			x"0000" when x"D7B0",
			x"0000" when x"D7B1",
			x"0000" when x"D7B2",
			x"0000" when x"D7B3",
			x"0000" when x"D7B4",
			x"0000" when x"D7B5",
			x"0000" when x"D7B6",
			x"0000" when x"D7B7",
			x"0000" when x"D7B8",
			x"0000" when x"D7B9",
			x"0000" when x"D7BA",
			x"0000" when x"D7BB",
			x"0000" when x"D7BC",
			x"0000" when x"D7BD",
			x"0000" when x"D7BE",
			x"0000" when x"D7BF",
			x"0000" when x"D7C0",
			x"0000" when x"D7C1",
			x"0000" when x"D7C2",
			x"0000" when x"D7C3",
			x"0000" when x"D7C4",
			x"0000" when x"D7C5",
			x"0000" when x"D7C6",
			x"0000" when x"D7C7",
			x"0000" when x"D7C8",
			x"0000" when x"D7C9",
			x"0000" when x"D7CA",
			x"0000" when x"D7CB",
			x"0000" when x"D7CC",
			x"0000" when x"D7CD",
			x"0000" when x"D7CE",
			x"0000" when x"D7CF",
			x"0000" when x"D7D0",
			x"0000" when x"D7D1",
			x"0000" when x"D7D2",
			x"0000" when x"D7D3",
			x"0000" when x"D7D4",
			x"0000" when x"D7D5",
			x"0000" when x"D7D6",
			x"0000" when x"D7D7",
			x"0000" when x"D7D8",
			x"0000" when x"D7D9",
			x"0000" when x"D7DA",
			x"0000" when x"D7DB",
			x"0000" when x"D7DC",
			x"0000" when x"D7DD",
			x"0000" when x"D7DE",
			x"0000" when x"D7DF",
			x"0000" when x"D7E0",
			x"0000" when x"D7E1",
			x"0000" when x"D7E2",
			x"0000" when x"D7E3",
			x"0000" when x"D7E4",
			x"0000" when x"D7E5",
			x"0000" when x"D7E6",
			x"0000" when x"D7E7",
			x"0000" when x"D7E8",
			x"0000" when x"D7E9",
			x"0000" when x"D7EA",
			x"0000" when x"D7EB",
			x"0000" when x"D7EC",
			x"0000" when x"D7ED",
			x"0000" when x"D7EE",
			x"0000" when x"D7EF",
			x"0000" when x"D7F0",
			x"0000" when x"D7F1",
			x"0000" when x"D7F2",
			x"0000" when x"D7F3",
			x"0000" when x"D7F4",
			x"0000" when x"D7F5",
			x"0000" when x"D7F6",
			x"0000" when x"D7F7",
			x"0000" when x"D7F8",
			x"0000" when x"D7F9",
			x"0000" when x"D7FA",
			x"0000" when x"D7FB",
			x"0000" when x"D7FC",
			x"0000" when x"D7FD",
			x"0000" when x"D7FE",
			x"0000" when x"D7FF",
			x"0000" when x"D800",
			x"0000" when x"D801",
			x"0000" when x"D802",
			x"0000" when x"D803",
			x"0000" when x"D804",
			x"0000" when x"D805",
			x"0000" when x"D806",
			x"0000" when x"D807",
			x"0000" when x"D808",
			x"0000" when x"D809",
			x"0000" when x"D80A",
			x"0000" when x"D80B",
			x"0000" when x"D80C",
			x"0000" when x"D80D",
			x"0000" when x"D80E",
			x"0000" when x"D80F",
			x"0000" when x"D810",
			x"0000" when x"D811",
			x"0000" when x"D812",
			x"0000" when x"D813",
			x"0000" when x"D814",
			x"0000" when x"D815",
			x"0000" when x"D816",
			x"0000" when x"D817",
			x"0000" when x"D818",
			x"0000" when x"D819",
			x"0000" when x"D81A",
			x"0000" when x"D81B",
			x"0000" when x"D81C",
			x"0000" when x"D81D",
			x"0000" when x"D81E",
			x"0000" when x"D81F",
			x"0000" when x"D820",
			x"0000" when x"D821",
			x"0000" when x"D822",
			x"0000" when x"D823",
			x"0000" when x"D824",
			x"0000" when x"D825",
			x"0000" when x"D826",
			x"0000" when x"D827",
			x"0000" when x"D828",
			x"0000" when x"D829",
			x"0000" when x"D82A",
			x"0000" when x"D82B",
			x"0000" when x"D82C",
			x"0000" when x"D82D",
			x"0000" when x"D82E",
			x"0000" when x"D82F",
			x"0000" when x"D830",
			x"0000" when x"D831",
			x"0000" when x"D832",
			x"0000" when x"D833",
			x"0000" when x"D834",
			x"0000" when x"D835",
			x"0000" when x"D836",
			x"0000" when x"D837",
			x"0000" when x"D838",
			x"0000" when x"D839",
			x"0000" when x"D83A",
			x"0000" when x"D83B",
			x"0000" when x"D83C",
			x"0000" when x"D83D",
			x"0000" when x"D83E",
			x"0000" when x"D83F",
			x"0000" when x"D840",
			x"0000" when x"D841",
			x"0000" when x"D842",
			x"0000" when x"D843",
			x"0000" when x"D844",
			x"0000" when x"D845",
			x"0000" when x"D846",
			x"0000" when x"D847",
			x"0000" when x"D848",
			x"0000" when x"D849",
			x"0000" when x"D84A",
			x"0000" when x"D84B",
			x"0000" when x"D84C",
			x"0000" when x"D84D",
			x"0000" when x"D84E",
			x"0000" when x"D84F",
			x"0000" when x"D850",
			x"0000" when x"D851",
			x"0000" when x"D852",
			x"0000" when x"D853",
			x"0000" when x"D854",
			x"0000" when x"D855",
			x"0000" when x"D856",
			x"0000" when x"D857",
			x"0000" when x"D858",
			x"0000" when x"D859",
			x"0000" when x"D85A",
			x"0000" when x"D85B",
			x"0000" when x"D85C",
			x"0000" when x"D85D",
			x"0000" when x"D85E",
			x"0000" when x"D85F",
			x"0000" when x"D860",
			x"0000" when x"D861",
			x"0000" when x"D862",
			x"0000" when x"D863",
			x"0000" when x"D864",
			x"0000" when x"D865",
			x"0000" when x"D866",
			x"0000" when x"D867",
			x"0000" when x"D868",
			x"0000" when x"D869",
			x"0000" when x"D86A",
			x"0000" when x"D86B",
			x"0000" when x"D86C",
			x"0000" when x"D86D",
			x"0000" when x"D86E",
			x"0000" when x"D86F",
			x"0000" when x"D870",
			x"0000" when x"D871",
			x"0000" when x"D872",
			x"0000" when x"D873",
			x"0000" when x"D874",
			x"0000" when x"D875",
			x"0000" when x"D876",
			x"0000" when x"D877",
			x"0000" when x"D878",
			x"0000" when x"D879",
			x"0000" when x"D87A",
			x"0000" when x"D87B",
			x"0000" when x"D87C",
			x"0000" when x"D87D",
			x"0000" when x"D87E",
			x"0000" when x"D87F",
			x"0000" when x"D880",
			x"0000" when x"D881",
			x"0000" when x"D882",
			x"0000" when x"D883",
			x"0000" when x"D884",
			x"0000" when x"D885",
			x"0000" when x"D886",
			x"0000" when x"D887",
			x"0000" when x"D888",
			x"0000" when x"D889",
			x"0000" when x"D88A",
			x"0000" when x"D88B",
			x"0000" when x"D88C",
			x"0000" when x"D88D",
			x"0000" when x"D88E",
			x"0000" when x"D88F",
			x"0000" when x"D890",
			x"0000" when x"D891",
			x"0000" when x"D892",
			x"0000" when x"D893",
			x"0000" when x"D894",
			x"0000" when x"D895",
			x"0000" when x"D896",
			x"0000" when x"D897",
			x"0000" when x"D898",
			x"0000" when x"D899",
			x"0000" when x"D89A",
			x"0000" when x"D89B",
			x"0000" when x"D89C",
			x"0000" when x"D89D",
			x"0000" when x"D89E",
			x"0000" when x"D89F",
			x"0000" when x"D8A0",
			x"0000" when x"D8A1",
			x"0000" when x"D8A2",
			x"0000" when x"D8A3",
			x"0000" when x"D8A4",
			x"0000" when x"D8A5",
			x"0000" when x"D8A6",
			x"0000" when x"D8A7",
			x"0000" when x"D8A8",
			x"0000" when x"D8A9",
			x"0000" when x"D8AA",
			x"0000" when x"D8AB",
			x"0000" when x"D8AC",
			x"0000" when x"D8AD",
			x"0000" when x"D8AE",
			x"0000" when x"D8AF",
			x"0000" when x"D8B0",
			x"0000" when x"D8B1",
			x"0000" when x"D8B2",
			x"0000" when x"D8B3",
			x"0000" when x"D8B4",
			x"0000" when x"D8B5",
			x"0000" when x"D8B6",
			x"0000" when x"D8B7",
			x"0000" when x"D8B8",
			x"0000" when x"D8B9",
			x"0000" when x"D8BA",
			x"0000" when x"D8BB",
			x"0000" when x"D8BC",
			x"0000" when x"D8BD",
			x"0000" when x"D8BE",
			x"0000" when x"D8BF",
			x"0000" when x"D8C0",
			x"0000" when x"D8C1",
			x"0000" when x"D8C2",
			x"0000" when x"D8C3",
			x"0000" when x"D8C4",
			x"0000" when x"D8C5",
			x"0000" when x"D8C6",
			x"0000" when x"D8C7",
			x"0000" when x"D8C8",
			x"0000" when x"D8C9",
			x"0000" when x"D8CA",
			x"0000" when x"D8CB",
			x"0000" when x"D8CC",
			x"0000" when x"D8CD",
			x"0000" when x"D8CE",
			x"0000" when x"D8CF",
			x"0000" when x"D8D0",
			x"0000" when x"D8D1",
			x"0000" when x"D8D2",
			x"0000" when x"D8D3",
			x"0000" when x"D8D4",
			x"0000" when x"D8D5",
			x"0000" when x"D8D6",
			x"0000" when x"D8D7",
			x"0000" when x"D8D8",
			x"0000" when x"D8D9",
			x"0000" when x"D8DA",
			x"0000" when x"D8DB",
			x"0000" when x"D8DC",
			x"0000" when x"D8DD",
			x"0000" when x"D8DE",
			x"0000" when x"D8DF",
			x"0000" when x"D8E0",
			x"0000" when x"D8E1",
			x"0000" when x"D8E2",
			x"0000" when x"D8E3",
			x"0000" when x"D8E4",
			x"0000" when x"D8E5",
			x"0000" when x"D8E6",
			x"0000" when x"D8E7",
			x"0000" when x"D8E8",
			x"0000" when x"D8E9",
			x"0000" when x"D8EA",
			x"0000" when x"D8EB",
			x"0000" when x"D8EC",
			x"0000" when x"D8ED",
			x"0000" when x"D8EE",
			x"0000" when x"D8EF",
			x"0000" when x"D8F0",
			x"0000" when x"D8F1",
			x"0000" when x"D8F2",
			x"0000" when x"D8F3",
			x"0000" when x"D8F4",
			x"0000" when x"D8F5",
			x"0000" when x"D8F6",
			x"0000" when x"D8F7",
			x"0000" when x"D8F8",
			x"0000" when x"D8F9",
			x"0000" when x"D8FA",
			x"0000" when x"D8FB",
			x"0000" when x"D8FC",
			x"0000" when x"D8FD",
			x"0000" when x"D8FE",
			x"0000" when x"D8FF",
			x"0000" when x"D900",
			x"0000" when x"D901",
			x"0000" when x"D902",
			x"0000" when x"D903",
			x"0000" when x"D904",
			x"0000" when x"D905",
			x"0000" when x"D906",
			x"0000" when x"D907",
			x"0000" when x"D908",
			x"0000" when x"D909",
			x"0000" when x"D90A",
			x"0000" when x"D90B",
			x"0000" when x"D90C",
			x"0000" when x"D90D",
			x"0000" when x"D90E",
			x"0000" when x"D90F",
			x"0000" when x"D910",
			x"0000" when x"D911",
			x"0000" when x"D912",
			x"0000" when x"D913",
			x"0000" when x"D914",
			x"0000" when x"D915",
			x"0000" when x"D916",
			x"0000" when x"D917",
			x"0000" when x"D918",
			x"0000" when x"D919",
			x"0000" when x"D91A",
			x"0000" when x"D91B",
			x"0000" when x"D91C",
			x"0000" when x"D91D",
			x"0000" when x"D91E",
			x"0000" when x"D91F",
			x"0000" when x"D920",
			x"0000" when x"D921",
			x"0000" when x"D922",
			x"0000" when x"D923",
			x"0000" when x"D924",
			x"0000" when x"D925",
			x"0000" when x"D926",
			x"0000" when x"D927",
			x"0000" when x"D928",
			x"0000" when x"D929",
			x"0000" when x"D92A",
			x"0000" when x"D92B",
			x"0000" when x"D92C",
			x"0000" when x"D92D",
			x"0000" when x"D92E",
			x"0000" when x"D92F",
			x"0000" when x"D930",
			x"0000" when x"D931",
			x"0000" when x"D932",
			x"0000" when x"D933",
			x"0000" when x"D934",
			x"0000" when x"D935",
			x"0000" when x"D936",
			x"0000" when x"D937",
			x"0000" when x"D938",
			x"0000" when x"D939",
			x"0000" when x"D93A",
			x"0000" when x"D93B",
			x"0000" when x"D93C",
			x"0000" when x"D93D",
			x"0000" when x"D93E",
			x"0000" when x"D93F",
			x"0000" when x"D940",
			x"0000" when x"D941",
			x"0000" when x"D942",
			x"0000" when x"D943",
			x"0000" when x"D944",
			x"0000" when x"D945",
			x"0000" when x"D946",
			x"0000" when x"D947",
			x"0000" when x"D948",
			x"0000" when x"D949",
			x"0000" when x"D94A",
			x"0000" when x"D94B",
			x"0000" when x"D94C",
			x"0000" when x"D94D",
			x"0000" when x"D94E",
			x"0000" when x"D94F",
			x"0000" when x"D950",
			x"0000" when x"D951",
			x"0000" when x"D952",
			x"0000" when x"D953",
			x"0000" when x"D954",
			x"0000" when x"D955",
			x"0000" when x"D956",
			x"0000" when x"D957",
			x"0000" when x"D958",
			x"0000" when x"D959",
			x"0000" when x"D95A",
			x"0000" when x"D95B",
			x"0000" when x"D95C",
			x"0000" when x"D95D",
			x"0000" when x"D95E",
			x"0000" when x"D95F",
			x"0000" when x"D960",
			x"0000" when x"D961",
			x"0000" when x"D962",
			x"0000" when x"D963",
			x"0000" when x"D964",
			x"0000" when x"D965",
			x"0000" when x"D966",
			x"0000" when x"D967",
			x"0000" when x"D968",
			x"0000" when x"D969",
			x"0000" when x"D96A",
			x"0000" when x"D96B",
			x"0000" when x"D96C",
			x"0000" when x"D96D",
			x"0000" when x"D96E",
			x"0000" when x"D96F",
			x"0000" when x"D970",
			x"0000" when x"D971",
			x"0000" when x"D972",
			x"0000" when x"D973",
			x"0000" when x"D974",
			x"0000" when x"D975",
			x"0000" when x"D976",
			x"0000" when x"D977",
			x"0000" when x"D978",
			x"0000" when x"D979",
			x"0000" when x"D97A",
			x"0000" when x"D97B",
			x"0000" when x"D97C",
			x"0000" when x"D97D",
			x"0000" when x"D97E",
			x"0000" when x"D97F",
			x"0000" when x"D980",
			x"0000" when x"D981",
			x"0000" when x"D982",
			x"0000" when x"D983",
			x"0000" when x"D984",
			x"0000" when x"D985",
			x"0000" when x"D986",
			x"0000" when x"D987",
			x"0000" when x"D988",
			x"0000" when x"D989",
			x"0000" when x"D98A",
			x"0000" when x"D98B",
			x"0000" when x"D98C",
			x"0000" when x"D98D",
			x"0000" when x"D98E",
			x"0000" when x"D98F",
			x"0000" when x"D990",
			x"0000" when x"D991",
			x"0000" when x"D992",
			x"0000" when x"D993",
			x"0000" when x"D994",
			x"0000" when x"D995",
			x"0000" when x"D996",
			x"0000" when x"D997",
			x"0000" when x"D998",
			x"0000" when x"D999",
			x"0000" when x"D99A",
			x"0000" when x"D99B",
			x"0000" when x"D99C",
			x"0000" when x"D99D",
			x"0000" when x"D99E",
			x"0000" when x"D99F",
			x"0000" when x"D9A0",
			x"0000" when x"D9A1",
			x"0000" when x"D9A2",
			x"0000" when x"D9A3",
			x"0000" when x"D9A4",
			x"0000" when x"D9A5",
			x"0000" when x"D9A6",
			x"0000" when x"D9A7",
			x"0000" when x"D9A8",
			x"0000" when x"D9A9",
			x"0000" when x"D9AA",
			x"0000" when x"D9AB",
			x"0000" when x"D9AC",
			x"0000" when x"D9AD",
			x"0000" when x"D9AE",
			x"0000" when x"D9AF",
			x"0000" when x"D9B0",
			x"0000" when x"D9B1",
			x"0000" when x"D9B2",
			x"0000" when x"D9B3",
			x"0000" when x"D9B4",
			x"0000" when x"D9B5",
			x"0000" when x"D9B6",
			x"0000" when x"D9B7",
			x"0000" when x"D9B8",
			x"0000" when x"D9B9",
			x"0000" when x"D9BA",
			x"0000" when x"D9BB",
			x"0000" when x"D9BC",
			x"0000" when x"D9BD",
			x"0000" when x"D9BE",
			x"0000" when x"D9BF",
			x"0000" when x"D9C0",
			x"0000" when x"D9C1",
			x"0000" when x"D9C2",
			x"0000" when x"D9C3",
			x"0000" when x"D9C4",
			x"0000" when x"D9C5",
			x"0000" when x"D9C6",
			x"0000" when x"D9C7",
			x"0000" when x"D9C8",
			x"0000" when x"D9C9",
			x"0000" when x"D9CA",
			x"0000" when x"D9CB",
			x"0000" when x"D9CC",
			x"0000" when x"D9CD",
			x"0000" when x"D9CE",
			x"0000" when x"D9CF",
			x"0000" when x"D9D0",
			x"0000" when x"D9D1",
			x"0000" when x"D9D2",
			x"0000" when x"D9D3",
			x"0000" when x"D9D4",
			x"0000" when x"D9D5",
			x"0000" when x"D9D6",
			x"0000" when x"D9D7",
			x"0000" when x"D9D8",
			x"0000" when x"D9D9",
			x"0000" when x"D9DA",
			x"0000" when x"D9DB",
			x"0000" when x"D9DC",
			x"0000" when x"D9DD",
			x"0000" when x"D9DE",
			x"0000" when x"D9DF",
			x"0000" when x"D9E0",
			x"0000" when x"D9E1",
			x"0000" when x"D9E2",
			x"0000" when x"D9E3",
			x"0000" when x"D9E4",
			x"0000" when x"D9E5",
			x"0000" when x"D9E6",
			x"0000" when x"D9E7",
			x"0000" when x"D9E8",
			x"0000" when x"D9E9",
			x"0000" when x"D9EA",
			x"0000" when x"D9EB",
			x"0000" when x"D9EC",
			x"0000" when x"D9ED",
			x"0000" when x"D9EE",
			x"0000" when x"D9EF",
			x"0000" when x"D9F0",
			x"0000" when x"D9F1",
			x"0000" when x"D9F2",
			x"0000" when x"D9F3",
			x"0000" when x"D9F4",
			x"0000" when x"D9F5",
			x"0000" when x"D9F6",
			x"0000" when x"D9F7",
			x"0000" when x"D9F8",
			x"0000" when x"D9F9",
			x"0000" when x"D9FA",
			x"0000" when x"D9FB",
			x"0000" when x"D9FC",
			x"0000" when x"D9FD",
			x"0000" when x"D9FE",
			x"0000" when x"D9FF",
			x"0000" when x"DA00",
			x"0000" when x"DA01",
			x"0000" when x"DA02",
			x"0000" when x"DA03",
			x"0000" when x"DA04",
			x"0000" when x"DA05",
			x"0000" when x"DA06",
			x"0000" when x"DA07",
			x"0000" when x"DA08",
			x"0000" when x"DA09",
			x"0000" when x"DA0A",
			x"0000" when x"DA0B",
			x"0000" when x"DA0C",
			x"0000" when x"DA0D",
			x"0000" when x"DA0E",
			x"0000" when x"DA0F",
			x"0000" when x"DA10",
			x"0000" when x"DA11",
			x"0000" when x"DA12",
			x"0000" when x"DA13",
			x"0000" when x"DA14",
			x"0000" when x"DA15",
			x"0000" when x"DA16",
			x"0000" when x"DA17",
			x"0000" when x"DA18",
			x"0000" when x"DA19",
			x"0000" when x"DA1A",
			x"0000" when x"DA1B",
			x"0000" when x"DA1C",
			x"0000" when x"DA1D",
			x"0000" when x"DA1E",
			x"0000" when x"DA1F",
			x"0000" when x"DA20",
			x"0000" when x"DA21",
			x"0000" when x"DA22",
			x"0000" when x"DA23",
			x"0000" when x"DA24",
			x"0000" when x"DA25",
			x"0000" when x"DA26",
			x"0000" when x"DA27",
			x"0000" when x"DA28",
			x"0000" when x"DA29",
			x"0000" when x"DA2A",
			x"0000" when x"DA2B",
			x"0000" when x"DA2C",
			x"0000" when x"DA2D",
			x"0000" when x"DA2E",
			x"0000" when x"DA2F",
			x"0000" when x"DA30",
			x"0000" when x"DA31",
			x"0000" when x"DA32",
			x"0000" when x"DA33",
			x"0000" when x"DA34",
			x"0000" when x"DA35",
			x"0000" when x"DA36",
			x"0000" when x"DA37",
			x"0000" when x"DA38",
			x"0000" when x"DA39",
			x"0000" when x"DA3A",
			x"0000" when x"DA3B",
			x"0000" when x"DA3C",
			x"0000" when x"DA3D",
			x"0000" when x"DA3E",
			x"0000" when x"DA3F",
			x"0000" when x"DA40",
			x"0000" when x"DA41",
			x"0000" when x"DA42",
			x"0000" when x"DA43",
			x"0000" when x"DA44",
			x"0000" when x"DA45",
			x"0000" when x"DA46",
			x"0000" when x"DA47",
			x"0000" when x"DA48",
			x"0000" when x"DA49",
			x"0000" when x"DA4A",
			x"0000" when x"DA4B",
			x"0000" when x"DA4C",
			x"0000" when x"DA4D",
			x"0000" when x"DA4E",
			x"0000" when x"DA4F",
			x"0000" when x"DA50",
			x"0000" when x"DA51",
			x"0000" when x"DA52",
			x"0000" when x"DA53",
			x"0000" when x"DA54",
			x"0000" when x"DA55",
			x"0000" when x"DA56",
			x"0000" when x"DA57",
			x"0000" when x"DA58",
			x"0000" when x"DA59",
			x"0000" when x"DA5A",
			x"0000" when x"DA5B",
			x"0000" when x"DA5C",
			x"0000" when x"DA5D",
			x"0000" when x"DA5E",
			x"0000" when x"DA5F",
			x"0000" when x"DA60",
			x"0000" when x"DA61",
			x"0000" when x"DA62",
			x"0000" when x"DA63",
			x"0000" when x"DA64",
			x"0000" when x"DA65",
			x"0000" when x"DA66",
			x"0000" when x"DA67",
			x"0000" when x"DA68",
			x"0000" when x"DA69",
			x"0000" when x"DA6A",
			x"0000" when x"DA6B",
			x"0000" when x"DA6C",
			x"0000" when x"DA6D",
			x"0000" when x"DA6E",
			x"0000" when x"DA6F",
			x"0000" when x"DA70",
			x"0000" when x"DA71",
			x"0000" when x"DA72",
			x"0000" when x"DA73",
			x"0000" when x"DA74",
			x"0000" when x"DA75",
			x"0000" when x"DA76",
			x"0000" when x"DA77",
			x"0000" when x"DA78",
			x"0000" when x"DA79",
			x"0000" when x"DA7A",
			x"0000" when x"DA7B",
			x"0000" when x"DA7C",
			x"0000" when x"DA7D",
			x"0000" when x"DA7E",
			x"0000" when x"DA7F",
			x"0000" when x"DA80",
			x"0000" when x"DA81",
			x"0000" when x"DA82",
			x"0000" when x"DA83",
			x"0000" when x"DA84",
			x"0000" when x"DA85",
			x"0000" when x"DA86",
			x"0000" when x"DA87",
			x"0000" when x"DA88",
			x"0000" when x"DA89",
			x"0000" when x"DA8A",
			x"0000" when x"DA8B",
			x"0000" when x"DA8C",
			x"0000" when x"DA8D",
			x"0000" when x"DA8E",
			x"0000" when x"DA8F",
			x"0000" when x"DA90",
			x"0000" when x"DA91",
			x"0000" when x"DA92",
			x"0000" when x"DA93",
			x"0000" when x"DA94",
			x"0000" when x"DA95",
			x"0000" when x"DA96",
			x"0000" when x"DA97",
			x"0000" when x"DA98",
			x"0000" when x"DA99",
			x"0000" when x"DA9A",
			x"0000" when x"DA9B",
			x"0000" when x"DA9C",
			x"0000" when x"DA9D",
			x"0000" when x"DA9E",
			x"0000" when x"DA9F",
			x"0000" when x"DAA0",
			x"0000" when x"DAA1",
			x"0000" when x"DAA2",
			x"0000" when x"DAA3",
			x"0000" when x"DAA4",
			x"0000" when x"DAA5",
			x"0000" when x"DAA6",
			x"0000" when x"DAA7",
			x"0000" when x"DAA8",
			x"0000" when x"DAA9",
			x"0000" when x"DAAA",
			x"0000" when x"DAAB",
			x"0000" when x"DAAC",
			x"0000" when x"DAAD",
			x"0000" when x"DAAE",
			x"0000" when x"DAAF",
			x"0000" when x"DAB0",
			x"0000" when x"DAB1",
			x"0000" when x"DAB2",
			x"0000" when x"DAB3",
			x"0000" when x"DAB4",
			x"0000" when x"DAB5",
			x"0000" when x"DAB6",
			x"0000" when x"DAB7",
			x"0000" when x"DAB8",
			x"0000" when x"DAB9",
			x"0000" when x"DABA",
			x"0000" when x"DABB",
			x"0000" when x"DABC",
			x"0000" when x"DABD",
			x"0000" when x"DABE",
			x"0000" when x"DABF",
			x"0000" when x"DAC0",
			x"0000" when x"DAC1",
			x"0000" when x"DAC2",
			x"0000" when x"DAC3",
			x"0000" when x"DAC4",
			x"0000" when x"DAC5",
			x"0000" when x"DAC6",
			x"0000" when x"DAC7",
			x"0000" when x"DAC8",
			x"0000" when x"DAC9",
			x"0000" when x"DACA",
			x"0000" when x"DACB",
			x"0000" when x"DACC",
			x"0000" when x"DACD",
			x"0000" when x"DACE",
			x"0000" when x"DACF",
			x"0000" when x"DAD0",
			x"0000" when x"DAD1",
			x"0000" when x"DAD2",
			x"0000" when x"DAD3",
			x"0000" when x"DAD4",
			x"0000" when x"DAD5",
			x"0000" when x"DAD6",
			x"0000" when x"DAD7",
			x"0000" when x"DAD8",
			x"0000" when x"DAD9",
			x"0000" when x"DADA",
			x"0000" when x"DADB",
			x"0000" when x"DADC",
			x"0000" when x"DADD",
			x"0000" when x"DADE",
			x"0000" when x"DADF",
			x"0000" when x"DAE0",
			x"0000" when x"DAE1",
			x"0000" when x"DAE2",
			x"0000" when x"DAE3",
			x"0000" when x"DAE4",
			x"0000" when x"DAE5",
			x"0000" when x"DAE6",
			x"0000" when x"DAE7",
			x"0000" when x"DAE8",
			x"0000" when x"DAE9",
			x"0000" when x"DAEA",
			x"0000" when x"DAEB",
			x"0000" when x"DAEC",
			x"0000" when x"DAED",
			x"0000" when x"DAEE",
			x"0000" when x"DAEF",
			x"0000" when x"DAF0",
			x"0000" when x"DAF1",
			x"0000" when x"DAF2",
			x"0000" when x"DAF3",
			x"0000" when x"DAF4",
			x"0000" when x"DAF5",
			x"0000" when x"DAF6",
			x"0000" when x"DAF7",
			x"0000" when x"DAF8",
			x"0000" when x"DAF9",
			x"0000" when x"DAFA",
			x"0000" when x"DAFB",
			x"0000" when x"DAFC",
			x"0000" when x"DAFD",
			x"0000" when x"DAFE",
			x"0000" when x"DAFF",
			x"0000" when x"DB00",
			x"0000" when x"DB01",
			x"0000" when x"DB02",
			x"0000" when x"DB03",
			x"0000" when x"DB04",
			x"0000" when x"DB05",
			x"0000" when x"DB06",
			x"0000" when x"DB07",
			x"0000" when x"DB08",
			x"0000" when x"DB09",
			x"0000" when x"DB0A",
			x"0000" when x"DB0B",
			x"0000" when x"DB0C",
			x"0000" when x"DB0D",
			x"0000" when x"DB0E",
			x"0000" when x"DB0F",
			x"0000" when x"DB10",
			x"0000" when x"DB11",
			x"0000" when x"DB12",
			x"0000" when x"DB13",
			x"0000" when x"DB14",
			x"0000" when x"DB15",
			x"0000" when x"DB16",
			x"0000" when x"DB17",
			x"0000" when x"DB18",
			x"0000" when x"DB19",
			x"0000" when x"DB1A",
			x"0000" when x"DB1B",
			x"0000" when x"DB1C",
			x"0000" when x"DB1D",
			x"0000" when x"DB1E",
			x"0000" when x"DB1F",
			x"0000" when x"DB20",
			x"0000" when x"DB21",
			x"0000" when x"DB22",
			x"0000" when x"DB23",
			x"0000" when x"DB24",
			x"0000" when x"DB25",
			x"0000" when x"DB26",
			x"0000" when x"DB27",
			x"0000" when x"DB28",
			x"0000" when x"DB29",
			x"0000" when x"DB2A",
			x"0000" when x"DB2B",
			x"0000" when x"DB2C",
			x"0000" when x"DB2D",
			x"0000" when x"DB2E",
			x"0000" when x"DB2F",
			x"0000" when x"DB30",
			x"0000" when x"DB31",
			x"0000" when x"DB32",
			x"0000" when x"DB33",
			x"0000" when x"DB34",
			x"0000" when x"DB35",
			x"0000" when x"DB36",
			x"0000" when x"DB37",
			x"0000" when x"DB38",
			x"0000" when x"DB39",
			x"0000" when x"DB3A",
			x"0000" when x"DB3B",
			x"0000" when x"DB3C",
			x"0000" when x"DB3D",
			x"0000" when x"DB3E",
			x"0000" when x"DB3F",
			x"0000" when x"DB40",
			x"0000" when x"DB41",
			x"0000" when x"DB42",
			x"0000" when x"DB43",
			x"0000" when x"DB44",
			x"0000" when x"DB45",
			x"0000" when x"DB46",
			x"0000" when x"DB47",
			x"0000" when x"DB48",
			x"0000" when x"DB49",
			x"0000" when x"DB4A",
			x"0000" when x"DB4B",
			x"0000" when x"DB4C",
			x"0000" when x"DB4D",
			x"0000" when x"DB4E",
			x"0000" when x"DB4F",
			x"0000" when x"DB50",
			x"0000" when x"DB51",
			x"0000" when x"DB52",
			x"0000" when x"DB53",
			x"0000" when x"DB54",
			x"0000" when x"DB55",
			x"0000" when x"DB56",
			x"0000" when x"DB57",
			x"0000" when x"DB58",
			x"0000" when x"DB59",
			x"0000" when x"DB5A",
			x"0000" when x"DB5B",
			x"0000" when x"DB5C",
			x"0000" when x"DB5D",
			x"0000" when x"DB5E",
			x"0000" when x"DB5F",
			x"0000" when x"DB60",
			x"0000" when x"DB61",
			x"0000" when x"DB62",
			x"0000" when x"DB63",
			x"0000" when x"DB64",
			x"0000" when x"DB65",
			x"0000" when x"DB66",
			x"0000" when x"DB67",
			x"0000" when x"DB68",
			x"0000" when x"DB69",
			x"0000" when x"DB6A",
			x"0000" when x"DB6B",
			x"0000" when x"DB6C",
			x"0000" when x"DB6D",
			x"0000" when x"DB6E",
			x"0000" when x"DB6F",
			x"0000" when x"DB70",
			x"0000" when x"DB71",
			x"0000" when x"DB72",
			x"0000" when x"DB73",
			x"0000" when x"DB74",
			x"0000" when x"DB75",
			x"0000" when x"DB76",
			x"0000" when x"DB77",
			x"0000" when x"DB78",
			x"0000" when x"DB79",
			x"0000" when x"DB7A",
			x"0000" when x"DB7B",
			x"0000" when x"DB7C",
			x"0000" when x"DB7D",
			x"0000" when x"DB7E",
			x"0000" when x"DB7F",
			x"0000" when x"DB80",
			x"0000" when x"DB81",
			x"0000" when x"DB82",
			x"0000" when x"DB83",
			x"0000" when x"DB84",
			x"0000" when x"DB85",
			x"0000" when x"DB86",
			x"0000" when x"DB87",
			x"0000" when x"DB88",
			x"0000" when x"DB89",
			x"0000" when x"DB8A",
			x"0000" when x"DB8B",
			x"0000" when x"DB8C",
			x"0000" when x"DB8D",
			x"0000" when x"DB8E",
			x"0000" when x"DB8F",
			x"0000" when x"DB90",
			x"0000" when x"DB91",
			x"0000" when x"DB92",
			x"0000" when x"DB93",
			x"0000" when x"DB94",
			x"0000" when x"DB95",
			x"0000" when x"DB96",
			x"0000" when x"DB97",
			x"0000" when x"DB98",
			x"0000" when x"DB99",
			x"0000" when x"DB9A",
			x"0000" when x"DB9B",
			x"0000" when x"DB9C",
			x"0000" when x"DB9D",
			x"0000" when x"DB9E",
			x"0000" when x"DB9F",
			x"0000" when x"DBA0",
			x"0000" when x"DBA1",
			x"0000" when x"DBA2",
			x"0000" when x"DBA3",
			x"0000" when x"DBA4",
			x"0000" when x"DBA5",
			x"0000" when x"DBA6",
			x"0000" when x"DBA7",
			x"0000" when x"DBA8",
			x"0000" when x"DBA9",
			x"0000" when x"DBAA",
			x"0000" when x"DBAB",
			x"0000" when x"DBAC",
			x"0000" when x"DBAD",
			x"0000" when x"DBAE",
			x"0000" when x"DBAF",
			x"0000" when x"DBB0",
			x"0000" when x"DBB1",
			x"0000" when x"DBB2",
			x"0000" when x"DBB3",
			x"0000" when x"DBB4",
			x"0000" when x"DBB5",
			x"0000" when x"DBB6",
			x"0000" when x"DBB7",
			x"0000" when x"DBB8",
			x"0000" when x"DBB9",
			x"0000" when x"DBBA",
			x"0000" when x"DBBB",
			x"0000" when x"DBBC",
			x"0000" when x"DBBD",
			x"0000" when x"DBBE",
			x"0000" when x"DBBF",
			x"0000" when x"DBC0",
			x"0000" when x"DBC1",
			x"0000" when x"DBC2",
			x"0000" when x"DBC3",
			x"0000" when x"DBC4",
			x"0000" when x"DBC5",
			x"0000" when x"DBC6",
			x"0000" when x"DBC7",
			x"0000" when x"DBC8",
			x"0000" when x"DBC9",
			x"0000" when x"DBCA",
			x"0000" when x"DBCB",
			x"0000" when x"DBCC",
			x"0000" when x"DBCD",
			x"0000" when x"DBCE",
			x"0000" when x"DBCF",
			x"0000" when x"DBD0",
			x"0000" when x"DBD1",
			x"0000" when x"DBD2",
			x"0000" when x"DBD3",
			x"0000" when x"DBD4",
			x"0000" when x"DBD5",
			x"0000" when x"DBD6",
			x"0000" when x"DBD7",
			x"0000" when x"DBD8",
			x"0000" when x"DBD9",
			x"0000" when x"DBDA",
			x"0000" when x"DBDB",
			x"0000" when x"DBDC",
			x"0000" when x"DBDD",
			x"0000" when x"DBDE",
			x"0000" when x"DBDF",
			x"0000" when x"DBE0",
			x"0000" when x"DBE1",
			x"0000" when x"DBE2",
			x"0000" when x"DBE3",
			x"0000" when x"DBE4",
			x"0000" when x"DBE5",
			x"0000" when x"DBE6",
			x"0000" when x"DBE7",
			x"0000" when x"DBE8",
			x"0000" when x"DBE9",
			x"0000" when x"DBEA",
			x"0000" when x"DBEB",
			x"0000" when x"DBEC",
			x"0000" when x"DBED",
			x"0000" when x"DBEE",
			x"0000" when x"DBEF",
			x"0000" when x"DBF0",
			x"0000" when x"DBF1",
			x"0000" when x"DBF2",
			x"0000" when x"DBF3",
			x"0000" when x"DBF4",
			x"0000" when x"DBF5",
			x"0000" when x"DBF6",
			x"0000" when x"DBF7",
			x"0000" when x"DBF8",
			x"0000" when x"DBF9",
			x"0000" when x"DBFA",
			x"0000" when x"DBFB",
			x"0000" when x"DBFC",
			x"0000" when x"DBFD",
			x"0000" when x"DBFE",
			x"0000" when x"DBFF",
			x"0000" when x"DC00",
			x"0000" when x"DC01",
			x"0000" when x"DC02",
			x"0000" when x"DC03",
			x"0000" when x"DC04",
			x"0000" when x"DC05",
			x"0000" when x"DC06",
			x"0000" when x"DC07",
			x"0000" when x"DC08",
			x"0000" when x"DC09",
			x"0000" when x"DC0A",
			x"0000" when x"DC0B",
			x"0000" when x"DC0C",
			x"0000" when x"DC0D",
			x"0000" when x"DC0E",
			x"0000" when x"DC0F",
			x"0000" when x"DC10",
			x"0000" when x"DC11",
			x"0000" when x"DC12",
			x"0000" when x"DC13",
			x"0000" when x"DC14",
			x"0000" when x"DC15",
			x"0000" when x"DC16",
			x"0000" when x"DC17",
			x"0000" when x"DC18",
			x"0000" when x"DC19",
			x"0000" when x"DC1A",
			x"0000" when x"DC1B",
			x"0000" when x"DC1C",
			x"0000" when x"DC1D",
			x"0000" when x"DC1E",
			x"0000" when x"DC1F",
			x"0000" when x"DC20",
			x"0000" when x"DC21",
			x"0000" when x"DC22",
			x"0000" when x"DC23",
			x"0000" when x"DC24",
			x"0000" when x"DC25",
			x"0000" when x"DC26",
			x"0000" when x"DC27",
			x"0000" when x"DC28",
			x"0000" when x"DC29",
			x"0000" when x"DC2A",
			x"0000" when x"DC2B",
			x"0000" when x"DC2C",
			x"0000" when x"DC2D",
			x"0000" when x"DC2E",
			x"0000" when x"DC2F",
			x"0000" when x"DC30",
			x"0000" when x"DC31",
			x"0000" when x"DC32",
			x"0000" when x"DC33",
			x"0000" when x"DC34",
			x"0000" when x"DC35",
			x"0000" when x"DC36",
			x"0000" when x"DC37",
			x"0000" when x"DC38",
			x"0000" when x"DC39",
			x"0000" when x"DC3A",
			x"0000" when x"DC3B",
			x"0000" when x"DC3C",
			x"0000" when x"DC3D",
			x"0000" when x"DC3E",
			x"0000" when x"DC3F",
			x"0000" when x"DC40",
			x"0000" when x"DC41",
			x"0000" when x"DC42",
			x"0000" when x"DC43",
			x"0000" when x"DC44",
			x"0000" when x"DC45",
			x"0000" when x"DC46",
			x"0000" when x"DC47",
			x"0000" when x"DC48",
			x"0000" when x"DC49",
			x"0000" when x"DC4A",
			x"0000" when x"DC4B",
			x"0000" when x"DC4C",
			x"0000" when x"DC4D",
			x"0000" when x"DC4E",
			x"0000" when x"DC4F",
			x"0000" when x"DC50",
			x"0000" when x"DC51",
			x"0000" when x"DC52",
			x"0000" when x"DC53",
			x"0000" when x"DC54",
			x"0000" when x"DC55",
			x"0000" when x"DC56",
			x"0000" when x"DC57",
			x"0000" when x"DC58",
			x"0000" when x"DC59",
			x"0000" when x"DC5A",
			x"0000" when x"DC5B",
			x"0000" when x"DC5C",
			x"0000" when x"DC5D",
			x"0000" when x"DC5E",
			x"0000" when x"DC5F",
			x"0000" when x"DC60",
			x"0000" when x"DC61",
			x"0000" when x"DC62",
			x"0000" when x"DC63",
			x"0000" when x"DC64",
			x"0000" when x"DC65",
			x"0000" when x"DC66",
			x"0000" when x"DC67",
			x"0000" when x"DC68",
			x"0000" when x"DC69",
			x"0000" when x"DC6A",
			x"0000" when x"DC6B",
			x"0000" when x"DC6C",
			x"0000" when x"DC6D",
			x"0000" when x"DC6E",
			x"0000" when x"DC6F",
			x"0000" when x"DC70",
			x"0000" when x"DC71",
			x"0000" when x"DC72",
			x"0000" when x"DC73",
			x"0000" when x"DC74",
			x"0000" when x"DC75",
			x"0000" when x"DC76",
			x"0000" when x"DC77",
			x"0000" when x"DC78",
			x"0000" when x"DC79",
			x"0000" when x"DC7A",
			x"0000" when x"DC7B",
			x"0000" when x"DC7C",
			x"0000" when x"DC7D",
			x"0000" when x"DC7E",
			x"0000" when x"DC7F",
			x"0000" when x"DC80",
			x"0000" when x"DC81",
			x"0000" when x"DC82",
			x"0000" when x"DC83",
			x"0000" when x"DC84",
			x"0000" when x"DC85",
			x"0000" when x"DC86",
			x"0000" when x"DC87",
			x"0000" when x"DC88",
			x"0000" when x"DC89",
			x"0000" when x"DC8A",
			x"0000" when x"DC8B",
			x"0000" when x"DC8C",
			x"0000" when x"DC8D",
			x"0000" when x"DC8E",
			x"0000" when x"DC8F",
			x"0000" when x"DC90",
			x"0000" when x"DC91",
			x"0000" when x"DC92",
			x"0000" when x"DC93",
			x"0000" when x"DC94",
			x"0000" when x"DC95",
			x"0000" when x"DC96",
			x"0000" when x"DC97",
			x"0000" when x"DC98",
			x"0000" when x"DC99",
			x"0000" when x"DC9A",
			x"0000" when x"DC9B",
			x"0000" when x"DC9C",
			x"0000" when x"DC9D",
			x"0000" when x"DC9E",
			x"0000" when x"DC9F",
			x"0000" when x"DCA0",
			x"0000" when x"DCA1",
			x"0000" when x"DCA2",
			x"0000" when x"DCA3",
			x"0000" when x"DCA4",
			x"0000" when x"DCA5",
			x"0000" when x"DCA6",
			x"0000" when x"DCA7",
			x"0000" when x"DCA8",
			x"0000" when x"DCA9",
			x"0000" when x"DCAA",
			x"0000" when x"DCAB",
			x"0000" when x"DCAC",
			x"0000" when x"DCAD",
			x"0000" when x"DCAE",
			x"0000" when x"DCAF",
			x"0000" when x"DCB0",
			x"0000" when x"DCB1",
			x"0000" when x"DCB2",
			x"0000" when x"DCB3",
			x"0000" when x"DCB4",
			x"0000" when x"DCB5",
			x"0000" when x"DCB6",
			x"0000" when x"DCB7",
			x"0000" when x"DCB8",
			x"0000" when x"DCB9",
			x"0000" when x"DCBA",
			x"0000" when x"DCBB",
			x"0000" when x"DCBC",
			x"0000" when x"DCBD",
			x"0000" when x"DCBE",
			x"0000" when x"DCBF",
			x"0000" when x"DCC0",
			x"0000" when x"DCC1",
			x"0000" when x"DCC2",
			x"0000" when x"DCC3",
			x"0000" when x"DCC4",
			x"0000" when x"DCC5",
			x"0000" when x"DCC6",
			x"0000" when x"DCC7",
			x"0000" when x"DCC8",
			x"0000" when x"DCC9",
			x"0000" when x"DCCA",
			x"0000" when x"DCCB",
			x"0000" when x"DCCC",
			x"0000" when x"DCCD",
			x"0000" when x"DCCE",
			x"0000" when x"DCCF",
			x"0000" when x"DCD0",
			x"0000" when x"DCD1",
			x"0000" when x"DCD2",
			x"0000" when x"DCD3",
			x"0000" when x"DCD4",
			x"0000" when x"DCD5",
			x"0000" when x"DCD6",
			x"0000" when x"DCD7",
			x"0000" when x"DCD8",
			x"0000" when x"DCD9",
			x"0000" when x"DCDA",
			x"0000" when x"DCDB",
			x"0000" when x"DCDC",
			x"0000" when x"DCDD",
			x"0000" when x"DCDE",
			x"0000" when x"DCDF",
			x"0000" when x"DCE0",
			x"0000" when x"DCE1",
			x"0000" when x"DCE2",
			x"0000" when x"DCE3",
			x"0000" when x"DCE4",
			x"0000" when x"DCE5",
			x"0000" when x"DCE6",
			x"0000" when x"DCE7",
			x"0000" when x"DCE8",
			x"0000" when x"DCE9",
			x"0000" when x"DCEA",
			x"0000" when x"DCEB",
			x"0000" when x"DCEC",
			x"0000" when x"DCED",
			x"0000" when x"DCEE",
			x"0000" when x"DCEF",
			x"0000" when x"DCF0",
			x"0000" when x"DCF1",
			x"0000" when x"DCF2",
			x"0000" when x"DCF3",
			x"0000" when x"DCF4",
			x"0000" when x"DCF5",
			x"0000" when x"DCF6",
			x"0000" when x"DCF7",
			x"0000" when x"DCF8",
			x"0000" when x"DCF9",
			x"0000" when x"DCFA",
			x"0000" when x"DCFB",
			x"0000" when x"DCFC",
			x"0000" when x"DCFD",
			x"0000" when x"DCFE",
			x"0000" when x"DCFF",
			x"0000" when x"DD00",
			x"0000" when x"DD01",
			x"0000" when x"DD02",
			x"0000" when x"DD03",
			x"0000" when x"DD04",
			x"0000" when x"DD05",
			x"0000" when x"DD06",
			x"0000" when x"DD07",
			x"0000" when x"DD08",
			x"0000" when x"DD09",
			x"0000" when x"DD0A",
			x"0000" when x"DD0B",
			x"0000" when x"DD0C",
			x"0000" when x"DD0D",
			x"0000" when x"DD0E",
			x"0000" when x"DD0F",
			x"0000" when x"DD10",
			x"0000" when x"DD11",
			x"0000" when x"DD12",
			x"0000" when x"DD13",
			x"0000" when x"DD14",
			x"0000" when x"DD15",
			x"0000" when x"DD16",
			x"0000" when x"DD17",
			x"0000" when x"DD18",
			x"0000" when x"DD19",
			x"0000" when x"DD1A",
			x"0000" when x"DD1B",
			x"0000" when x"DD1C",
			x"0000" when x"DD1D",
			x"0000" when x"DD1E",
			x"0000" when x"DD1F",
			x"0000" when x"DD20",
			x"0000" when x"DD21",
			x"0000" when x"DD22",
			x"0000" when x"DD23",
			x"0000" when x"DD24",
			x"0000" when x"DD25",
			x"0000" when x"DD26",
			x"0000" when x"DD27",
			x"0000" when x"DD28",
			x"0000" when x"DD29",
			x"0000" when x"DD2A",
			x"0000" when x"DD2B",
			x"0000" when x"DD2C",
			x"0000" when x"DD2D",
			x"0000" when x"DD2E",
			x"0000" when x"DD2F",
			x"0000" when x"DD30",
			x"0000" when x"DD31",
			x"0000" when x"DD32",
			x"0000" when x"DD33",
			x"0000" when x"DD34",
			x"0000" when x"DD35",
			x"0000" when x"DD36",
			x"0000" when x"DD37",
			x"0000" when x"DD38",
			x"0000" when x"DD39",
			x"0000" when x"DD3A",
			x"0000" when x"DD3B",
			x"0000" when x"DD3C",
			x"0000" when x"DD3D",
			x"0000" when x"DD3E",
			x"0000" when x"DD3F",
			x"0000" when x"DD40",
			x"0000" when x"DD41",
			x"0000" when x"DD42",
			x"0000" when x"DD43",
			x"0000" when x"DD44",
			x"0000" when x"DD45",
			x"0000" when x"DD46",
			x"0000" when x"DD47",
			x"0000" when x"DD48",
			x"0000" when x"DD49",
			x"0000" when x"DD4A",
			x"0000" when x"DD4B",
			x"0000" when x"DD4C",
			x"0000" when x"DD4D",
			x"0000" when x"DD4E",
			x"0000" when x"DD4F",
			x"0000" when x"DD50",
			x"0000" when x"DD51",
			x"0000" when x"DD52",
			x"0000" when x"DD53",
			x"0000" when x"DD54",
			x"0000" when x"DD55",
			x"0000" when x"DD56",
			x"0000" when x"DD57",
			x"0000" when x"DD58",
			x"0000" when x"DD59",
			x"0000" when x"DD5A",
			x"0000" when x"DD5B",
			x"0000" when x"DD5C",
			x"0000" when x"DD5D",
			x"0000" when x"DD5E",
			x"0000" when x"DD5F",
			x"0000" when x"DD60",
			x"0000" when x"DD61",
			x"0000" when x"DD62",
			x"0000" when x"DD63",
			x"0000" when x"DD64",
			x"0000" when x"DD65",
			x"0000" when x"DD66",
			x"0000" when x"DD67",
			x"0000" when x"DD68",
			x"0000" when x"DD69",
			x"0000" when x"DD6A",
			x"0000" when x"DD6B",
			x"0000" when x"DD6C",
			x"0000" when x"DD6D",
			x"0000" when x"DD6E",
			x"0000" when x"DD6F",
			x"0000" when x"DD70",
			x"0000" when x"DD71",
			x"0000" when x"DD72",
			x"0000" when x"DD73",
			x"0000" when x"DD74",
			x"0000" when x"DD75",
			x"0000" when x"DD76",
			x"0000" when x"DD77",
			x"0000" when x"DD78",
			x"0000" when x"DD79",
			x"0000" when x"DD7A",
			x"0000" when x"DD7B",
			x"0000" when x"DD7C",
			x"0000" when x"DD7D",
			x"0000" when x"DD7E",
			x"0000" when x"DD7F",
			x"0000" when x"DD80",
			x"0000" when x"DD81",
			x"0000" when x"DD82",
			x"0000" when x"DD83",
			x"0000" when x"DD84",
			x"0000" when x"DD85",
			x"0000" when x"DD86",
			x"0000" when x"DD87",
			x"0000" when x"DD88",
			x"0000" when x"DD89",
			x"0000" when x"DD8A",
			x"0000" when x"DD8B",
			x"0000" when x"DD8C",
			x"0000" when x"DD8D",
			x"0000" when x"DD8E",
			x"0000" when x"DD8F",
			x"0000" when x"DD90",
			x"0000" when x"DD91",
			x"0000" when x"DD92",
			x"0000" when x"DD93",
			x"0000" when x"DD94",
			x"0000" when x"DD95",
			x"0000" when x"DD96",
			x"0000" when x"DD97",
			x"0000" when x"DD98",
			x"0000" when x"DD99",
			x"0000" when x"DD9A",
			x"0000" when x"DD9B",
			x"0000" when x"DD9C",
			x"0000" when x"DD9D",
			x"0000" when x"DD9E",
			x"0000" when x"DD9F",
			x"0000" when x"DDA0",
			x"0000" when x"DDA1",
			x"0000" when x"DDA2",
			x"0000" when x"DDA3",
			x"0000" when x"DDA4",
			x"0000" when x"DDA5",
			x"0000" when x"DDA6",
			x"0000" when x"DDA7",
			x"0000" when x"DDA8",
			x"0000" when x"DDA9",
			x"0000" when x"DDAA",
			x"0000" when x"DDAB",
			x"0000" when x"DDAC",
			x"0000" when x"DDAD",
			x"0000" when x"DDAE",
			x"0000" when x"DDAF",
			x"0000" when x"DDB0",
			x"0000" when x"DDB1",
			x"0000" when x"DDB2",
			x"0000" when x"DDB3",
			x"0000" when x"DDB4",
			x"0000" when x"DDB5",
			x"0000" when x"DDB6",
			x"0000" when x"DDB7",
			x"0000" when x"DDB8",
			x"0000" when x"DDB9",
			x"0000" when x"DDBA",
			x"0000" when x"DDBB",
			x"0000" when x"DDBC",
			x"0000" when x"DDBD",
			x"0000" when x"DDBE",
			x"0000" when x"DDBF",
			x"0000" when x"DDC0",
			x"0000" when x"DDC1",
			x"0000" when x"DDC2",
			x"0000" when x"DDC3",
			x"0000" when x"DDC4",
			x"0000" when x"DDC5",
			x"0000" when x"DDC6",
			x"0000" when x"DDC7",
			x"0000" when x"DDC8",
			x"0000" when x"DDC9",
			x"0000" when x"DDCA",
			x"0000" when x"DDCB",
			x"0000" when x"DDCC",
			x"0000" when x"DDCD",
			x"0000" when x"DDCE",
			x"0000" when x"DDCF",
			x"0000" when x"DDD0",
			x"0000" when x"DDD1",
			x"0000" when x"DDD2",
			x"0000" when x"DDD3",
			x"0000" when x"DDD4",
			x"0000" when x"DDD5",
			x"0000" when x"DDD6",
			x"0000" when x"DDD7",
			x"0000" when x"DDD8",
			x"0000" when x"DDD9",
			x"0000" when x"DDDA",
			x"0000" when x"DDDB",
			x"0000" when x"DDDC",
			x"0000" when x"DDDD",
			x"0000" when x"DDDE",
			x"0000" when x"DDDF",
			x"0000" when x"DDE0",
			x"0000" when x"DDE1",
			x"0000" when x"DDE2",
			x"0000" when x"DDE3",
			x"0000" when x"DDE4",
			x"0000" when x"DDE5",
			x"0000" when x"DDE6",
			x"0000" when x"DDE7",
			x"0000" when x"DDE8",
			x"0000" when x"DDE9",
			x"0000" when x"DDEA",
			x"0000" when x"DDEB",
			x"0000" when x"DDEC",
			x"0000" when x"DDED",
			x"0000" when x"DDEE",
			x"0000" when x"DDEF",
			x"0000" when x"DDF0",
			x"0000" when x"DDF1",
			x"0000" when x"DDF2",
			x"0000" when x"DDF3",
			x"0000" when x"DDF4",
			x"0000" when x"DDF5",
			x"0000" when x"DDF6",
			x"0000" when x"DDF7",
			x"0000" when x"DDF8",
			x"0000" when x"DDF9",
			x"0000" when x"DDFA",
			x"0000" when x"DDFB",
			x"0000" when x"DDFC",
			x"0000" when x"DDFD",
			x"0000" when x"DDFE",
			x"0000" when x"DDFF",
			x"0000" when x"DE00",
			x"0000" when x"DE01",
			x"0000" when x"DE02",
			x"0000" when x"DE03",
			x"0000" when x"DE04",
			x"0000" when x"DE05",
			x"0000" when x"DE06",
			x"0000" when x"DE07",
			x"0000" when x"DE08",
			x"0000" when x"DE09",
			x"0000" when x"DE0A",
			x"0000" when x"DE0B",
			x"0000" when x"DE0C",
			x"0000" when x"DE0D",
			x"0000" when x"DE0E",
			x"0000" when x"DE0F",
			x"0000" when x"DE10",
			x"0000" when x"DE11",
			x"0000" when x"DE12",
			x"0000" when x"DE13",
			x"0000" when x"DE14",
			x"0000" when x"DE15",
			x"0000" when x"DE16",
			x"0000" when x"DE17",
			x"0000" when x"DE18",
			x"0000" when x"DE19",
			x"0000" when x"DE1A",
			x"0000" when x"DE1B",
			x"0000" when x"DE1C",
			x"0000" when x"DE1D",
			x"0000" when x"DE1E",
			x"0000" when x"DE1F",
			x"0000" when x"DE20",
			x"0000" when x"DE21",
			x"0000" when x"DE22",
			x"0000" when x"DE23",
			x"0000" when x"DE24",
			x"0000" when x"DE25",
			x"0000" when x"DE26",
			x"0000" when x"DE27",
			x"0000" when x"DE28",
			x"0000" when x"DE29",
			x"0000" when x"DE2A",
			x"0000" when x"DE2B",
			x"0000" when x"DE2C",
			x"0000" when x"DE2D",
			x"0000" when x"DE2E",
			x"0000" when x"DE2F",
			x"0000" when x"DE30",
			x"0000" when x"DE31",
			x"0000" when x"DE32",
			x"0000" when x"DE33",
			x"0000" when x"DE34",
			x"0000" when x"DE35",
			x"0000" when x"DE36",
			x"0000" when x"DE37",
			x"0000" when x"DE38",
			x"0000" when x"DE39",
			x"0000" when x"DE3A",
			x"0000" when x"DE3B",
			x"0000" when x"DE3C",
			x"0000" when x"DE3D",
			x"0000" when x"DE3E",
			x"0000" when x"DE3F",
			x"0000" when x"DE40",
			x"0000" when x"DE41",
			x"0000" when x"DE42",
			x"0000" when x"DE43",
			x"0000" when x"DE44",
			x"0000" when x"DE45",
			x"0000" when x"DE46",
			x"0000" when x"DE47",
			x"0000" when x"DE48",
			x"0000" when x"DE49",
			x"0000" when x"DE4A",
			x"0000" when x"DE4B",
			x"0000" when x"DE4C",
			x"0000" when x"DE4D",
			x"0000" when x"DE4E",
			x"0000" when x"DE4F",
			x"0000" when x"DE50",
			x"0000" when x"DE51",
			x"0000" when x"DE52",
			x"0000" when x"DE53",
			x"0000" when x"DE54",
			x"0000" when x"DE55",
			x"0000" when x"DE56",
			x"0000" when x"DE57",
			x"0000" when x"DE58",
			x"0000" when x"DE59",
			x"0000" when x"DE5A",
			x"0000" when x"DE5B",
			x"0000" when x"DE5C",
			x"0000" when x"DE5D",
			x"0000" when x"DE5E",
			x"0000" when x"DE5F",
			x"0000" when x"DE60",
			x"0000" when x"DE61",
			x"0000" when x"DE62",
			x"0000" when x"DE63",
			x"0000" when x"DE64",
			x"0000" when x"DE65",
			x"0000" when x"DE66",
			x"0000" when x"DE67",
			x"0000" when x"DE68",
			x"0000" when x"DE69",
			x"0000" when x"DE6A",
			x"0000" when x"DE6B",
			x"0000" when x"DE6C",
			x"0000" when x"DE6D",
			x"0000" when x"DE6E",
			x"0000" when x"DE6F",
			x"0000" when x"DE70",
			x"0000" when x"DE71",
			x"0000" when x"DE72",
			x"0000" when x"DE73",
			x"0000" when x"DE74",
			x"0000" when x"DE75",
			x"0000" when x"DE76",
			x"0000" when x"DE77",
			x"0000" when x"DE78",
			x"0000" when x"DE79",
			x"0000" when x"DE7A",
			x"0000" when x"DE7B",
			x"0000" when x"DE7C",
			x"0000" when x"DE7D",
			x"0000" when x"DE7E",
			x"0000" when x"DE7F",
			x"0000" when x"DE80",
			x"0000" when x"DE81",
			x"0000" when x"DE82",
			x"0000" when x"DE83",
			x"0000" when x"DE84",
			x"0000" when x"DE85",
			x"0000" when x"DE86",
			x"0000" when x"DE87",
			x"0000" when x"DE88",
			x"0000" when x"DE89",
			x"0000" when x"DE8A",
			x"0000" when x"DE8B",
			x"0000" when x"DE8C",
			x"0000" when x"DE8D",
			x"0000" when x"DE8E",
			x"0000" when x"DE8F",
			x"0000" when x"DE90",
			x"0000" when x"DE91",
			x"0000" when x"DE92",
			x"0000" when x"DE93",
			x"0000" when x"DE94",
			x"0000" when x"DE95",
			x"0000" when x"DE96",
			x"0000" when x"DE97",
			x"0000" when x"DE98",
			x"0000" when x"DE99",
			x"0000" when x"DE9A",
			x"0000" when x"DE9B",
			x"0000" when x"DE9C",
			x"0000" when x"DE9D",
			x"0000" when x"DE9E",
			x"0000" when x"DE9F",
			x"0000" when x"DEA0",
			x"0000" when x"DEA1",
			x"0000" when x"DEA2",
			x"0000" when x"DEA3",
			x"0000" when x"DEA4",
			x"0000" when x"DEA5",
			x"0000" when x"DEA6",
			x"0000" when x"DEA7",
			x"0000" when x"DEA8",
			x"0000" when x"DEA9",
			x"0000" when x"DEAA",
			x"0000" when x"DEAB",
			x"0000" when x"DEAC",
			x"0000" when x"DEAD",
			x"0000" when x"DEAE",
			x"0000" when x"DEAF",
			x"0000" when x"DEB0",
			x"0000" when x"DEB1",
			x"0000" when x"DEB2",
			x"0000" when x"DEB3",
			x"0000" when x"DEB4",
			x"0000" when x"DEB5",
			x"0000" when x"DEB6",
			x"0000" when x"DEB7",
			x"0000" when x"DEB8",
			x"0000" when x"DEB9",
			x"0000" when x"DEBA",
			x"0000" when x"DEBB",
			x"0000" when x"DEBC",
			x"0000" when x"DEBD",
			x"0000" when x"DEBE",
			x"0000" when x"DEBF",
			x"0000" when x"DEC0",
			x"0000" when x"DEC1",
			x"0000" when x"DEC2",
			x"0000" when x"DEC3",
			x"0000" when x"DEC4",
			x"0000" when x"DEC5",
			x"0000" when x"DEC6",
			x"0000" when x"DEC7",
			x"0000" when x"DEC8",
			x"0000" when x"DEC9",
			x"0000" when x"DECA",
			x"0000" when x"DECB",
			x"0000" when x"DECC",
			x"0000" when x"DECD",
			x"0000" when x"DECE",
			x"0000" when x"DECF",
			x"0000" when x"DED0",
			x"0000" when x"DED1",
			x"0000" when x"DED2",
			x"0000" when x"DED3",
			x"0000" when x"DED4",
			x"0000" when x"DED5",
			x"0000" when x"DED6",
			x"0000" when x"DED7",
			x"0000" when x"DED8",
			x"0000" when x"DED9",
			x"0000" when x"DEDA",
			x"0000" when x"DEDB",
			x"0000" when x"DEDC",
			x"0000" when x"DEDD",
			x"0000" when x"DEDE",
			x"0000" when x"DEDF",
			x"0000" when x"DEE0",
			x"0000" when x"DEE1",
			x"0000" when x"DEE2",
			x"0000" when x"DEE3",
			x"0000" when x"DEE4",
			x"0000" when x"DEE5",
			x"0000" when x"DEE6",
			x"0000" when x"DEE7",
			x"0000" when x"DEE8",
			x"0000" when x"DEE9",
			x"0000" when x"DEEA",
			x"0000" when x"DEEB",
			x"0000" when x"DEEC",
			x"0000" when x"DEED",
			x"0000" when x"DEEE",
			x"0000" when x"DEEF",
			x"0000" when x"DEF0",
			x"0000" when x"DEF1",
			x"0000" when x"DEF2",
			x"0000" when x"DEF3",
			x"0000" when x"DEF4",
			x"0000" when x"DEF5",
			x"0000" when x"DEF6",
			x"0000" when x"DEF7",
			x"0000" when x"DEF8",
			x"0000" when x"DEF9",
			x"0000" when x"DEFA",
			x"0000" when x"DEFB",
			x"0000" when x"DEFC",
			x"0000" when x"DEFD",
			x"0000" when x"DEFE",
			x"0000" when x"DEFF",
			x"0000" when x"DF00",
			x"0000" when x"DF01",
			x"0000" when x"DF02",
			x"0000" when x"DF03",
			x"0000" when x"DF04",
			x"0000" when x"DF05",
			x"0000" when x"DF06",
			x"0000" when x"DF07",
			x"0000" when x"DF08",
			x"0000" when x"DF09",
			x"0000" when x"DF0A",
			x"0000" when x"DF0B",
			x"0000" when x"DF0C",
			x"0000" when x"DF0D",
			x"0000" when x"DF0E",
			x"0000" when x"DF0F",
			x"0000" when x"DF10",
			x"0000" when x"DF11",
			x"0000" when x"DF12",
			x"0000" when x"DF13",
			x"0000" when x"DF14",
			x"0000" when x"DF15",
			x"0000" when x"DF16",
			x"0000" when x"DF17",
			x"0000" when x"DF18",
			x"0000" when x"DF19",
			x"0000" when x"DF1A",
			x"0000" when x"DF1B",
			x"0000" when x"DF1C",
			x"0000" when x"DF1D",
			x"0000" when x"DF1E",
			x"0000" when x"DF1F",
			x"0000" when x"DF20",
			x"0000" when x"DF21",
			x"0000" when x"DF22",
			x"0000" when x"DF23",
			x"0000" when x"DF24",
			x"0000" when x"DF25",
			x"0000" when x"DF26",
			x"0000" when x"DF27",
			x"0000" when x"DF28",
			x"0000" when x"DF29",
			x"0000" when x"DF2A",
			x"0000" when x"DF2B",
			x"0000" when x"DF2C",
			x"0000" when x"DF2D",
			x"0000" when x"DF2E",
			x"0000" when x"DF2F",
			x"0000" when x"DF30",
			x"0000" when x"DF31",
			x"0000" when x"DF32",
			x"0000" when x"DF33",
			x"0000" when x"DF34",
			x"0000" when x"DF35",
			x"0000" when x"DF36",
			x"0000" when x"DF37",
			x"0000" when x"DF38",
			x"0000" when x"DF39",
			x"0000" when x"DF3A",
			x"0000" when x"DF3B",
			x"0000" when x"DF3C",
			x"0000" when x"DF3D",
			x"0000" when x"DF3E",
			x"0000" when x"DF3F",
			x"0000" when x"DF40",
			x"0000" when x"DF41",
			x"0000" when x"DF42",
			x"0000" when x"DF43",
			x"0000" when x"DF44",
			x"0000" when x"DF45",
			x"0000" when x"DF46",
			x"0000" when x"DF47",
			x"0000" when x"DF48",
			x"0000" when x"DF49",
			x"0000" when x"DF4A",
			x"0000" when x"DF4B",
			x"0000" when x"DF4C",
			x"0000" when x"DF4D",
			x"0000" when x"DF4E",
			x"0000" when x"DF4F",
			x"0000" when x"DF50",
			x"0000" when x"DF51",
			x"0000" when x"DF52",
			x"0000" when x"DF53",
			x"0000" when x"DF54",
			x"0000" when x"DF55",
			x"0000" when x"DF56",
			x"0000" when x"DF57",
			x"0000" when x"DF58",
			x"0000" when x"DF59",
			x"0000" when x"DF5A",
			x"0000" when x"DF5B",
			x"0000" when x"DF5C",
			x"0000" when x"DF5D",
			x"0000" when x"DF5E",
			x"0000" when x"DF5F",
			x"0000" when x"DF60",
			x"0000" when x"DF61",
			x"0000" when x"DF62",
			x"0000" when x"DF63",
			x"0000" when x"DF64",
			x"0000" when x"DF65",
			x"0000" when x"DF66",
			x"0000" when x"DF67",
			x"0000" when x"DF68",
			x"0000" when x"DF69",
			x"0000" when x"DF6A",
			x"0000" when x"DF6B",
			x"0000" when x"DF6C",
			x"0000" when x"DF6D",
			x"0000" when x"DF6E",
			x"0000" when x"DF6F",
			x"0000" when x"DF70",
			x"0000" when x"DF71",
			x"0000" when x"DF72",
			x"0000" when x"DF73",
			x"0000" when x"DF74",
			x"0000" when x"DF75",
			x"0000" when x"DF76",
			x"0000" when x"DF77",
			x"0000" when x"DF78",
			x"0000" when x"DF79",
			x"0000" when x"DF7A",
			x"0000" when x"DF7B",
			x"0000" when x"DF7C",
			x"0000" when x"DF7D",
			x"0000" when x"DF7E",
			x"0000" when x"DF7F",
			x"0000" when x"DF80",
			x"0000" when x"DF81",
			x"0000" when x"DF82",
			x"0000" when x"DF83",
			x"0000" when x"DF84",
			x"0000" when x"DF85",
			x"0000" when x"DF86",
			x"0000" when x"DF87",
			x"0000" when x"DF88",
			x"0000" when x"DF89",
			x"0000" when x"DF8A",
			x"0000" when x"DF8B",
			x"0000" when x"DF8C",
			x"0000" when x"DF8D",
			x"0000" when x"DF8E",
			x"0000" when x"DF8F",
			x"0000" when x"DF90",
			x"0000" when x"DF91",
			x"0000" when x"DF92",
			x"0000" when x"DF93",
			x"0000" when x"DF94",
			x"0000" when x"DF95",
			x"0000" when x"DF96",
			x"0000" when x"DF97",
			x"0000" when x"DF98",
			x"0000" when x"DF99",
			x"0000" when x"DF9A",
			x"0000" when x"DF9B",
			x"0000" when x"DF9C",
			x"0000" when x"DF9D",
			x"0000" when x"DF9E",
			x"0000" when x"DF9F",
			x"0000" when x"DFA0",
			x"0000" when x"DFA1",
			x"0000" when x"DFA2",
			x"0000" when x"DFA3",
			x"0000" when x"DFA4",
			x"0000" when x"DFA5",
			x"0000" when x"DFA6",
			x"0000" when x"DFA7",
			x"0000" when x"DFA8",
			x"0000" when x"DFA9",
			x"0000" when x"DFAA",
			x"0000" when x"DFAB",
			x"0000" when x"DFAC",
			x"0000" when x"DFAD",
			x"0000" when x"DFAE",
			x"0000" when x"DFAF",
			x"0000" when x"DFB0",
			x"0000" when x"DFB1",
			x"0000" when x"DFB2",
			x"0000" when x"DFB3",
			x"0000" when x"DFB4",
			x"0000" when x"DFB5",
			x"0000" when x"DFB6",
			x"0000" when x"DFB7",
			x"0000" when x"DFB8",
			x"0000" when x"DFB9",
			x"0000" when x"DFBA",
			x"0000" when x"DFBB",
			x"0000" when x"DFBC",
			x"0000" when x"DFBD",
			x"0000" when x"DFBE",
			x"0000" when x"DFBF",
			x"0000" when x"DFC0",
			x"0000" when x"DFC1",
			x"0000" when x"DFC2",
			x"0000" when x"DFC3",
			x"0000" when x"DFC4",
			x"0000" when x"DFC5",
			x"0000" when x"DFC6",
			x"0000" when x"DFC7",
			x"0000" when x"DFC8",
			x"0000" when x"DFC9",
			x"0000" when x"DFCA",
			x"0000" when x"DFCB",
			x"0000" when x"DFCC",
			x"0000" when x"DFCD",
			x"0000" when x"DFCE",
			x"0000" when x"DFCF",
			x"0000" when x"DFD0",
			x"0000" when x"DFD1",
			x"0000" when x"DFD2",
			x"0000" when x"DFD3",
			x"0000" when x"DFD4",
			x"0000" when x"DFD5",
			x"0000" when x"DFD6",
			x"0000" when x"DFD7",
			x"0000" when x"DFD8",
			x"0000" when x"DFD9",
			x"0000" when x"DFDA",
			x"0000" when x"DFDB",
			x"0000" when x"DFDC",
			x"0000" when x"DFDD",
			x"0000" when x"DFDE",
			x"0000" when x"DFDF",
			x"0000" when x"DFE0",
			x"0000" when x"DFE1",
			x"0000" when x"DFE2",
			x"0000" when x"DFE3",
			x"0000" when x"DFE4",
			x"0000" when x"DFE5",
			x"0000" when x"DFE6",
			x"0000" when x"DFE7",
			x"0000" when x"DFE8",
			x"0000" when x"DFE9",
			x"0000" when x"DFEA",
			x"0000" when x"DFEB",
			x"0000" when x"DFEC",
			x"0000" when x"DFED",
			x"0000" when x"DFEE",
			x"0000" when x"DFEF",
			x"0000" when x"DFF0",
			x"0000" when x"DFF1",
			x"0000" when x"DFF2",
			x"0000" when x"DFF3",
			x"0000" when x"DFF4",
			x"0000" when x"DFF5",
			x"0000" when x"DFF6",
			x"0000" when x"DFF7",
			x"0000" when x"DFF8",
			x"0000" when x"DFF9",
			x"0000" when x"DFFA",
			x"0000" when x"DFFB",
			x"0000" when x"DFFC",
			x"0000" when x"DFFD",
			x"0000" when x"DFFE",
			x"0000" when x"DFFF",
			x"0000" when x"E000",
			x"0000" when x"E001",
			x"0000" when x"E002",
			x"0000" when x"E003",
			x"0000" when x"E004",
			x"0000" when x"E005",
			x"0000" when x"E006",
			x"0000" when x"E007",
			x"0000" when x"E008",
			x"0000" when x"E009",
			x"0000" when x"E00A",
			x"0000" when x"E00B",
			x"0000" when x"E00C",
			x"0000" when x"E00D",
			x"0000" when x"E00E",
			x"0000" when x"E00F",
			x"0000" when x"E010",
			x"0000" when x"E011",
			x"0000" when x"E012",
			x"0000" when x"E013",
			x"0000" when x"E014",
			x"0000" when x"E015",
			x"0000" when x"E016",
			x"0000" when x"E017",
			x"0000" when x"E018",
			x"0000" when x"E019",
			x"0000" when x"E01A",
			x"0000" when x"E01B",
			x"0000" when x"E01C",
			x"0000" when x"E01D",
			x"0000" when x"E01E",
			x"0000" when x"E01F",
			x"0000" when x"E020",
			x"0000" when x"E021",
			x"0000" when x"E022",
			x"0000" when x"E023",
			x"0000" when x"E024",
			x"0000" when x"E025",
			x"0000" when x"E026",
			x"0000" when x"E027",
			x"0000" when x"E028",
			x"0000" when x"E029",
			x"0000" when x"E02A",
			x"0000" when x"E02B",
			x"0000" when x"E02C",
			x"0000" when x"E02D",
			x"0000" when x"E02E",
			x"0000" when x"E02F",
			x"0000" when x"E030",
			x"0000" when x"E031",
			x"0000" when x"E032",
			x"0000" when x"E033",
			x"0000" when x"E034",
			x"0000" when x"E035",
			x"0000" when x"E036",
			x"0000" when x"E037",
			x"0000" when x"E038",
			x"0000" when x"E039",
			x"0000" when x"E03A",
			x"0000" when x"E03B",
			x"0000" when x"E03C",
			x"0000" when x"E03D",
			x"0000" when x"E03E",
			x"0000" when x"E03F",
			x"0000" when x"E040",
			x"0000" when x"E041",
			x"0000" when x"E042",
			x"0000" when x"E043",
			x"0000" when x"E044",
			x"0000" when x"E045",
			x"0000" when x"E046",
			x"0000" when x"E047",
			x"0000" when x"E048",
			x"0000" when x"E049",
			x"0000" when x"E04A",
			x"0000" when x"E04B",
			x"0000" when x"E04C",
			x"0000" when x"E04D",
			x"0000" when x"E04E",
			x"0000" when x"E04F",
			x"0000" when x"E050",
			x"0000" when x"E051",
			x"0000" when x"E052",
			x"0000" when x"E053",
			x"0000" when x"E054",
			x"0000" when x"E055",
			x"0000" when x"E056",
			x"0000" when x"E057",
			x"0000" when x"E058",
			x"0000" when x"E059",
			x"0000" when x"E05A",
			x"0000" when x"E05B",
			x"0000" when x"E05C",
			x"0000" when x"E05D",
			x"0000" when x"E05E",
			x"0000" when x"E05F",
			x"0000" when x"E060",
			x"0000" when x"E061",
			x"0000" when x"E062",
			x"0000" when x"E063",
			x"0000" when x"E064",
			x"0000" when x"E065",
			x"0000" when x"E066",
			x"0000" when x"E067",
			x"0000" when x"E068",
			x"0000" when x"E069",
			x"0000" when x"E06A",
			x"0000" when x"E06B",
			x"0000" when x"E06C",
			x"0000" when x"E06D",
			x"0000" when x"E06E",
			x"0000" when x"E06F",
			x"0000" when x"E070",
			x"0000" when x"E071",
			x"0000" when x"E072",
			x"0000" when x"E073",
			x"0000" when x"E074",
			x"0000" when x"E075",
			x"0000" when x"E076",
			x"0000" when x"E077",
			x"0000" when x"E078",
			x"0000" when x"E079",
			x"0000" when x"E07A",
			x"0000" when x"E07B",
			x"0000" when x"E07C",
			x"0000" when x"E07D",
			x"0000" when x"E07E",
			x"0000" when x"E07F",
			x"0000" when x"E080",
			x"0000" when x"E081",
			x"0000" when x"E082",
			x"0000" when x"E083",
			x"0000" when x"E084",
			x"0000" when x"E085",
			x"0000" when x"E086",
			x"0000" when x"E087",
			x"0000" when x"E088",
			x"0000" when x"E089",
			x"0000" when x"E08A",
			x"0000" when x"E08B",
			x"0000" when x"E08C",
			x"0000" when x"E08D",
			x"0000" when x"E08E",
			x"0000" when x"E08F",
			x"0000" when x"E090",
			x"0000" when x"E091",
			x"0000" when x"E092",
			x"0000" when x"E093",
			x"0000" when x"E094",
			x"0000" when x"E095",
			x"0000" when x"E096",
			x"0000" when x"E097",
			x"0000" when x"E098",
			x"0000" when x"E099",
			x"0000" when x"E09A",
			x"0000" when x"E09B",
			x"0000" when x"E09C",
			x"0000" when x"E09D",
			x"0000" when x"E09E",
			x"0000" when x"E09F",
			x"0000" when x"E0A0",
			x"0000" when x"E0A1",
			x"0000" when x"E0A2",
			x"0000" when x"E0A3",
			x"0000" when x"E0A4",
			x"0000" when x"E0A5",
			x"0000" when x"E0A6",
			x"0000" when x"E0A7",
			x"0000" when x"E0A8",
			x"0000" when x"E0A9",
			x"0000" when x"E0AA",
			x"0000" when x"E0AB",
			x"0000" when x"E0AC",
			x"0000" when x"E0AD",
			x"0000" when x"E0AE",
			x"0000" when x"E0AF",
			x"0000" when x"E0B0",
			x"0000" when x"E0B1",
			x"0000" when x"E0B2",
			x"0000" when x"E0B3",
			x"0000" when x"E0B4",
			x"0000" when x"E0B5",
			x"0000" when x"E0B6",
			x"0000" when x"E0B7",
			x"0000" when x"E0B8",
			x"0000" when x"E0B9",
			x"0000" when x"E0BA",
			x"0000" when x"E0BB",
			x"0000" when x"E0BC",
			x"0000" when x"E0BD",
			x"0000" when x"E0BE",
			x"0000" when x"E0BF",
			x"0000" when x"E0C0",
			x"0000" when x"E0C1",
			x"0000" when x"E0C2",
			x"0000" when x"E0C3",
			x"0000" when x"E0C4",
			x"0000" when x"E0C5",
			x"0000" when x"E0C6",
			x"0000" when x"E0C7",
			x"0000" when x"E0C8",
			x"0000" when x"E0C9",
			x"0000" when x"E0CA",
			x"0000" when x"E0CB",
			x"0000" when x"E0CC",
			x"0000" when x"E0CD",
			x"0000" when x"E0CE",
			x"0000" when x"E0CF",
			x"0000" when x"E0D0",
			x"0000" when x"E0D1",
			x"0000" when x"E0D2",
			x"0000" when x"E0D3",
			x"0000" when x"E0D4",
			x"0000" when x"E0D5",
			x"0000" when x"E0D6",
			x"0000" when x"E0D7",
			x"0000" when x"E0D8",
			x"0000" when x"E0D9",
			x"0000" when x"E0DA",
			x"0000" when x"E0DB",
			x"0000" when x"E0DC",
			x"0000" when x"E0DD",
			x"0000" when x"E0DE",
			x"0000" when x"E0DF",
			x"0000" when x"E0E0",
			x"0000" when x"E0E1",
			x"0000" when x"E0E2",
			x"0000" when x"E0E3",
			x"0000" when x"E0E4",
			x"0000" when x"E0E5",
			x"0000" when x"E0E6",
			x"0000" when x"E0E7",
			x"0000" when x"E0E8",
			x"0000" when x"E0E9",
			x"0000" when x"E0EA",
			x"0000" when x"E0EB",
			x"0000" when x"E0EC",
			x"0000" when x"E0ED",
			x"0000" when x"E0EE",
			x"0000" when x"E0EF",
			x"0000" when x"E0F0",
			x"0000" when x"E0F1",
			x"0000" when x"E0F2",
			x"0000" when x"E0F3",
			x"0000" when x"E0F4",
			x"0000" when x"E0F5",
			x"0000" when x"E0F6",
			x"0000" when x"E0F7",
			x"0000" when x"E0F8",
			x"0000" when x"E0F9",
			x"0000" when x"E0FA",
			x"0000" when x"E0FB",
			x"0000" when x"E0FC",
			x"0000" when x"E0FD",
			x"0000" when x"E0FE",
			x"0000" when x"E0FF",
			x"0000" when x"E100",
			x"0000" when x"E101",
			x"0000" when x"E102",
			x"0000" when x"E103",
			x"0000" when x"E104",
			x"0000" when x"E105",
			x"0000" when x"E106",
			x"0000" when x"E107",
			x"0000" when x"E108",
			x"0000" when x"E109",
			x"0000" when x"E10A",
			x"0000" when x"E10B",
			x"0000" when x"E10C",
			x"0000" when x"E10D",
			x"0000" when x"E10E",
			x"0000" when x"E10F",
			x"0000" when x"E110",
			x"0000" when x"E111",
			x"0000" when x"E112",
			x"0000" when x"E113",
			x"0000" when x"E114",
			x"0000" when x"E115",
			x"0000" when x"E116",
			x"0000" when x"E117",
			x"0000" when x"E118",
			x"0000" when x"E119",
			x"0000" when x"E11A",
			x"0000" when x"E11B",
			x"0000" when x"E11C",
			x"0000" when x"E11D",
			x"0000" when x"E11E",
			x"0000" when x"E11F",
			x"0000" when x"E120",
			x"0000" when x"E121",
			x"0000" when x"E122",
			x"0000" when x"E123",
			x"0000" when x"E124",
			x"0000" when x"E125",
			x"0000" when x"E126",
			x"0000" when x"E127",
			x"0000" when x"E128",
			x"0000" when x"E129",
			x"0000" when x"E12A",
			x"0000" when x"E12B",
			x"0000" when x"E12C",
			x"0000" when x"E12D",
			x"0000" when x"E12E",
			x"0000" when x"E12F",
			x"0000" when x"E130",
			x"0000" when x"E131",
			x"0000" when x"E132",
			x"0000" when x"E133",
			x"0000" when x"E134",
			x"0000" when x"E135",
			x"0000" when x"E136",
			x"0000" when x"E137",
			x"0000" when x"E138",
			x"0000" when x"E139",
			x"0000" when x"E13A",
			x"0000" when x"E13B",
			x"0000" when x"E13C",
			x"0000" when x"E13D",
			x"0000" when x"E13E",
			x"0000" when x"E13F",
			x"0000" when x"E140",
			x"0000" when x"E141",
			x"0000" when x"E142",
			x"0000" when x"E143",
			x"0000" when x"E144",
			x"0000" when x"E145",
			x"0000" when x"E146",
			x"0000" when x"E147",
			x"0000" when x"E148",
			x"0000" when x"E149",
			x"0000" when x"E14A",
			x"0000" when x"E14B",
			x"0000" when x"E14C",
			x"0000" when x"E14D",
			x"0000" when x"E14E",
			x"0000" when x"E14F",
			x"0000" when x"E150",
			x"0000" when x"E151",
			x"0000" when x"E152",
			x"0000" when x"E153",
			x"0000" when x"E154",
			x"0000" when x"E155",
			x"0000" when x"E156",
			x"0000" when x"E157",
			x"0000" when x"E158",
			x"0000" when x"E159",
			x"0000" when x"E15A",
			x"0000" when x"E15B",
			x"0000" when x"E15C",
			x"0000" when x"E15D",
			x"0000" when x"E15E",
			x"0000" when x"E15F",
			x"0000" when x"E160",
			x"0000" when x"E161",
			x"0000" when x"E162",
			x"0000" when x"E163",
			x"0000" when x"E164",
			x"0000" when x"E165",
			x"0000" when x"E166",
			x"0000" when x"E167",
			x"0000" when x"E168",
			x"0000" when x"E169",
			x"0000" when x"E16A",
			x"0000" when x"E16B",
			x"0000" when x"E16C",
			x"0000" when x"E16D",
			x"0000" when x"E16E",
			x"0000" when x"E16F",
			x"0000" when x"E170",
			x"0000" when x"E171",
			x"0000" when x"E172",
			x"0000" when x"E173",
			x"0000" when x"E174",
			x"0000" when x"E175",
			x"0000" when x"E176",
			x"0000" when x"E177",
			x"0000" when x"E178",
			x"0000" when x"E179",
			x"0000" when x"E17A",
			x"0000" when x"E17B",
			x"0000" when x"E17C",
			x"0000" when x"E17D",
			x"0000" when x"E17E",
			x"0000" when x"E17F",
			x"0000" when x"E180",
			x"0000" when x"E181",
			x"0000" when x"E182",
			x"0000" when x"E183",
			x"0000" when x"E184",
			x"0000" when x"E185",
			x"0000" when x"E186",
			x"0000" when x"E187",
			x"0000" when x"E188",
			x"0000" when x"E189",
			x"0000" when x"E18A",
			x"0000" when x"E18B",
			x"0000" when x"E18C",
			x"0000" when x"E18D",
			x"0000" when x"E18E",
			x"0000" when x"E18F",
			x"0000" when x"E190",
			x"0000" when x"E191",
			x"0000" when x"E192",
			x"0000" when x"E193",
			x"0000" when x"E194",
			x"0000" when x"E195",
			x"0000" when x"E196",
			x"0000" when x"E197",
			x"0000" when x"E198",
			x"0000" when x"E199",
			x"0000" when x"E19A",
			x"0000" when x"E19B",
			x"0000" when x"E19C",
			x"0000" when x"E19D",
			x"0000" when x"E19E",
			x"0000" when x"E19F",
			x"0000" when x"E1A0",
			x"0000" when x"E1A1",
			x"0000" when x"E1A2",
			x"0000" when x"E1A3",
			x"0000" when x"E1A4",
			x"0000" when x"E1A5",
			x"0000" when x"E1A6",
			x"0000" when x"E1A7",
			x"0000" when x"E1A8",
			x"0000" when x"E1A9",
			x"0000" when x"E1AA",
			x"0000" when x"E1AB",
			x"0000" when x"E1AC",
			x"0000" when x"E1AD",
			x"0000" when x"E1AE",
			x"0000" when x"E1AF",
			x"0000" when x"E1B0",
			x"0000" when x"E1B1",
			x"0000" when x"E1B2",
			x"0000" when x"E1B3",
			x"0000" when x"E1B4",
			x"0000" when x"E1B5",
			x"0000" when x"E1B6",
			x"0000" when x"E1B7",
			x"0000" when x"E1B8",
			x"0000" when x"E1B9",
			x"0000" when x"E1BA",
			x"0000" when x"E1BB",
			x"0000" when x"E1BC",
			x"0000" when x"E1BD",
			x"0000" when x"E1BE",
			x"0000" when x"E1BF",
			x"0000" when x"E1C0",
			x"0000" when x"E1C1",
			x"0000" when x"E1C2",
			x"0000" when x"E1C3",
			x"0000" when x"E1C4",
			x"0000" when x"E1C5",
			x"0000" when x"E1C6",
			x"0000" when x"E1C7",
			x"0000" when x"E1C8",
			x"0000" when x"E1C9",
			x"0000" when x"E1CA",
			x"0000" when x"E1CB",
			x"0000" when x"E1CC",
			x"0000" when x"E1CD",
			x"0000" when x"E1CE",
			x"0000" when x"E1CF",
			x"0000" when x"E1D0",
			x"0000" when x"E1D1",
			x"0000" when x"E1D2",
			x"0000" when x"E1D3",
			x"0000" when x"E1D4",
			x"0000" when x"E1D5",
			x"0000" when x"E1D6",
			x"0000" when x"E1D7",
			x"0000" when x"E1D8",
			x"0000" when x"E1D9",
			x"0000" when x"E1DA",
			x"0000" when x"E1DB",
			x"0000" when x"E1DC",
			x"0000" when x"E1DD",
			x"0000" when x"E1DE",
			x"0000" when x"E1DF",
			x"0000" when x"E1E0",
			x"0000" when x"E1E1",
			x"0000" when x"E1E2",
			x"0000" when x"E1E3",
			x"0000" when x"E1E4",
			x"0000" when x"E1E5",
			x"0000" when x"E1E6",
			x"0000" when x"E1E7",
			x"0000" when x"E1E8",
			x"0000" when x"E1E9",
			x"0000" when x"E1EA",
			x"0000" when x"E1EB",
			x"0000" when x"E1EC",
			x"0000" when x"E1ED",
			x"0000" when x"E1EE",
			x"0000" when x"E1EF",
			x"0000" when x"E1F0",
			x"0000" when x"E1F1",
			x"0000" when x"E1F2",
			x"0000" when x"E1F3",
			x"0000" when x"E1F4",
			x"0000" when x"E1F5",
			x"0000" when x"E1F6",
			x"0000" when x"E1F7",
			x"0000" when x"E1F8",
			x"0000" when x"E1F9",
			x"0000" when x"E1FA",
			x"0000" when x"E1FB",
			x"0000" when x"E1FC",
			x"0000" when x"E1FD",
			x"0000" when x"E1FE",
			x"0000" when x"E1FF",
			x"0000" when x"E200",
			x"0000" when x"E201",
			x"0000" when x"E202",
			x"0000" when x"E203",
			x"0000" when x"E204",
			x"0000" when x"E205",
			x"0000" when x"E206",
			x"0000" when x"E207",
			x"0000" when x"E208",
			x"0000" when x"E209",
			x"0000" when x"E20A",
			x"0000" when x"E20B",
			x"0000" when x"E20C",
			x"0000" when x"E20D",
			x"0000" when x"E20E",
			x"0000" when x"E20F",
			x"0000" when x"E210",
			x"0000" when x"E211",
			x"0000" when x"E212",
			x"0000" when x"E213",
			x"0000" when x"E214",
			x"0000" when x"E215",
			x"0000" when x"E216",
			x"0000" when x"E217",
			x"0000" when x"E218",
			x"0000" when x"E219",
			x"0000" when x"E21A",
			x"0000" when x"E21B",
			x"0000" when x"E21C",
			x"0000" when x"E21D",
			x"0000" when x"E21E",
			x"0000" when x"E21F",
			x"0000" when x"E220",
			x"0000" when x"E221",
			x"0000" when x"E222",
			x"0000" when x"E223",
			x"0000" when x"E224",
			x"0000" when x"E225",
			x"0000" when x"E226",
			x"0000" when x"E227",
			x"0000" when x"E228",
			x"0000" when x"E229",
			x"0000" when x"E22A",
			x"0000" when x"E22B",
			x"0000" when x"E22C",
			x"0000" when x"E22D",
			x"0000" when x"E22E",
			x"0000" when x"E22F",
			x"0000" when x"E230",
			x"0000" when x"E231",
			x"0000" when x"E232",
			x"0000" when x"E233",
			x"0000" when x"E234",
			x"0000" when x"E235",
			x"0000" when x"E236",
			x"0000" when x"E237",
			x"0000" when x"E238",
			x"0000" when x"E239",
			x"0000" when x"E23A",
			x"0000" when x"E23B",
			x"0000" when x"E23C",
			x"0000" when x"E23D",
			x"0000" when x"E23E",
			x"0000" when x"E23F",
			x"0000" when x"E240",
			x"0000" when x"E241",
			x"0000" when x"E242",
			x"0000" when x"E243",
			x"0000" when x"E244",
			x"0000" when x"E245",
			x"0000" when x"E246",
			x"0000" when x"E247",
			x"0000" when x"E248",
			x"0000" when x"E249",
			x"0000" when x"E24A",
			x"0000" when x"E24B",
			x"0000" when x"E24C",
			x"0000" when x"E24D",
			x"0000" when x"E24E",
			x"0000" when x"E24F",
			x"0000" when x"E250",
			x"0000" when x"E251",
			x"0000" when x"E252",
			x"0000" when x"E253",
			x"0000" when x"E254",
			x"0000" when x"E255",
			x"0000" when x"E256",
			x"0000" when x"E257",
			x"0000" when x"E258",
			x"0000" when x"E259",
			x"0000" when x"E25A",
			x"0000" when x"E25B",
			x"0000" when x"E25C",
			x"0000" when x"E25D",
			x"0000" when x"E25E",
			x"0000" when x"E25F",
			x"0000" when x"E260",
			x"0000" when x"E261",
			x"0000" when x"E262",
			x"0000" when x"E263",
			x"0000" when x"E264",
			x"0000" when x"E265",
			x"0000" when x"E266",
			x"0000" when x"E267",
			x"0000" when x"E268",
			x"0000" when x"E269",
			x"0000" when x"E26A",
			x"0000" when x"E26B",
			x"0000" when x"E26C",
			x"0000" when x"E26D",
			x"0000" when x"E26E",
			x"0000" when x"E26F",
			x"0000" when x"E270",
			x"0000" when x"E271",
			x"0000" when x"E272",
			x"0000" when x"E273",
			x"0000" when x"E274",
			x"0000" when x"E275",
			x"0000" when x"E276",
			x"0000" when x"E277",
			x"0000" when x"E278",
			x"0000" when x"E279",
			x"0000" when x"E27A",
			x"0000" when x"E27B",
			x"0000" when x"E27C",
			x"0000" when x"E27D",
			x"0000" when x"E27E",
			x"0000" when x"E27F",
			x"0000" when x"E280",
			x"0000" when x"E281",
			x"0000" when x"E282",
			x"0000" when x"E283",
			x"0000" when x"E284",
			x"0000" when x"E285",
			x"0000" when x"E286",
			x"0000" when x"E287",
			x"0000" when x"E288",
			x"0000" when x"E289",
			x"0000" when x"E28A",
			x"0000" when x"E28B",
			x"0000" when x"E28C",
			x"0000" when x"E28D",
			x"0000" when x"E28E",
			x"0000" when x"E28F",
			x"0000" when x"E290",
			x"0000" when x"E291",
			x"0000" when x"E292",
			x"0000" when x"E293",
			x"0000" when x"E294",
			x"0000" when x"E295",
			x"0000" when x"E296",
			x"0000" when x"E297",
			x"0000" when x"E298",
			x"0000" when x"E299",
			x"0000" when x"E29A",
			x"0000" when x"E29B",
			x"0000" when x"E29C",
			x"0000" when x"E29D",
			x"0000" when x"E29E",
			x"0000" when x"E29F",
			x"0000" when x"E2A0",
			x"0000" when x"E2A1",
			x"0000" when x"E2A2",
			x"0000" when x"E2A3",
			x"0000" when x"E2A4",
			x"0000" when x"E2A5",
			x"0000" when x"E2A6",
			x"0000" when x"E2A7",
			x"0000" when x"E2A8",
			x"0000" when x"E2A9",
			x"0000" when x"E2AA",
			x"0000" when x"E2AB",
			x"0000" when x"E2AC",
			x"0000" when x"E2AD",
			x"0000" when x"E2AE",
			x"0000" when x"E2AF",
			x"0000" when x"E2B0",
			x"0000" when x"E2B1",
			x"0000" when x"E2B2",
			x"0000" when x"E2B3",
			x"0000" when x"E2B4",
			x"0000" when x"E2B5",
			x"0000" when x"E2B6",
			x"0000" when x"E2B7",
			x"0000" when x"E2B8",
			x"0000" when x"E2B9",
			x"0000" when x"E2BA",
			x"0000" when x"E2BB",
			x"0000" when x"E2BC",
			x"0000" when x"E2BD",
			x"0000" when x"E2BE",
			x"0000" when x"E2BF",
			x"0000" when x"E2C0",
			x"0000" when x"E2C1",
			x"0000" when x"E2C2",
			x"0000" when x"E2C3",
			x"0000" when x"E2C4",
			x"0000" when x"E2C5",
			x"0000" when x"E2C6",
			x"0000" when x"E2C7",
			x"0000" when x"E2C8",
			x"0000" when x"E2C9",
			x"0000" when x"E2CA",
			x"0000" when x"E2CB",
			x"0000" when x"E2CC",
			x"0000" when x"E2CD",
			x"0000" when x"E2CE",
			x"0000" when x"E2CF",
			x"0000" when x"E2D0",
			x"0000" when x"E2D1",
			x"0000" when x"E2D2",
			x"0000" when x"E2D3",
			x"0000" when x"E2D4",
			x"0000" when x"E2D5",
			x"0000" when x"E2D6",
			x"0000" when x"E2D7",
			x"0000" when x"E2D8",
			x"0000" when x"E2D9",
			x"0000" when x"E2DA",
			x"0000" when x"E2DB",
			x"0000" when x"E2DC",
			x"0000" when x"E2DD",
			x"0000" when x"E2DE",
			x"0000" when x"E2DF",
			x"0000" when x"E2E0",
			x"0000" when x"E2E1",
			x"0000" when x"E2E2",
			x"0000" when x"E2E3",
			x"0000" when x"E2E4",
			x"0000" when x"E2E5",
			x"0000" when x"E2E6",
			x"0000" when x"E2E7",
			x"0000" when x"E2E8",
			x"0000" when x"E2E9",
			x"0000" when x"E2EA",
			x"0000" when x"E2EB",
			x"0000" when x"E2EC",
			x"0000" when x"E2ED",
			x"0000" when x"E2EE",
			x"0000" when x"E2EF",
			x"0000" when x"E2F0",
			x"0000" when x"E2F1",
			x"0000" when x"E2F2",
			x"0000" when x"E2F3",
			x"0000" when x"E2F4",
			x"0000" when x"E2F5",
			x"0000" when x"E2F6",
			x"0000" when x"E2F7",
			x"0000" when x"E2F8",
			x"0000" when x"E2F9",
			x"0000" when x"E2FA",
			x"0000" when x"E2FB",
			x"0000" when x"E2FC",
			x"0000" when x"E2FD",
			x"0000" when x"E2FE",
			x"0000" when x"E2FF",
			x"0000" when x"E300",
			x"0000" when x"E301",
			x"0000" when x"E302",
			x"0000" when x"E303",
			x"0000" when x"E304",
			x"0000" when x"E305",
			x"0000" when x"E306",
			x"0000" when x"E307",
			x"0000" when x"E308",
			x"0000" when x"E309",
			x"0000" when x"E30A",
			x"0000" when x"E30B",
			x"0000" when x"E30C",
			x"0000" when x"E30D",
			x"0000" when x"E30E",
			x"0000" when x"E30F",
			x"0000" when x"E310",
			x"0000" when x"E311",
			x"0000" when x"E312",
			x"0000" when x"E313",
			x"0000" when x"E314",
			x"0000" when x"E315",
			x"0000" when x"E316",
			x"0000" when x"E317",
			x"0000" when x"E318",
			x"0000" when x"E319",
			x"0000" when x"E31A",
			x"0000" when x"E31B",
			x"0000" when x"E31C",
			x"0000" when x"E31D",
			x"0000" when x"E31E",
			x"0000" when x"E31F",
			x"0000" when x"E320",
			x"0000" when x"E321",
			x"0000" when x"E322",
			x"0000" when x"E323",
			x"0000" when x"E324",
			x"0000" when x"E325",
			x"0000" when x"E326",
			x"0000" when x"E327",
			x"0000" when x"E328",
			x"0000" when x"E329",
			x"0000" when x"E32A",
			x"0000" when x"E32B",
			x"0000" when x"E32C",
			x"0000" when x"E32D",
			x"0000" when x"E32E",
			x"0000" when x"E32F",
			x"0000" when x"E330",
			x"0000" when x"E331",
			x"0000" when x"E332",
			x"0000" when x"E333",
			x"0000" when x"E334",
			x"0000" when x"E335",
			x"0000" when x"E336",
			x"0000" when x"E337",
			x"0000" when x"E338",
			x"0000" when x"E339",
			x"0000" when x"E33A",
			x"0000" when x"E33B",
			x"0000" when x"E33C",
			x"0000" when x"E33D",
			x"0000" when x"E33E",
			x"0000" when x"E33F",
			x"0000" when x"E340",
			x"0000" when x"E341",
			x"0000" when x"E342",
			x"0000" when x"E343",
			x"0000" when x"E344",
			x"0000" when x"E345",
			x"0000" when x"E346",
			x"0000" when x"E347",
			x"0000" when x"E348",
			x"0000" when x"E349",
			x"0000" when x"E34A",
			x"0000" when x"E34B",
			x"0000" when x"E34C",
			x"0000" when x"E34D",
			x"0000" when x"E34E",
			x"0000" when x"E34F",
			x"0000" when x"E350",
			x"0000" when x"E351",
			x"0000" when x"E352",
			x"0000" when x"E353",
			x"0000" when x"E354",
			x"0000" when x"E355",
			x"0000" when x"E356",
			x"0000" when x"E357",
			x"0000" when x"E358",
			x"0000" when x"E359",
			x"0000" when x"E35A",
			x"0000" when x"E35B",
			x"0000" when x"E35C",
			x"0000" when x"E35D",
			x"0000" when x"E35E",
			x"0000" when x"E35F",
			x"0000" when x"E360",
			x"0000" when x"E361",
			x"0000" when x"E362",
			x"0000" when x"E363",
			x"0000" when x"E364",
			x"0000" when x"E365",
			x"0000" when x"E366",
			x"0000" when x"E367",
			x"0000" when x"E368",
			x"0000" when x"E369",
			x"0000" when x"E36A",
			x"0000" when x"E36B",
			x"0000" when x"E36C",
			x"0000" when x"E36D",
			x"0000" when x"E36E",
			x"0000" when x"E36F",
			x"0000" when x"E370",
			x"0000" when x"E371",
			x"0000" when x"E372",
			x"0000" when x"E373",
			x"0000" when x"E374",
			x"0000" when x"E375",
			x"0000" when x"E376",
			x"0000" when x"E377",
			x"0000" when x"E378",
			x"0000" when x"E379",
			x"0000" when x"E37A",
			x"0000" when x"E37B",
			x"0000" when x"E37C",
			x"0000" when x"E37D",
			x"0000" when x"E37E",
			x"0000" when x"E37F",
			x"0000" when x"E380",
			x"0000" when x"E381",
			x"0000" when x"E382",
			x"0000" when x"E383",
			x"0000" when x"E384",
			x"0000" when x"E385",
			x"0000" when x"E386",
			x"0000" when x"E387",
			x"0000" when x"E388",
			x"0000" when x"E389",
			x"0000" when x"E38A",
			x"0000" when x"E38B",
			x"0000" when x"E38C",
			x"0000" when x"E38D",
			x"0000" when x"E38E",
			x"0000" when x"E38F",
			x"0000" when x"E390",
			x"0000" when x"E391",
			x"0000" when x"E392",
			x"0000" when x"E393",
			x"0000" when x"E394",
			x"0000" when x"E395",
			x"0000" when x"E396",
			x"0000" when x"E397",
			x"0000" when x"E398",
			x"0000" when x"E399",
			x"0000" when x"E39A",
			x"0000" when x"E39B",
			x"0000" when x"E39C",
			x"0000" when x"E39D",
			x"0000" when x"E39E",
			x"0000" when x"E39F",
			x"0000" when x"E3A0",
			x"0000" when x"E3A1",
			x"0000" when x"E3A2",
			x"0000" when x"E3A3",
			x"0000" when x"E3A4",
			x"0000" when x"E3A5",
			x"0000" when x"E3A6",
			x"0000" when x"E3A7",
			x"0000" when x"E3A8",
			x"0000" when x"E3A9",
			x"0000" when x"E3AA",
			x"0000" when x"E3AB",
			x"0000" when x"E3AC",
			x"0000" when x"E3AD",
			x"0000" when x"E3AE",
			x"0000" when x"E3AF",
			x"0000" when x"E3B0",
			x"0000" when x"E3B1",
			x"0000" when x"E3B2",
			x"0000" when x"E3B3",
			x"0000" when x"E3B4",
			x"0000" when x"E3B5",
			x"0000" when x"E3B6",
			x"0000" when x"E3B7",
			x"0000" when x"E3B8",
			x"0000" when x"E3B9",
			x"0000" when x"E3BA",
			x"0000" when x"E3BB",
			x"0000" when x"E3BC",
			x"0000" when x"E3BD",
			x"0000" when x"E3BE",
			x"0000" when x"E3BF",
			x"0000" when x"E3C0",
			x"0000" when x"E3C1",
			x"0000" when x"E3C2",
			x"0000" when x"E3C3",
			x"0000" when x"E3C4",
			x"0000" when x"E3C5",
			x"0000" when x"E3C6",
			x"0000" when x"E3C7",
			x"0000" when x"E3C8",
			x"0000" when x"E3C9",
			x"0000" when x"E3CA",
			x"0000" when x"E3CB",
			x"0000" when x"E3CC",
			x"0000" when x"E3CD",
			x"0000" when x"E3CE",
			x"0000" when x"E3CF",
			x"0000" when x"E3D0",
			x"0000" when x"E3D1",
			x"0000" when x"E3D2",
			x"0000" when x"E3D3",
			x"0000" when x"E3D4",
			x"0000" when x"E3D5",
			x"0000" when x"E3D6",
			x"0000" when x"E3D7",
			x"0000" when x"E3D8",
			x"0000" when x"E3D9",
			x"0000" when x"E3DA",
			x"0000" when x"E3DB",
			x"0000" when x"E3DC",
			x"0000" when x"E3DD",
			x"0000" when x"E3DE",
			x"0000" when x"E3DF",
			x"0000" when x"E3E0",
			x"0000" when x"E3E1",
			x"0000" when x"E3E2",
			x"0000" when x"E3E3",
			x"0000" when x"E3E4",
			x"0000" when x"E3E5",
			x"0000" when x"E3E6",
			x"0000" when x"E3E7",
			x"0000" when x"E3E8",
			x"0000" when x"E3E9",
			x"0000" when x"E3EA",
			x"0000" when x"E3EB",
			x"0000" when x"E3EC",
			x"0000" when x"E3ED",
			x"0000" when x"E3EE",
			x"0000" when x"E3EF",
			x"0000" when x"E3F0",
			x"0000" when x"E3F1",
			x"0000" when x"E3F2",
			x"0000" when x"E3F3",
			x"0000" when x"E3F4",
			x"0000" when x"E3F5",
			x"0000" when x"E3F6",
			x"0000" when x"E3F7",
			x"0000" when x"E3F8",
			x"0000" when x"E3F9",
			x"0000" when x"E3FA",
			x"0000" when x"E3FB",
			x"0000" when x"E3FC",
			x"0000" when x"E3FD",
			x"0000" when x"E3FE",
			x"0000" when x"E3FF",
			x"0000" when x"E400",
			x"0000" when x"E401",
			x"0000" when x"E402",
			x"0000" when x"E403",
			x"0000" when x"E404",
			x"0000" when x"E405",
			x"0000" when x"E406",
			x"0000" when x"E407",
			x"0000" when x"E408",
			x"0000" when x"E409",
			x"0000" when x"E40A",
			x"0000" when x"E40B",
			x"0000" when x"E40C",
			x"0000" when x"E40D",
			x"0000" when x"E40E",
			x"0000" when x"E40F",
			x"0000" when x"E410",
			x"0000" when x"E411",
			x"0000" when x"E412",
			x"0000" when x"E413",
			x"0000" when x"E414",
			x"0000" when x"E415",
			x"0000" when x"E416",
			x"0000" when x"E417",
			x"0000" when x"E418",
			x"0000" when x"E419",
			x"0000" when x"E41A",
			x"0000" when x"E41B",
			x"0000" when x"E41C",
			x"0000" when x"E41D",
			x"0000" when x"E41E",
			x"0000" when x"E41F",
			x"0000" when x"E420",
			x"0000" when x"E421",
			x"0000" when x"E422",
			x"0000" when x"E423",
			x"0000" when x"E424",
			x"0000" when x"E425",
			x"0000" when x"E426",
			x"0000" when x"E427",
			x"0000" when x"E428",
			x"0000" when x"E429",
			x"0000" when x"E42A",
			x"0000" when x"E42B",
			x"0000" when x"E42C",
			x"0000" when x"E42D",
			x"0000" when x"E42E",
			x"0000" when x"E42F",
			x"0000" when x"E430",
			x"0000" when x"E431",
			x"0000" when x"E432",
			x"0000" when x"E433",
			x"0000" when x"E434",
			x"0000" when x"E435",
			x"0000" when x"E436",
			x"0000" when x"E437",
			x"0000" when x"E438",
			x"0000" when x"E439",
			x"0000" when x"E43A",
			x"0000" when x"E43B",
			x"0000" when x"E43C",
			x"0000" when x"E43D",
			x"0000" when x"E43E",
			x"0000" when x"E43F",
			x"0000" when x"E440",
			x"0000" when x"E441",
			x"0000" when x"E442",
			x"0000" when x"E443",
			x"0000" when x"E444",
			x"0000" when x"E445",
			x"0000" when x"E446",
			x"0000" when x"E447",
			x"0000" when x"E448",
			x"0000" when x"E449",
			x"0000" when x"E44A",
			x"0000" when x"E44B",
			x"0000" when x"E44C",
			x"0000" when x"E44D",
			x"0000" when x"E44E",
			x"0000" when x"E44F",
			x"0000" when x"E450",
			x"0000" when x"E451",
			x"0000" when x"E452",
			x"0000" when x"E453",
			x"0000" when x"E454",
			x"0000" when x"E455",
			x"0000" when x"E456",
			x"0000" when x"E457",
			x"0000" when x"E458",
			x"0000" when x"E459",
			x"0000" when x"E45A",
			x"0000" when x"E45B",
			x"0000" when x"E45C",
			x"0000" when x"E45D",
			x"0000" when x"E45E",
			x"0000" when x"E45F",
			x"0000" when x"E460",
			x"0000" when x"E461",
			x"0000" when x"E462",
			x"0000" when x"E463",
			x"0000" when x"E464",
			x"0000" when x"E465",
			x"0000" when x"E466",
			x"0000" when x"E467",
			x"0000" when x"E468",
			x"0000" when x"E469",
			x"0000" when x"E46A",
			x"0000" when x"E46B",
			x"0000" when x"E46C",
			x"0000" when x"E46D",
			x"0000" when x"E46E",
			x"0000" when x"E46F",
			x"0000" when x"E470",
			x"0000" when x"E471",
			x"0000" when x"E472",
			x"0000" when x"E473",
			x"0000" when x"E474",
			x"0000" when x"E475",
			x"0000" when x"E476",
			x"0000" when x"E477",
			x"0000" when x"E478",
			x"0000" when x"E479",
			x"0000" when x"E47A",
			x"0000" when x"E47B",
			x"0000" when x"E47C",
			x"0000" when x"E47D",
			x"0000" when x"E47E",
			x"0000" when x"E47F",
			x"0000" when x"E480",
			x"0000" when x"E481",
			x"0000" when x"E482",
			x"0000" when x"E483",
			x"0000" when x"E484",
			x"0000" when x"E485",
			x"0000" when x"E486",
			x"0000" when x"E487",
			x"0000" when x"E488",
			x"0000" when x"E489",
			x"0000" when x"E48A",
			x"0000" when x"E48B",
			x"0000" when x"E48C",
			x"0000" when x"E48D",
			x"0000" when x"E48E",
			x"0000" when x"E48F",
			x"0000" when x"E490",
			x"0000" when x"E491",
			x"0000" when x"E492",
			x"0000" when x"E493",
			x"0000" when x"E494",
			x"0000" when x"E495",
			x"0000" when x"E496",
			x"0000" when x"E497",
			x"0000" when x"E498",
			x"0000" when x"E499",
			x"0000" when x"E49A",
			x"0000" when x"E49B",
			x"0000" when x"E49C",
			x"0000" when x"E49D",
			x"0000" when x"E49E",
			x"0000" when x"E49F",
			x"0000" when x"E4A0",
			x"0000" when x"E4A1",
			x"0000" when x"E4A2",
			x"0000" when x"E4A3",
			x"0000" when x"E4A4",
			x"0000" when x"E4A5",
			x"0000" when x"E4A6",
			x"0000" when x"E4A7",
			x"0000" when x"E4A8",
			x"0000" when x"E4A9",
			x"0000" when x"E4AA",
			x"0000" when x"E4AB",
			x"0000" when x"E4AC",
			x"0000" when x"E4AD",
			x"0000" when x"E4AE",
			x"0000" when x"E4AF",
			x"0000" when x"E4B0",
			x"0000" when x"E4B1",
			x"0000" when x"E4B2",
			x"0000" when x"E4B3",
			x"0000" when x"E4B4",
			x"0000" when x"E4B5",
			x"0000" when x"E4B6",
			x"0000" when x"E4B7",
			x"0000" when x"E4B8",
			x"0000" when x"E4B9",
			x"0000" when x"E4BA",
			x"0000" when x"E4BB",
			x"0000" when x"E4BC",
			x"0000" when x"E4BD",
			x"0000" when x"E4BE",
			x"0000" when x"E4BF",
			x"0000" when x"E4C0",
			x"0000" when x"E4C1",
			x"0000" when x"E4C2",
			x"0000" when x"E4C3",
			x"0000" when x"E4C4",
			x"0000" when x"E4C5",
			x"0000" when x"E4C6",
			x"0000" when x"E4C7",
			x"0000" when x"E4C8",
			x"0000" when x"E4C9",
			x"0000" when x"E4CA",
			x"0000" when x"E4CB",
			x"0000" when x"E4CC",
			x"0000" when x"E4CD",
			x"0000" when x"E4CE",
			x"0000" when x"E4CF",
			x"0000" when x"E4D0",
			x"0000" when x"E4D1",
			x"0000" when x"E4D2",
			x"0000" when x"E4D3",
			x"0000" when x"E4D4",
			x"0000" when x"E4D5",
			x"0000" when x"E4D6",
			x"0000" when x"E4D7",
			x"0000" when x"E4D8",
			x"0000" when x"E4D9",
			x"0000" when x"E4DA",
			x"0000" when x"E4DB",
			x"0000" when x"E4DC",
			x"0000" when x"E4DD",
			x"0000" when x"E4DE",
			x"0000" when x"E4DF",
			x"0000" when x"E4E0",
			x"0000" when x"E4E1",
			x"0000" when x"E4E2",
			x"0000" when x"E4E3",
			x"0000" when x"E4E4",
			x"0000" when x"E4E5",
			x"0000" when x"E4E6",
			x"0000" when x"E4E7",
			x"0000" when x"E4E8",
			x"0000" when x"E4E9",
			x"0000" when x"E4EA",
			x"0000" when x"E4EB",
			x"0000" when x"E4EC",
			x"0000" when x"E4ED",
			x"0000" when x"E4EE",
			x"0000" when x"E4EF",
			x"0000" when x"E4F0",
			x"0000" when x"E4F1",
			x"0000" when x"E4F2",
			x"0000" when x"E4F3",
			x"0000" when x"E4F4",
			x"0000" when x"E4F5",
			x"0000" when x"E4F6",
			x"0000" when x"E4F7",
			x"0000" when x"E4F8",
			x"0000" when x"E4F9",
			x"0000" when x"E4FA",
			x"0000" when x"E4FB",
			x"0000" when x"E4FC",
			x"0000" when x"E4FD",
			x"0000" when x"E4FE",
			x"0000" when x"E4FF",
			x"0000" when x"E500",
			x"0000" when x"E501",
			x"0000" when x"E502",
			x"0000" when x"E503",
			x"0000" when x"E504",
			x"0000" when x"E505",
			x"0000" when x"E506",
			x"0000" when x"E507",
			x"0000" when x"E508",
			x"0000" when x"E509",
			x"0000" when x"E50A",
			x"0000" when x"E50B",
			x"0000" when x"E50C",
			x"0000" when x"E50D",
			x"0000" when x"E50E",
			x"0000" when x"E50F",
			x"0000" when x"E510",
			x"0000" when x"E511",
			x"0000" when x"E512",
			x"0000" when x"E513",
			x"0000" when x"E514",
			x"0000" when x"E515",
			x"0000" when x"E516",
			x"0000" when x"E517",
			x"0000" when x"E518",
			x"0000" when x"E519",
			x"0000" when x"E51A",
			x"0000" when x"E51B",
			x"0000" when x"E51C",
			x"0000" when x"E51D",
			x"0000" when x"E51E",
			x"0000" when x"E51F",
			x"0000" when x"E520",
			x"0000" when x"E521",
			x"0000" when x"E522",
			x"0000" when x"E523",
			x"0000" when x"E524",
			x"0000" when x"E525",
			x"0000" when x"E526",
			x"0000" when x"E527",
			x"0000" when x"E528",
			x"0000" when x"E529",
			x"0000" when x"E52A",
			x"0000" when x"E52B",
			x"0000" when x"E52C",
			x"0000" when x"E52D",
			x"0000" when x"E52E",
			x"0000" when x"E52F",
			x"0000" when x"E530",
			x"0000" when x"E531",
			x"0000" when x"E532",
			x"0000" when x"E533",
			x"0000" when x"E534",
			x"0000" when x"E535",
			x"0000" when x"E536",
			x"0000" when x"E537",
			x"0000" when x"E538",
			x"0000" when x"E539",
			x"0000" when x"E53A",
			x"0000" when x"E53B",
			x"0000" when x"E53C",
			x"0000" when x"E53D",
			x"0000" when x"E53E",
			x"0000" when x"E53F",
			x"0000" when x"E540",
			x"0000" when x"E541",
			x"0000" when x"E542",
			x"0000" when x"E543",
			x"0000" when x"E544",
			x"0000" when x"E545",
			x"0000" when x"E546",
			x"0000" when x"E547",
			x"0000" when x"E548",
			x"0000" when x"E549",
			x"0000" when x"E54A",
			x"0000" when x"E54B",
			x"0000" when x"E54C",
			x"0000" when x"E54D",
			x"0000" when x"E54E",
			x"0000" when x"E54F",
			x"0000" when x"E550",
			x"0000" when x"E551",
			x"0000" when x"E552",
			x"0000" when x"E553",
			x"0000" when x"E554",
			x"0000" when x"E555",
			x"0000" when x"E556",
			x"0000" when x"E557",
			x"0000" when x"E558",
			x"0000" when x"E559",
			x"0000" when x"E55A",
			x"0000" when x"E55B",
			x"0000" when x"E55C",
			x"0000" when x"E55D",
			x"0000" when x"E55E",
			x"0000" when x"E55F",
			x"0000" when x"E560",
			x"0000" when x"E561",
			x"0000" when x"E562",
			x"0000" when x"E563",
			x"0000" when x"E564",
			x"0000" when x"E565",
			x"0000" when x"E566",
			x"0000" when x"E567",
			x"0000" when x"E568",
			x"0000" when x"E569",
			x"0000" when x"E56A",
			x"0000" when x"E56B",
			x"0000" when x"E56C",
			x"0000" when x"E56D",
			x"0000" when x"E56E",
			x"0000" when x"E56F",
			x"0000" when x"E570",
			x"0000" when x"E571",
			x"0000" when x"E572",
			x"0000" when x"E573",
			x"0000" when x"E574",
			x"0000" when x"E575",
			x"0000" when x"E576",
			x"0000" when x"E577",
			x"0000" when x"E578",
			x"0000" when x"E579",
			x"0000" when x"E57A",
			x"0000" when x"E57B",
			x"0000" when x"E57C",
			x"0000" when x"E57D",
			x"0000" when x"E57E",
			x"0000" when x"E57F",
			x"0000" when x"E580",
			x"0000" when x"E581",
			x"0000" when x"E582",
			x"0000" when x"E583",
			x"0000" when x"E584",
			x"0000" when x"E585",
			x"0000" when x"E586",
			x"0000" when x"E587",
			x"0000" when x"E588",
			x"0000" when x"E589",
			x"0000" when x"E58A",
			x"0000" when x"E58B",
			x"0000" when x"E58C",
			x"0000" when x"E58D",
			x"0000" when x"E58E",
			x"0000" when x"E58F",
			x"0000" when x"E590",
			x"0000" when x"E591",
			x"0000" when x"E592",
			x"0000" when x"E593",
			x"0000" when x"E594",
			x"0000" when x"E595",
			x"0000" when x"E596",
			x"0000" when x"E597",
			x"0000" when x"E598",
			x"0000" when x"E599",
			x"0000" when x"E59A",
			x"0000" when x"E59B",
			x"0000" when x"E59C",
			x"0000" when x"E59D",
			x"0000" when x"E59E",
			x"0000" when x"E59F",
			x"0000" when x"E5A0",
			x"0000" when x"E5A1",
			x"0000" when x"E5A2",
			x"0000" when x"E5A3",
			x"0000" when x"E5A4",
			x"0000" when x"E5A5",
			x"0000" when x"E5A6",
			x"0000" when x"E5A7",
			x"0000" when x"E5A8",
			x"0000" when x"E5A9",
			x"0000" when x"E5AA",
			x"0000" when x"E5AB",
			x"0000" when x"E5AC",
			x"0000" when x"E5AD",
			x"0000" when x"E5AE",
			x"0000" when x"E5AF",
			x"0000" when x"E5B0",
			x"0000" when x"E5B1",
			x"0000" when x"E5B2",
			x"0000" when x"E5B3",
			x"0000" when x"E5B4",
			x"0000" when x"E5B5",
			x"0000" when x"E5B6",
			x"0000" when x"E5B7",
			x"0000" when x"E5B8",
			x"0000" when x"E5B9",
			x"0000" when x"E5BA",
			x"0000" when x"E5BB",
			x"0000" when x"E5BC",
			x"0000" when x"E5BD",
			x"0000" when x"E5BE",
			x"0000" when x"E5BF",
			x"0000" when x"E5C0",
			x"0000" when x"E5C1",
			x"0000" when x"E5C2",
			x"0000" when x"E5C3",
			x"0000" when x"E5C4",
			x"0000" when x"E5C5",
			x"0000" when x"E5C6",
			x"0000" when x"E5C7",
			x"0000" when x"E5C8",
			x"0000" when x"E5C9",
			x"0000" when x"E5CA",
			x"0000" when x"E5CB",
			x"0000" when x"E5CC",
			x"0000" when x"E5CD",
			x"0000" when x"E5CE",
			x"0000" when x"E5CF",
			x"0000" when x"E5D0",
			x"0000" when x"E5D1",
			x"0000" when x"E5D2",
			x"0000" when x"E5D3",
			x"0000" when x"E5D4",
			x"0000" when x"E5D5",
			x"0000" when x"E5D6",
			x"0000" when x"E5D7",
			x"0000" when x"E5D8",
			x"0000" when x"E5D9",
			x"0000" when x"E5DA",
			x"0000" when x"E5DB",
			x"0000" when x"E5DC",
			x"0000" when x"E5DD",
			x"0000" when x"E5DE",
			x"0000" when x"E5DF",
			x"0000" when x"E5E0",
			x"0000" when x"E5E1",
			x"0000" when x"E5E2",
			x"0000" when x"E5E3",
			x"0000" when x"E5E4",
			x"0000" when x"E5E5",
			x"0000" when x"E5E6",
			x"0000" when x"E5E7",
			x"0000" when x"E5E8",
			x"0000" when x"E5E9",
			x"0000" when x"E5EA",
			x"0000" when x"E5EB",
			x"0000" when x"E5EC",
			x"0000" when x"E5ED",
			x"0000" when x"E5EE",
			x"0000" when x"E5EF",
			x"0000" when x"E5F0",
			x"0000" when x"E5F1",
			x"0000" when x"E5F2",
			x"0000" when x"E5F3",
			x"0000" when x"E5F4",
			x"0000" when x"E5F5",
			x"0000" when x"E5F6",
			x"0000" when x"E5F7",
			x"0000" when x"E5F8",
			x"0000" when x"E5F9",
			x"0000" when x"E5FA",
			x"0000" when x"E5FB",
			x"0000" when x"E5FC",
			x"0000" when x"E5FD",
			x"0000" when x"E5FE",
			x"0000" when x"E5FF",
			x"0000" when x"E600",
			x"0000" when x"E601",
			x"0000" when x"E602",
			x"0000" when x"E603",
			x"0000" when x"E604",
			x"0000" when x"E605",
			x"0000" when x"E606",
			x"0000" when x"E607",
			x"0000" when x"E608",
			x"0000" when x"E609",
			x"0000" when x"E60A",
			x"0000" when x"E60B",
			x"0000" when x"E60C",
			x"0000" when x"E60D",
			x"0000" when x"E60E",
			x"0000" when x"E60F",
			x"0000" when x"E610",
			x"0000" when x"E611",
			x"0000" when x"E612",
			x"0000" when x"E613",
			x"0000" when x"E614",
			x"0000" when x"E615",
			x"0000" when x"E616",
			x"0000" when x"E617",
			x"0000" when x"E618",
			x"0000" when x"E619",
			x"0000" when x"E61A",
			x"0000" when x"E61B",
			x"0000" when x"E61C",
			x"0000" when x"E61D",
			x"0000" when x"E61E",
			x"0000" when x"E61F",
			x"0000" when x"E620",
			x"0000" when x"E621",
			x"0000" when x"E622",
			x"0000" when x"E623",
			x"0000" when x"E624",
			x"0000" when x"E625",
			x"0000" when x"E626",
			x"0000" when x"E627",
			x"0000" when x"E628",
			x"0000" when x"E629",
			x"0000" when x"E62A",
			x"0000" when x"E62B",
			x"0000" when x"E62C",
			x"0000" when x"E62D",
			x"0000" when x"E62E",
			x"0000" when x"E62F",
			x"0000" when x"E630",
			x"0000" when x"E631",
			x"0000" when x"E632",
			x"0000" when x"E633",
			x"0000" when x"E634",
			x"0000" when x"E635",
			x"0000" when x"E636",
			x"0000" when x"E637",
			x"0000" when x"E638",
			x"0000" when x"E639",
			x"0000" when x"E63A",
			x"0000" when x"E63B",
			x"0000" when x"E63C",
			x"0000" when x"E63D",
			x"0000" when x"E63E",
			x"0000" when x"E63F",
			x"0000" when x"E640",
			x"0000" when x"E641",
			x"0000" when x"E642",
			x"0000" when x"E643",
			x"0000" when x"E644",
			x"0000" when x"E645",
			x"0000" when x"E646",
			x"0000" when x"E647",
			x"0000" when x"E648",
			x"0000" when x"E649",
			x"0000" when x"E64A",
			x"0000" when x"E64B",
			x"0000" when x"E64C",
			x"0000" when x"E64D",
			x"0000" when x"E64E",
			x"0000" when x"E64F",
			x"0000" when x"E650",
			x"0000" when x"E651",
			x"0000" when x"E652",
			x"0000" when x"E653",
			x"0000" when x"E654",
			x"0000" when x"E655",
			x"0000" when x"E656",
			x"0000" when x"E657",
			x"0000" when x"E658",
			x"0000" when x"E659",
			x"0000" when x"E65A",
			x"0000" when x"E65B",
			x"0000" when x"E65C",
			x"0000" when x"E65D",
			x"0000" when x"E65E",
			x"0000" when x"E65F",
			x"0000" when x"E660",
			x"0000" when x"E661",
			x"0000" when x"E662",
			x"0000" when x"E663",
			x"0000" when x"E664",
			x"0000" when x"E665",
			x"0000" when x"E666",
			x"0000" when x"E667",
			x"0000" when x"E668",
			x"0000" when x"E669",
			x"0000" when x"E66A",
			x"0000" when x"E66B",
			x"0000" when x"E66C",
			x"0000" when x"E66D",
			x"0000" when x"E66E",
			x"0000" when x"E66F",
			x"0000" when x"E670",
			x"0000" when x"E671",
			x"0000" when x"E672",
			x"0000" when x"E673",
			x"0000" when x"E674",
			x"0000" when x"E675",
			x"0000" when x"E676",
			x"0000" when x"E677",
			x"0000" when x"E678",
			x"0000" when x"E679",
			x"0000" when x"E67A",
			x"0000" when x"E67B",
			x"0000" when x"E67C",
			x"0000" when x"E67D",
			x"0000" when x"E67E",
			x"0000" when x"E67F",
			x"0000" when x"E680",
			x"0000" when x"E681",
			x"0000" when x"E682",
			x"0000" when x"E683",
			x"0000" when x"E684",
			x"0000" when x"E685",
			x"0000" when x"E686",
			x"0000" when x"E687",
			x"0000" when x"E688",
			x"0000" when x"E689",
			x"0000" when x"E68A",
			x"0000" when x"E68B",
			x"0000" when x"E68C",
			x"0000" when x"E68D",
			x"0000" when x"E68E",
			x"0000" when x"E68F",
			x"0000" when x"E690",
			x"0000" when x"E691",
			x"0000" when x"E692",
			x"0000" when x"E693",
			x"0000" when x"E694",
			x"0000" when x"E695",
			x"0000" when x"E696",
			x"0000" when x"E697",
			x"0000" when x"E698",
			x"0000" when x"E699",
			x"0000" when x"E69A",
			x"0000" when x"E69B",
			x"0000" when x"E69C",
			x"0000" when x"E69D",
			x"0000" when x"E69E",
			x"0000" when x"E69F",
			x"0000" when x"E6A0",
			x"0000" when x"E6A1",
			x"0000" when x"E6A2",
			x"0000" when x"E6A3",
			x"0000" when x"E6A4",
			x"0000" when x"E6A5",
			x"0000" when x"E6A6",
			x"0000" when x"E6A7",
			x"0000" when x"E6A8",
			x"0000" when x"E6A9",
			x"0000" when x"E6AA",
			x"0000" when x"E6AB",
			x"0000" when x"E6AC",
			x"0000" when x"E6AD",
			x"0000" when x"E6AE",
			x"0000" when x"E6AF",
			x"0000" when x"E6B0",
			x"0000" when x"E6B1",
			x"0000" when x"E6B2",
			x"0000" when x"E6B3",
			x"0000" when x"E6B4",
			x"0000" when x"E6B5",
			x"0000" when x"E6B6",
			x"0000" when x"E6B7",
			x"0000" when x"E6B8",
			x"0000" when x"E6B9",
			x"0000" when x"E6BA",
			x"0000" when x"E6BB",
			x"0000" when x"E6BC",
			x"0000" when x"E6BD",
			x"0000" when x"E6BE",
			x"0000" when x"E6BF",
			x"0000" when x"E6C0",
			x"0000" when x"E6C1",
			x"0000" when x"E6C2",
			x"0000" when x"E6C3",
			x"0000" when x"E6C4",
			x"0000" when x"E6C5",
			x"0000" when x"E6C6",
			x"0000" when x"E6C7",
			x"0000" when x"E6C8",
			x"0000" when x"E6C9",
			x"0000" when x"E6CA",
			x"0000" when x"E6CB",
			x"0000" when x"E6CC",
			x"0000" when x"E6CD",
			x"0000" when x"E6CE",
			x"0000" when x"E6CF",
			x"0000" when x"E6D0",
			x"0000" when x"E6D1",
			x"0000" when x"E6D2",
			x"0000" when x"E6D3",
			x"0000" when x"E6D4",
			x"0000" when x"E6D5",
			x"0000" when x"E6D6",
			x"0000" when x"E6D7",
			x"0000" when x"E6D8",
			x"0000" when x"E6D9",
			x"0000" when x"E6DA",
			x"0000" when x"E6DB",
			x"0000" when x"E6DC",
			x"0000" when x"E6DD",
			x"0000" when x"E6DE",
			x"0000" when x"E6DF",
			x"0000" when x"E6E0",
			x"0000" when x"E6E1",
			x"0000" when x"E6E2",
			x"0000" when x"E6E3",
			x"0000" when x"E6E4",
			x"0000" when x"E6E5",
			x"0000" when x"E6E6",
			x"0000" when x"E6E7",
			x"0000" when x"E6E8",
			x"0000" when x"E6E9",
			x"0000" when x"E6EA",
			x"0000" when x"E6EB",
			x"0000" when x"E6EC",
			x"0000" when x"E6ED",
			x"0000" when x"E6EE",
			x"0000" when x"E6EF",
			x"0000" when x"E6F0",
			x"0000" when x"E6F1",
			x"0000" when x"E6F2",
			x"0000" when x"E6F3",
			x"0000" when x"E6F4",
			x"0000" when x"E6F5",
			x"0000" when x"E6F6",
			x"0000" when x"E6F7",
			x"0000" when x"E6F8",
			x"0000" when x"E6F9",
			x"0000" when x"E6FA",
			x"0000" when x"E6FB",
			x"0000" when x"E6FC",
			x"0000" when x"E6FD",
			x"0000" when x"E6FE",
			x"0000" when x"E6FF",
			x"0000" when x"E700",
			x"0000" when x"E701",
			x"0000" when x"E702",
			x"0000" when x"E703",
			x"0000" when x"E704",
			x"0000" when x"E705",
			x"0000" when x"E706",
			x"0000" when x"E707",
			x"0000" when x"E708",
			x"0000" when x"E709",
			x"0000" when x"E70A",
			x"0000" when x"E70B",
			x"0000" when x"E70C",
			x"0000" when x"E70D",
			x"0000" when x"E70E",
			x"0000" when x"E70F",
			x"0000" when x"E710",
			x"0000" when x"E711",
			x"0000" when x"E712",
			x"0000" when x"E713",
			x"0000" when x"E714",
			x"0000" when x"E715",
			x"0000" when x"E716",
			x"0000" when x"E717",
			x"0000" when x"E718",
			x"0000" when x"E719",
			x"0000" when x"E71A",
			x"0000" when x"E71B",
			x"0000" when x"E71C",
			x"0000" when x"E71D",
			x"0000" when x"E71E",
			x"0000" when x"E71F",
			x"0000" when x"E720",
			x"0000" when x"E721",
			x"0000" when x"E722",
			x"0000" when x"E723",
			x"0000" when x"E724",
			x"0000" when x"E725",
			x"0000" when x"E726",
			x"0000" when x"E727",
			x"0000" when x"E728",
			x"0000" when x"E729",
			x"0000" when x"E72A",
			x"0000" when x"E72B",
			x"0000" when x"E72C",
			x"0000" when x"E72D",
			x"0000" when x"E72E",
			x"0000" when x"E72F",
			x"0000" when x"E730",
			x"0000" when x"E731",
			x"0000" when x"E732",
			x"0000" when x"E733",
			x"0000" when x"E734",
			x"0000" when x"E735",
			x"0000" when x"E736",
			x"0000" when x"E737",
			x"0000" when x"E738",
			x"0000" when x"E739",
			x"0000" when x"E73A",
			x"0000" when x"E73B",
			x"0000" when x"E73C",
			x"0000" when x"E73D",
			x"0000" when x"E73E",
			x"0000" when x"E73F",
			x"0000" when x"E740",
			x"0000" when x"E741",
			x"0000" when x"E742",
			x"0000" when x"E743",
			x"0000" when x"E744",
			x"0000" when x"E745",
			x"0000" when x"E746",
			x"0000" when x"E747",
			x"0000" when x"E748",
			x"0000" when x"E749",
			x"0000" when x"E74A",
			x"0000" when x"E74B",
			x"0000" when x"E74C",
			x"0000" when x"E74D",
			x"0000" when x"E74E",
			x"0000" when x"E74F",
			x"0000" when x"E750",
			x"0000" when x"E751",
			x"0000" when x"E752",
			x"0000" when x"E753",
			x"0000" when x"E754",
			x"0000" when x"E755",
			x"0000" when x"E756",
			x"0000" when x"E757",
			x"0000" when x"E758",
			x"0000" when x"E759",
			x"0000" when x"E75A",
			x"0000" when x"E75B",
			x"0000" when x"E75C",
			x"0000" when x"E75D",
			x"0000" when x"E75E",
			x"0000" when x"E75F",
			x"0000" when x"E760",
			x"0000" when x"E761",
			x"0000" when x"E762",
			x"0000" when x"E763",
			x"0000" when x"E764",
			x"0000" when x"E765",
			x"0000" when x"E766",
			x"0000" when x"E767",
			x"0000" when x"E768",
			x"0000" when x"E769",
			x"0000" when x"E76A",
			x"0000" when x"E76B",
			x"0000" when x"E76C",
			x"0000" when x"E76D",
			x"0000" when x"E76E",
			x"0000" when x"E76F",
			x"0000" when x"E770",
			x"0000" when x"E771",
			x"0000" when x"E772",
			x"0000" when x"E773",
			x"0000" when x"E774",
			x"0000" when x"E775",
			x"0000" when x"E776",
			x"0000" when x"E777",
			x"0000" when x"E778",
			x"0000" when x"E779",
			x"0000" when x"E77A",
			x"0000" when x"E77B",
			x"0000" when x"E77C",
			x"0000" when x"E77D",
			x"0000" when x"E77E",
			x"0000" when x"E77F",
			x"0000" when x"E780",
			x"0000" when x"E781",
			x"0000" when x"E782",
			x"0000" when x"E783",
			x"0000" when x"E784",
			x"0000" when x"E785",
			x"0000" when x"E786",
			x"0000" when x"E787",
			x"0000" when x"E788",
			x"0000" when x"E789",
			x"0000" when x"E78A",
			x"0000" when x"E78B",
			x"0000" when x"E78C",
			x"0000" when x"E78D",
			x"0000" when x"E78E",
			x"0000" when x"E78F",
			x"0000" when x"E790",
			x"0000" when x"E791",
			x"0000" when x"E792",
			x"0000" when x"E793",
			x"0000" when x"E794",
			x"0000" when x"E795",
			x"0000" when x"E796",
			x"0000" when x"E797",
			x"0000" when x"E798",
			x"0000" when x"E799",
			x"0000" when x"E79A",
			x"0000" when x"E79B",
			x"0000" when x"E79C",
			x"0000" when x"E79D",
			x"0000" when x"E79E",
			x"0000" when x"E79F",
			x"0000" when x"E7A0",
			x"0000" when x"E7A1",
			x"0000" when x"E7A2",
			x"0000" when x"E7A3",
			x"0000" when x"E7A4",
			x"0000" when x"E7A5",
			x"0000" when x"E7A6",
			x"0000" when x"E7A7",
			x"0000" when x"E7A8",
			x"0000" when x"E7A9",
			x"0000" when x"E7AA",
			x"0000" when x"E7AB",
			x"0000" when x"E7AC",
			x"0000" when x"E7AD",
			x"0000" when x"E7AE",
			x"0000" when x"E7AF",
			x"0000" when x"E7B0",
			x"0000" when x"E7B1",
			x"0000" when x"E7B2",
			x"0000" when x"E7B3",
			x"0000" when x"E7B4",
			x"0000" when x"E7B5",
			x"0000" when x"E7B6",
			x"0000" when x"E7B7",
			x"0000" when x"E7B8",
			x"0000" when x"E7B9",
			x"0000" when x"E7BA",
			x"0000" when x"E7BB",
			x"0000" when x"E7BC",
			x"0000" when x"E7BD",
			x"0000" when x"E7BE",
			x"0000" when x"E7BF",
			x"0000" when x"E7C0",
			x"0000" when x"E7C1",
			x"0000" when x"E7C2",
			x"0000" when x"E7C3",
			x"0000" when x"E7C4",
			x"0000" when x"E7C5",
			x"0000" when x"E7C6",
			x"0000" when x"E7C7",
			x"0000" when x"E7C8",
			x"0000" when x"E7C9",
			x"0000" when x"E7CA",
			x"0000" when x"E7CB",
			x"0000" when x"E7CC",
			x"0000" when x"E7CD",
			x"0000" when x"E7CE",
			x"0000" when x"E7CF",
			x"0000" when x"E7D0",
			x"0000" when x"E7D1",
			x"0000" when x"E7D2",
			x"0000" when x"E7D3",
			x"0000" when x"E7D4",
			x"0000" when x"E7D5",
			x"0000" when x"E7D6",
			x"0000" when x"E7D7",
			x"0000" when x"E7D8",
			x"0000" when x"E7D9",
			x"0000" when x"E7DA",
			x"0000" when x"E7DB",
			x"0000" when x"E7DC",
			x"0000" when x"E7DD",
			x"0000" when x"E7DE",
			x"0000" when x"E7DF",
			x"0000" when x"E7E0",
			x"0000" when x"E7E1",
			x"0000" when x"E7E2",
			x"0000" when x"E7E3",
			x"0000" when x"E7E4",
			x"0000" when x"E7E5",
			x"0000" when x"E7E6",
			x"0000" when x"E7E7",
			x"0000" when x"E7E8",
			x"0000" when x"E7E9",
			x"0000" when x"E7EA",
			x"0000" when x"E7EB",
			x"0000" when x"E7EC",
			x"0000" when x"E7ED",
			x"0000" when x"E7EE",
			x"0000" when x"E7EF",
			x"0000" when x"E7F0",
			x"0000" when x"E7F1",
			x"0000" when x"E7F2",
			x"0000" when x"E7F3",
			x"0000" when x"E7F4",
			x"0000" when x"E7F5",
			x"0000" when x"E7F6",
			x"0000" when x"E7F7",
			x"0000" when x"E7F8",
			x"0000" when x"E7F9",
			x"0000" when x"E7FA",
			x"0000" when x"E7FB",
			x"0000" when x"E7FC",
			x"0000" when x"E7FD",
			x"0000" when x"E7FE",
			x"0000" when x"E7FF",
			x"0000" when x"E800",
			x"0000" when x"E801",
			x"0000" when x"E802",
			x"0000" when x"E803",
			x"0000" when x"E804",
			x"0000" when x"E805",
			x"0000" when x"E806",
			x"0000" when x"E807",
			x"0000" when x"E808",
			x"0000" when x"E809",
			x"0000" when x"E80A",
			x"0000" when x"E80B",
			x"0000" when x"E80C",
			x"0000" when x"E80D",
			x"0000" when x"E80E",
			x"0000" when x"E80F",
			x"0000" when x"E810",
			x"0000" when x"E811",
			x"0000" when x"E812",
			x"0000" when x"E813",
			x"0000" when x"E814",
			x"0000" when x"E815",
			x"0000" when x"E816",
			x"0000" when x"E817",
			x"0000" when x"E818",
			x"0000" when x"E819",
			x"0000" when x"E81A",
			x"0000" when x"E81B",
			x"0000" when x"E81C",
			x"0000" when x"E81D",
			x"0000" when x"E81E",
			x"0000" when x"E81F",
			x"0000" when x"E820",
			x"0000" when x"E821",
			x"0000" when x"E822",
			x"0000" when x"E823",
			x"0000" when x"E824",
			x"0000" when x"E825",
			x"0000" when x"E826",
			x"0000" when x"E827",
			x"0000" when x"E828",
			x"0000" when x"E829",
			x"0000" when x"E82A",
			x"0000" when x"E82B",
			x"0000" when x"E82C",
			x"0000" when x"E82D",
			x"0000" when x"E82E",
			x"0000" when x"E82F",
			x"0000" when x"E830",
			x"0000" when x"E831",
			x"0000" when x"E832",
			x"0000" when x"E833",
			x"0000" when x"E834",
			x"0000" when x"E835",
			x"0000" when x"E836",
			x"0000" when x"E837",
			x"0000" when x"E838",
			x"0000" when x"E839",
			x"0000" when x"E83A",
			x"0000" when x"E83B",
			x"0000" when x"E83C",
			x"0000" when x"E83D",
			x"0000" when x"E83E",
			x"0000" when x"E83F",
			x"0000" when x"E840",
			x"0000" when x"E841",
			x"0000" when x"E842",
			x"0000" when x"E843",
			x"0000" when x"E844",
			x"0000" when x"E845",
			x"0000" when x"E846",
			x"0000" when x"E847",
			x"0000" when x"E848",
			x"0000" when x"E849",
			x"0000" when x"E84A",
			x"0000" when x"E84B",
			x"0000" when x"E84C",
			x"0000" when x"E84D",
			x"0000" when x"E84E",
			x"0000" when x"E84F",
			x"0000" when x"E850",
			x"0000" when x"E851",
			x"0000" when x"E852",
			x"0000" when x"E853",
			x"0000" when x"E854",
			x"0000" when x"E855",
			x"0000" when x"E856",
			x"0000" when x"E857",
			x"0000" when x"E858",
			x"0000" when x"E859",
			x"0000" when x"E85A",
			x"0000" when x"E85B",
			x"0000" when x"E85C",
			x"0000" when x"E85D",
			x"0000" when x"E85E",
			x"0000" when x"E85F",
			x"0000" when x"E860",
			x"0000" when x"E861",
			x"0000" when x"E862",
			x"0000" when x"E863",
			x"0000" when x"E864",
			x"0000" when x"E865",
			x"0000" when x"E866",
			x"0000" when x"E867",
			x"0000" when x"E868",
			x"0000" when x"E869",
			x"0000" when x"E86A",
			x"0000" when x"E86B",
			x"0000" when x"E86C",
			x"0000" when x"E86D",
			x"0000" when x"E86E",
			x"0000" when x"E86F",
			x"0000" when x"E870",
			x"0000" when x"E871",
			x"0000" when x"E872",
			x"0000" when x"E873",
			x"0000" when x"E874",
			x"0000" when x"E875",
			x"0000" when x"E876",
			x"0000" when x"E877",
			x"0000" when x"E878",
			x"0000" when x"E879",
			x"0000" when x"E87A",
			x"0000" when x"E87B",
			x"0000" when x"E87C",
			x"0000" when x"E87D",
			x"0000" when x"E87E",
			x"0000" when x"E87F",
			x"0000" when x"E880",
			x"0000" when x"E881",
			x"0000" when x"E882",
			x"0000" when x"E883",
			x"0000" when x"E884",
			x"0000" when x"E885",
			x"0000" when x"E886",
			x"0000" when x"E887",
			x"0000" when x"E888",
			x"0000" when x"E889",
			x"0000" when x"E88A",
			x"0000" when x"E88B",
			x"0000" when x"E88C",
			x"0000" when x"E88D",
			x"0000" when x"E88E",
			x"0000" when x"E88F",
			x"0000" when x"E890",
			x"0000" when x"E891",
			x"0000" when x"E892",
			x"0000" when x"E893",
			x"0000" when x"E894",
			x"0000" when x"E895",
			x"0000" when x"E896",
			x"0000" when x"E897",
			x"0000" when x"E898",
			x"0000" when x"E899",
			x"0000" when x"E89A",
			x"0000" when x"E89B",
			x"0000" when x"E89C",
			x"0000" when x"E89D",
			x"0000" when x"E89E",
			x"0000" when x"E89F",
			x"0000" when x"E8A0",
			x"0000" when x"E8A1",
			x"0000" when x"E8A2",
			x"0000" when x"E8A3",
			x"0000" when x"E8A4",
			x"0000" when x"E8A5",
			x"0000" when x"E8A6",
			x"0000" when x"E8A7",
			x"0000" when x"E8A8",
			x"0000" when x"E8A9",
			x"0000" when x"E8AA",
			x"0000" when x"E8AB",
			x"0000" when x"E8AC",
			x"0000" when x"E8AD",
			x"0000" when x"E8AE",
			x"0000" when x"E8AF",
			x"0000" when x"E8B0",
			x"0000" when x"E8B1",
			x"0000" when x"E8B2",
			x"0000" when x"E8B3",
			x"0000" when x"E8B4",
			x"0000" when x"E8B5",
			x"0000" when x"E8B6",
			x"0000" when x"E8B7",
			x"0000" when x"E8B8",
			x"0000" when x"E8B9",
			x"0000" when x"E8BA",
			x"0000" when x"E8BB",
			x"0000" when x"E8BC",
			x"0000" when x"E8BD",
			x"0000" when x"E8BE",
			x"0000" when x"E8BF",
			x"0000" when x"E8C0",
			x"0000" when x"E8C1",
			x"0000" when x"E8C2",
			x"0000" when x"E8C3",
			x"0000" when x"E8C4",
			x"0000" when x"E8C5",
			x"0000" when x"E8C6",
			x"0000" when x"E8C7",
			x"0000" when x"E8C8",
			x"0000" when x"E8C9",
			x"0000" when x"E8CA",
			x"0000" when x"E8CB",
			x"0000" when x"E8CC",
			x"0000" when x"E8CD",
			x"0000" when x"E8CE",
			x"0000" when x"E8CF",
			x"0000" when x"E8D0",
			x"0000" when x"E8D1",
			x"0000" when x"E8D2",
			x"0000" when x"E8D3",
			x"0000" when x"E8D4",
			x"0000" when x"E8D5",
			x"0000" when x"E8D6",
			x"0000" when x"E8D7",
			x"0000" when x"E8D8",
			x"0000" when x"E8D9",
			x"0000" when x"E8DA",
			x"0000" when x"E8DB",
			x"0000" when x"E8DC",
			x"0000" when x"E8DD",
			x"0000" when x"E8DE",
			x"0000" when x"E8DF",
			x"0000" when x"E8E0",
			x"0000" when x"E8E1",
			x"0000" when x"E8E2",
			x"0000" when x"E8E3",
			x"0000" when x"E8E4",
			x"0000" when x"E8E5",
			x"0000" when x"E8E6",
			x"0000" when x"E8E7",
			x"0000" when x"E8E8",
			x"0000" when x"E8E9",
			x"0000" when x"E8EA",
			x"0000" when x"E8EB",
			x"0000" when x"E8EC",
			x"0000" when x"E8ED",
			x"0000" when x"E8EE",
			x"0000" when x"E8EF",
			x"0000" when x"E8F0",
			x"0000" when x"E8F1",
			x"0000" when x"E8F2",
			x"0000" when x"E8F3",
			x"0000" when x"E8F4",
			x"0000" when x"E8F5",
			x"0000" when x"E8F6",
			x"0000" when x"E8F7",
			x"0000" when x"E8F8",
			x"0000" when x"E8F9",
			x"0000" when x"E8FA",
			x"0000" when x"E8FB",
			x"0000" when x"E8FC",
			x"0000" when x"E8FD",
			x"0000" when x"E8FE",
			x"0000" when x"E8FF",
			x"0000" when x"E900",
			x"0000" when x"E901",
			x"0000" when x"E902",
			x"0000" when x"E903",
			x"0000" when x"E904",
			x"0000" when x"E905",
			x"0000" when x"E906",
			x"0000" when x"E907",
			x"0000" when x"E908",
			x"0000" when x"E909",
			x"0000" when x"E90A",
			x"0000" when x"E90B",
			x"0000" when x"E90C",
			x"0000" when x"E90D",
			x"0000" when x"E90E",
			x"0000" when x"E90F",
			x"0000" when x"E910",
			x"0000" when x"E911",
			x"0000" when x"E912",
			x"0000" when x"E913",
			x"0000" when x"E914",
			x"0000" when x"E915",
			x"0000" when x"E916",
			x"0000" when x"E917",
			x"0000" when x"E918",
			x"0000" when x"E919",
			x"0000" when x"E91A",
			x"0000" when x"E91B",
			x"0000" when x"E91C",
			x"0000" when x"E91D",
			x"0000" when x"E91E",
			x"0000" when x"E91F",
			x"0000" when x"E920",
			x"0000" when x"E921",
			x"0000" when x"E922",
			x"0000" when x"E923",
			x"0000" when x"E924",
			x"0000" when x"E925",
			x"0000" when x"E926",
			x"0000" when x"E927",
			x"0000" when x"E928",
			x"0000" when x"E929",
			x"0000" when x"E92A",
			x"0000" when x"E92B",
			x"0000" when x"E92C",
			x"0000" when x"E92D",
			x"0000" when x"E92E",
			x"0000" when x"E92F",
			x"0000" when x"E930",
			x"0000" when x"E931",
			x"0000" when x"E932",
			x"0000" when x"E933",
			x"0000" when x"E934",
			x"0000" when x"E935",
			x"0000" when x"E936",
			x"0000" when x"E937",
			x"0000" when x"E938",
			x"0000" when x"E939",
			x"0000" when x"E93A",
			x"0000" when x"E93B",
			x"0000" when x"E93C",
			x"0000" when x"E93D",
			x"0000" when x"E93E",
			x"0000" when x"E93F",
			x"0000" when x"E940",
			x"0000" when x"E941",
			x"0000" when x"E942",
			x"0000" when x"E943",
			x"0000" when x"E944",
			x"0000" when x"E945",
			x"0000" when x"E946",
			x"0000" when x"E947",
			x"0000" when x"E948",
			x"0000" when x"E949",
			x"0000" when x"E94A",
			x"0000" when x"E94B",
			x"0000" when x"E94C",
			x"0000" when x"E94D",
			x"0000" when x"E94E",
			x"0000" when x"E94F",
			x"0000" when x"E950",
			x"0000" when x"E951",
			x"0000" when x"E952",
			x"0000" when x"E953",
			x"0000" when x"E954",
			x"0000" when x"E955",
			x"0000" when x"E956",
			x"0000" when x"E957",
			x"0000" when x"E958",
			x"0000" when x"E959",
			x"0000" when x"E95A",
			x"0000" when x"E95B",
			x"0000" when x"E95C",
			x"0000" when x"E95D",
			x"0000" when x"E95E",
			x"0000" when x"E95F",
			x"0000" when x"E960",
			x"0000" when x"E961",
			x"0000" when x"E962",
			x"0000" when x"E963",
			x"0000" when x"E964",
			x"0000" when x"E965",
			x"0000" when x"E966",
			x"0000" when x"E967",
			x"0000" when x"E968",
			x"0000" when x"E969",
			x"0000" when x"E96A",
			x"0000" when x"E96B",
			x"0000" when x"E96C",
			x"0000" when x"E96D",
			x"0000" when x"E96E",
			x"0000" when x"E96F",
			x"0000" when x"E970",
			x"0000" when x"E971",
			x"0000" when x"E972",
			x"0000" when x"E973",
			x"0000" when x"E974",
			x"0000" when x"E975",
			x"0000" when x"E976",
			x"0000" when x"E977",
			x"0000" when x"E978",
			x"0000" when x"E979",
			x"0000" when x"E97A",
			x"0000" when x"E97B",
			x"0000" when x"E97C",
			x"0000" when x"E97D",
			x"0000" when x"E97E",
			x"0000" when x"E97F",
			x"0000" when x"E980",
			x"0000" when x"E981",
			x"0000" when x"E982",
			x"0000" when x"E983",
			x"0000" when x"E984",
			x"0000" when x"E985",
			x"0000" when x"E986",
			x"0000" when x"E987",
			x"0000" when x"E988",
			x"0000" when x"E989",
			x"0000" when x"E98A",
			x"0000" when x"E98B",
			x"0000" when x"E98C",
			x"0000" when x"E98D",
			x"0000" when x"E98E",
			x"0000" when x"E98F",
			x"0000" when x"E990",
			x"0000" when x"E991",
			x"0000" when x"E992",
			x"0000" when x"E993",
			x"0000" when x"E994",
			x"0000" when x"E995",
			x"0000" when x"E996",
			x"0000" when x"E997",
			x"0000" when x"E998",
			x"0000" when x"E999",
			x"0000" when x"E99A",
			x"0000" when x"E99B",
			x"0000" when x"E99C",
			x"0000" when x"E99D",
			x"0000" when x"E99E",
			x"0000" when x"E99F",
			x"0000" when x"E9A0",
			x"0000" when x"E9A1",
			x"0000" when x"E9A2",
			x"0000" when x"E9A3",
			x"0000" when x"E9A4",
			x"0000" when x"E9A5",
			x"0000" when x"E9A6",
			x"0000" when x"E9A7",
			x"0000" when x"E9A8",
			x"0000" when x"E9A9",
			x"0000" when x"E9AA",
			x"0000" when x"E9AB",
			x"0000" when x"E9AC",
			x"0000" when x"E9AD",
			x"0000" when x"E9AE",
			x"0000" when x"E9AF",
			x"0000" when x"E9B0",
			x"0000" when x"E9B1",
			x"0000" when x"E9B2",
			x"0000" when x"E9B3",
			x"0000" when x"E9B4",
			x"0000" when x"E9B5",
			x"0000" when x"E9B6",
			x"0000" when x"E9B7",
			x"0000" when x"E9B8",
			x"0000" when x"E9B9",
			x"0000" when x"E9BA",
			x"0000" when x"E9BB",
			x"0000" when x"E9BC",
			x"0000" when x"E9BD",
			x"0000" when x"E9BE",
			x"0000" when x"E9BF",
			x"0000" when x"E9C0",
			x"0000" when x"E9C1",
			x"0000" when x"E9C2",
			x"0000" when x"E9C3",
			x"0000" when x"E9C4",
			x"0000" when x"E9C5",
			x"0000" when x"E9C6",
			x"0000" when x"E9C7",
			x"0000" when x"E9C8",
			x"0000" when x"E9C9",
			x"0000" when x"E9CA",
			x"0000" when x"E9CB",
			x"0000" when x"E9CC",
			x"0000" when x"E9CD",
			x"0000" when x"E9CE",
			x"0000" when x"E9CF",
			x"0000" when x"E9D0",
			x"0000" when x"E9D1",
			x"0000" when x"E9D2",
			x"0000" when x"E9D3",
			x"0000" when x"E9D4",
			x"0000" when x"E9D5",
			x"0000" when x"E9D6",
			x"0000" when x"E9D7",
			x"0000" when x"E9D8",
			x"0000" when x"E9D9",
			x"0000" when x"E9DA",
			x"0000" when x"E9DB",
			x"0000" when x"E9DC",
			x"0000" when x"E9DD",
			x"0000" when x"E9DE",
			x"0000" when x"E9DF",
			x"0000" when x"E9E0",
			x"0000" when x"E9E1",
			x"0000" when x"E9E2",
			x"0000" when x"E9E3",
			x"0000" when x"E9E4",
			x"0000" when x"E9E5",
			x"0000" when x"E9E6",
			x"0000" when x"E9E7",
			x"0000" when x"E9E8",
			x"0000" when x"E9E9",
			x"0000" when x"E9EA",
			x"0000" when x"E9EB",
			x"0000" when x"E9EC",
			x"0000" when x"E9ED",
			x"0000" when x"E9EE",
			x"0000" when x"E9EF",
			x"0000" when x"E9F0",
			x"0000" when x"E9F1",
			x"0000" when x"E9F2",
			x"0000" when x"E9F3",
			x"0000" when x"E9F4",
			x"0000" when x"E9F5",
			x"0000" when x"E9F6",
			x"0000" when x"E9F7",
			x"0000" when x"E9F8",
			x"0000" when x"E9F9",
			x"0000" when x"E9FA",
			x"0000" when x"E9FB",
			x"0000" when x"E9FC",
			x"0000" when x"E9FD",
			x"0000" when x"E9FE",
			x"0000" when x"E9FF",
			x"0000" when x"EA00",
			x"0000" when x"EA01",
			x"0000" when x"EA02",
			x"0000" when x"EA03",
			x"0000" when x"EA04",
			x"0000" when x"EA05",
			x"0000" when x"EA06",
			x"0000" when x"EA07",
			x"0000" when x"EA08",
			x"0000" when x"EA09",
			x"0000" when x"EA0A",
			x"0000" when x"EA0B",
			x"0000" when x"EA0C",
			x"0000" when x"EA0D",
			x"0000" when x"EA0E",
			x"0000" when x"EA0F",
			x"0000" when x"EA10",
			x"0000" when x"EA11",
			x"0000" when x"EA12",
			x"0000" when x"EA13",
			x"0000" when x"EA14",
			x"0000" when x"EA15",
			x"0000" when x"EA16",
			x"0000" when x"EA17",
			x"0000" when x"EA18",
			x"0000" when x"EA19",
			x"0000" when x"EA1A",
			x"0000" when x"EA1B",
			x"0000" when x"EA1C",
			x"0000" when x"EA1D",
			x"0000" when x"EA1E",
			x"0000" when x"EA1F",
			x"0000" when x"EA20",
			x"0000" when x"EA21",
			x"0000" when x"EA22",
			x"0000" when x"EA23",
			x"0000" when x"EA24",
			x"0000" when x"EA25",
			x"0000" when x"EA26",
			x"0000" when x"EA27",
			x"0000" when x"EA28",
			x"0000" when x"EA29",
			x"0000" when x"EA2A",
			x"0000" when x"EA2B",
			x"0000" when x"EA2C",
			x"0000" when x"EA2D",
			x"0000" when x"EA2E",
			x"0000" when x"EA2F",
			x"0000" when x"EA30",
			x"0000" when x"EA31",
			x"0000" when x"EA32",
			x"0000" when x"EA33",
			x"0000" when x"EA34",
			x"0000" when x"EA35",
			x"0000" when x"EA36",
			x"0000" when x"EA37",
			x"0000" when x"EA38",
			x"0000" when x"EA39",
			x"0000" when x"EA3A",
			x"0000" when x"EA3B",
			x"0000" when x"EA3C",
			x"0000" when x"EA3D",
			x"0000" when x"EA3E",
			x"0000" when x"EA3F",
			x"0000" when x"EA40",
			x"0000" when x"EA41",
			x"0000" when x"EA42",
			x"0000" when x"EA43",
			x"0000" when x"EA44",
			x"0000" when x"EA45",
			x"0000" when x"EA46",
			x"0000" when x"EA47",
			x"0000" when x"EA48",
			x"0000" when x"EA49",
			x"0000" when x"EA4A",
			x"0000" when x"EA4B",
			x"0000" when x"EA4C",
			x"0000" when x"EA4D",
			x"0000" when x"EA4E",
			x"0000" when x"EA4F",
			x"0000" when x"EA50",
			x"0000" when x"EA51",
			x"0000" when x"EA52",
			x"0000" when x"EA53",
			x"0000" when x"EA54",
			x"0000" when x"EA55",
			x"0000" when x"EA56",
			x"0000" when x"EA57",
			x"0000" when x"EA58",
			x"0000" when x"EA59",
			x"0000" when x"EA5A",
			x"0000" when x"EA5B",
			x"0000" when x"EA5C",
			x"0000" when x"EA5D",
			x"0000" when x"EA5E",
			x"0000" when x"EA5F",
			x"0000" when x"EA60",
			x"0000" when x"EA61",
			x"0000" when x"EA62",
			x"0000" when x"EA63",
			x"0000" when x"EA64",
			x"0000" when x"EA65",
			x"0000" when x"EA66",
			x"0000" when x"EA67",
			x"0000" when x"EA68",
			x"0000" when x"EA69",
			x"0000" when x"EA6A",
			x"0000" when x"EA6B",
			x"0000" when x"EA6C",
			x"0000" when x"EA6D",
			x"0000" when x"EA6E",
			x"0000" when x"EA6F",
			x"0000" when x"EA70",
			x"0000" when x"EA71",
			x"0000" when x"EA72",
			x"0000" when x"EA73",
			x"0000" when x"EA74",
			x"0000" when x"EA75",
			x"0000" when x"EA76",
			x"0000" when x"EA77",
			x"0000" when x"EA78",
			x"0000" when x"EA79",
			x"0000" when x"EA7A",
			x"0000" when x"EA7B",
			x"0000" when x"EA7C",
			x"0000" when x"EA7D",
			x"0000" when x"EA7E",
			x"0000" when x"EA7F",
			x"0000" when x"EA80",
			x"0000" when x"EA81",
			x"0000" when x"EA82",
			x"0000" when x"EA83",
			x"0000" when x"EA84",
			x"0000" when x"EA85",
			x"0000" when x"EA86",
			x"0000" when x"EA87",
			x"0000" when x"EA88",
			x"0000" when x"EA89",
			x"0000" when x"EA8A",
			x"0000" when x"EA8B",
			x"0000" when x"EA8C",
			x"0000" when x"EA8D",
			x"0000" when x"EA8E",
			x"0000" when x"EA8F",
			x"0000" when x"EA90",
			x"0000" when x"EA91",
			x"0000" when x"EA92",
			x"0000" when x"EA93",
			x"0000" when x"EA94",
			x"0000" when x"EA95",
			x"0000" when x"EA96",
			x"0000" when x"EA97",
			x"0000" when x"EA98",
			x"0000" when x"EA99",
			x"0000" when x"EA9A",
			x"0000" when x"EA9B",
			x"0000" when x"EA9C",
			x"0000" when x"EA9D",
			x"0000" when x"EA9E",
			x"0000" when x"EA9F",
			x"0000" when x"EAA0",
			x"0000" when x"EAA1",
			x"0000" when x"EAA2",
			x"0000" when x"EAA3",
			x"0000" when x"EAA4",
			x"0000" when x"EAA5",
			x"0000" when x"EAA6",
			x"0000" when x"EAA7",
			x"0000" when x"EAA8",
			x"0000" when x"EAA9",
			x"0000" when x"EAAA",
			x"0000" when x"EAAB",
			x"0000" when x"EAAC",
			x"0000" when x"EAAD",
			x"0000" when x"EAAE",
			x"0000" when x"EAAF",
			x"0000" when x"EAB0",
			x"0000" when x"EAB1",
			x"0000" when x"EAB2",
			x"0000" when x"EAB3",
			x"0000" when x"EAB4",
			x"0000" when x"EAB5",
			x"0000" when x"EAB6",
			x"0000" when x"EAB7",
			x"0000" when x"EAB8",
			x"0000" when x"EAB9",
			x"0000" when x"EABA",
			x"0000" when x"EABB",
			x"0000" when x"EABC",
			x"0000" when x"EABD",
			x"0000" when x"EABE",
			x"0000" when x"EABF",
			x"0000" when x"EAC0",
			x"0000" when x"EAC1",
			x"0000" when x"EAC2",
			x"0000" when x"EAC3",
			x"0000" when x"EAC4",
			x"0000" when x"EAC5",
			x"0000" when x"EAC6",
			x"0000" when x"EAC7",
			x"0000" when x"EAC8",
			x"0000" when x"EAC9",
			x"0000" when x"EACA",
			x"0000" when x"EACB",
			x"0000" when x"EACC",
			x"0000" when x"EACD",
			x"0000" when x"EACE",
			x"0000" when x"EACF",
			x"0000" when x"EAD0",
			x"0000" when x"EAD1",
			x"0000" when x"EAD2",
			x"0000" when x"EAD3",
			x"0000" when x"EAD4",
			x"0000" when x"EAD5",
			x"0000" when x"EAD6",
			x"0000" when x"EAD7",
			x"0000" when x"EAD8",
			x"0000" when x"EAD9",
			x"0000" when x"EADA",
			x"0000" when x"EADB",
			x"0000" when x"EADC",
			x"0000" when x"EADD",
			x"0000" when x"EADE",
			x"0000" when x"EADF",
			x"0000" when x"EAE0",
			x"0000" when x"EAE1",
			x"0000" when x"EAE2",
			x"0000" when x"EAE3",
			x"0000" when x"EAE4",
			x"0000" when x"EAE5",
			x"0000" when x"EAE6",
			x"0000" when x"EAE7",
			x"0000" when x"EAE8",
			x"0000" when x"EAE9",
			x"0000" when x"EAEA",
			x"0000" when x"EAEB",
			x"0000" when x"EAEC",
			x"0000" when x"EAED",
			x"0000" when x"EAEE",
			x"0000" when x"EAEF",
			x"0000" when x"EAF0",
			x"0000" when x"EAF1",
			x"0000" when x"EAF2",
			x"0000" when x"EAF3",
			x"0000" when x"EAF4",
			x"0000" when x"EAF5",
			x"0000" when x"EAF6",
			x"0000" when x"EAF7",
			x"0000" when x"EAF8",
			x"0000" when x"EAF9",
			x"0000" when x"EAFA",
			x"0000" when x"EAFB",
			x"0000" when x"EAFC",
			x"0000" when x"EAFD",
			x"0000" when x"EAFE",
			x"0000" when x"EAFF",
			x"0000" when x"EB00",
			x"0000" when x"EB01",
			x"0000" when x"EB02",
			x"0000" when x"EB03",
			x"0000" when x"EB04",
			x"0000" when x"EB05",
			x"0000" when x"EB06",
			x"0000" when x"EB07",
			x"0000" when x"EB08",
			x"0000" when x"EB09",
			x"0000" when x"EB0A",
			x"0000" when x"EB0B",
			x"0000" when x"EB0C",
			x"0000" when x"EB0D",
			x"0000" when x"EB0E",
			x"0000" when x"EB0F",
			x"0000" when x"EB10",
			x"0000" when x"EB11",
			x"0000" when x"EB12",
			x"0000" when x"EB13",
			x"0000" when x"EB14",
			x"0000" when x"EB15",
			x"0000" when x"EB16",
			x"0000" when x"EB17",
			x"0000" when x"EB18",
			x"0000" when x"EB19",
			x"0000" when x"EB1A",
			x"0000" when x"EB1B",
			x"0000" when x"EB1C",
			x"0000" when x"EB1D",
			x"0000" when x"EB1E",
			x"0000" when x"EB1F",
			x"0000" when x"EB20",
			x"0000" when x"EB21",
			x"0000" when x"EB22",
			x"0000" when x"EB23",
			x"0000" when x"EB24",
			x"0000" when x"EB25",
			x"0000" when x"EB26",
			x"0000" when x"EB27",
			x"0000" when x"EB28",
			x"0000" when x"EB29",
			x"0000" when x"EB2A",
			x"0000" when x"EB2B",
			x"0000" when x"EB2C",
			x"0000" when x"EB2D",
			x"0000" when x"EB2E",
			x"0000" when x"EB2F",
			x"0000" when x"EB30",
			x"0000" when x"EB31",
			x"0000" when x"EB32",
			x"0000" when x"EB33",
			x"0000" when x"EB34",
			x"0000" when x"EB35",
			x"0000" when x"EB36",
			x"0000" when x"EB37",
			x"0000" when x"EB38",
			x"0000" when x"EB39",
			x"0000" when x"EB3A",
			x"0000" when x"EB3B",
			x"0000" when x"EB3C",
			x"0000" when x"EB3D",
			x"0000" when x"EB3E",
			x"0000" when x"EB3F",
			x"0000" when x"EB40",
			x"0000" when x"EB41",
			x"0000" when x"EB42",
			x"0000" when x"EB43",
			x"0000" when x"EB44",
			x"0000" when x"EB45",
			x"0000" when x"EB46",
			x"0000" when x"EB47",
			x"0000" when x"EB48",
			x"0000" when x"EB49",
			x"0000" when x"EB4A",
			x"0000" when x"EB4B",
			x"0000" when x"EB4C",
			x"0000" when x"EB4D",
			x"0000" when x"EB4E",
			x"0000" when x"EB4F",
			x"0000" when x"EB50",
			x"0000" when x"EB51",
			x"0000" when x"EB52",
			x"0000" when x"EB53",
			x"0000" when x"EB54",
			x"0000" when x"EB55",
			x"0000" when x"EB56",
			x"0000" when x"EB57",
			x"0000" when x"EB58",
			x"0000" when x"EB59",
			x"0000" when x"EB5A",
			x"0000" when x"EB5B",
			x"0000" when x"EB5C",
			x"0000" when x"EB5D",
			x"0000" when x"EB5E",
			x"0000" when x"EB5F",
			x"0000" when x"EB60",
			x"0000" when x"EB61",
			x"0000" when x"EB62",
			x"0000" when x"EB63",
			x"0000" when x"EB64",
			x"0000" when x"EB65",
			x"0000" when x"EB66",
			x"0000" when x"EB67",
			x"0000" when x"EB68",
			x"0000" when x"EB69",
			x"0000" when x"EB6A",
			x"0000" when x"EB6B",
			x"0000" when x"EB6C",
			x"0000" when x"EB6D",
			x"0000" when x"EB6E",
			x"0000" when x"EB6F",
			x"0000" when x"EB70",
			x"0000" when x"EB71",
			x"0000" when x"EB72",
			x"0000" when x"EB73",
			x"0000" when x"EB74",
			x"0000" when x"EB75",
			x"0000" when x"EB76",
			x"0000" when x"EB77",
			x"0000" when x"EB78",
			x"0000" when x"EB79",
			x"0000" when x"EB7A",
			x"0000" when x"EB7B",
			x"0000" when x"EB7C",
			x"0000" when x"EB7D",
			x"0000" when x"EB7E",
			x"0000" when x"EB7F",
			x"0000" when x"EB80",
			x"0000" when x"EB81",
			x"0000" when x"EB82",
			x"0000" when x"EB83",
			x"0000" when x"EB84",
			x"0000" when x"EB85",
			x"0000" when x"EB86",
			x"0000" when x"EB87",
			x"0000" when x"EB88",
			x"0000" when x"EB89",
			x"0000" when x"EB8A",
			x"0000" when x"EB8B",
			x"0000" when x"EB8C",
			x"0000" when x"EB8D",
			x"0000" when x"EB8E",
			x"0000" when x"EB8F",
			x"0000" when x"EB90",
			x"0000" when x"EB91",
			x"0000" when x"EB92",
			x"0000" when x"EB93",
			x"0000" when x"EB94",
			x"0000" when x"EB95",
			x"0000" when x"EB96",
			x"0000" when x"EB97",
			x"0000" when x"EB98",
			x"0000" when x"EB99",
			x"0000" when x"EB9A",
			x"0000" when x"EB9B",
			x"0000" when x"EB9C",
			x"0000" when x"EB9D",
			x"0000" when x"EB9E",
			x"0000" when x"EB9F",
			x"0000" when x"EBA0",
			x"0000" when x"EBA1",
			x"0000" when x"EBA2",
			x"0000" when x"EBA3",
			x"0000" when x"EBA4",
			x"0000" when x"EBA5",
			x"0000" when x"EBA6",
			x"0000" when x"EBA7",
			x"0000" when x"EBA8",
			x"0000" when x"EBA9",
			x"0000" when x"EBAA",
			x"0000" when x"EBAB",
			x"0000" when x"EBAC",
			x"0000" when x"EBAD",
			x"0000" when x"EBAE",
			x"0000" when x"EBAF",
			x"0000" when x"EBB0",
			x"0000" when x"EBB1",
			x"0000" when x"EBB2",
			x"0000" when x"EBB3",
			x"0000" when x"EBB4",
			x"0000" when x"EBB5",
			x"0000" when x"EBB6",
			x"0000" when x"EBB7",
			x"0000" when x"EBB8",
			x"0000" when x"EBB9",
			x"0000" when x"EBBA",
			x"0000" when x"EBBB",
			x"0000" when x"EBBC",
			x"0000" when x"EBBD",
			x"0000" when x"EBBE",
			x"0000" when x"EBBF",
			x"0000" when x"EBC0",
			x"0000" when x"EBC1",
			x"0000" when x"EBC2",
			x"0000" when x"EBC3",
			x"0000" when x"EBC4",
			x"0000" when x"EBC5",
			x"0000" when x"EBC6",
			x"0000" when x"EBC7",
			x"0000" when x"EBC8",
			x"0000" when x"EBC9",
			x"0000" when x"EBCA",
			x"0000" when x"EBCB",
			x"0000" when x"EBCC",
			x"0000" when x"EBCD",
			x"0000" when x"EBCE",
			x"0000" when x"EBCF",
			x"0000" when x"EBD0",
			x"0000" when x"EBD1",
			x"0000" when x"EBD2",
			x"0000" when x"EBD3",
			x"0000" when x"EBD4",
			x"0000" when x"EBD5",
			x"0000" when x"EBD6",
			x"0000" when x"EBD7",
			x"0000" when x"EBD8",
			x"0000" when x"EBD9",
			x"0000" when x"EBDA",
			x"0000" when x"EBDB",
			x"0000" when x"EBDC",
			x"0000" when x"EBDD",
			x"0000" when x"EBDE",
			x"0000" when x"EBDF",
			x"0000" when x"EBE0",
			x"0000" when x"EBE1",
			x"0000" when x"EBE2",
			x"0000" when x"EBE3",
			x"0000" when x"EBE4",
			x"0000" when x"EBE5",
			x"0000" when x"EBE6",
			x"0000" when x"EBE7",
			x"0000" when x"EBE8",
			x"0000" when x"EBE9",
			x"0000" when x"EBEA",
			x"0000" when x"EBEB",
			x"0000" when x"EBEC",
			x"0000" when x"EBED",
			x"0000" when x"EBEE",
			x"0000" when x"EBEF",
			x"0000" when x"EBF0",
			x"0000" when x"EBF1",
			x"0000" when x"EBF2",
			x"0000" when x"EBF3",
			x"0000" when x"EBF4",
			x"0000" when x"EBF5",
			x"0000" when x"EBF6",
			x"0000" when x"EBF7",
			x"0000" when x"EBF8",
			x"0000" when x"EBF9",
			x"0000" when x"EBFA",
			x"0000" when x"EBFB",
			x"0000" when x"EBFC",
			x"0000" when x"EBFD",
			x"0000" when x"EBFE",
			x"0000" when x"EBFF",
			x"0000" when x"EC00",
			x"0000" when x"EC01",
			x"0000" when x"EC02",
			x"0000" when x"EC03",
			x"0000" when x"EC04",
			x"0000" when x"EC05",
			x"0000" when x"EC06",
			x"0000" when x"EC07",
			x"0000" when x"EC08",
			x"0000" when x"EC09",
			x"0000" when x"EC0A",
			x"0000" when x"EC0B",
			x"0000" when x"EC0C",
			x"0000" when x"EC0D",
			x"0000" when x"EC0E",
			x"0000" when x"EC0F",
			x"0000" when x"EC10",
			x"0000" when x"EC11",
			x"0000" when x"EC12",
			x"0000" when x"EC13",
			x"0000" when x"EC14",
			x"0000" when x"EC15",
			x"0000" when x"EC16",
			x"0000" when x"EC17",
			x"0000" when x"EC18",
			x"0000" when x"EC19",
			x"0000" when x"EC1A",
			x"0000" when x"EC1B",
			x"0000" when x"EC1C",
			x"0000" when x"EC1D",
			x"0000" when x"EC1E",
			x"0000" when x"EC1F",
			x"0000" when x"EC20",
			x"0000" when x"EC21",
			x"0000" when x"EC22",
			x"0000" when x"EC23",
			x"0000" when x"EC24",
			x"0000" when x"EC25",
			x"0000" when x"EC26",
			x"0000" when x"EC27",
			x"0000" when x"EC28",
			x"0000" when x"EC29",
			x"0000" when x"EC2A",
			x"0000" when x"EC2B",
			x"0000" when x"EC2C",
			x"0000" when x"EC2D",
			x"0000" when x"EC2E",
			x"0000" when x"EC2F",
			x"0000" when x"EC30",
			x"0000" when x"EC31",
			x"0000" when x"EC32",
			x"0000" when x"EC33",
			x"0000" when x"EC34",
			x"0000" when x"EC35",
			x"0000" when x"EC36",
			x"0000" when x"EC37",
			x"0000" when x"EC38",
			x"0000" when x"EC39",
			x"0000" when x"EC3A",
			x"0000" when x"EC3B",
			x"0000" when x"EC3C",
			x"0000" when x"EC3D",
			x"0000" when x"EC3E",
			x"0000" when x"EC3F",
			x"0000" when x"EC40",
			x"0000" when x"EC41",
			x"0000" when x"EC42",
			x"0000" when x"EC43",
			x"0000" when x"EC44",
			x"0000" when x"EC45",
			x"0000" when x"EC46",
			x"0000" when x"EC47",
			x"0000" when x"EC48",
			x"0000" when x"EC49",
			x"0000" when x"EC4A",
			x"0000" when x"EC4B",
			x"0000" when x"EC4C",
			x"0000" when x"EC4D",
			x"0000" when x"EC4E",
			x"0000" when x"EC4F",
			x"0000" when x"EC50",
			x"0000" when x"EC51",
			x"0000" when x"EC52",
			x"0000" when x"EC53",
			x"0000" when x"EC54",
			x"0000" when x"EC55",
			x"0000" when x"EC56",
			x"0000" when x"EC57",
			x"0000" when x"EC58",
			x"0000" when x"EC59",
			x"0000" when x"EC5A",
			x"0000" when x"EC5B",
			x"0000" when x"EC5C",
			x"0000" when x"EC5D",
			x"0000" when x"EC5E",
			x"0000" when x"EC5F",
			x"0000" when x"EC60",
			x"0000" when x"EC61",
			x"0000" when x"EC62",
			x"0000" when x"EC63",
			x"0000" when x"EC64",
			x"0000" when x"EC65",
			x"0000" when x"EC66",
			x"0000" when x"EC67",
			x"0000" when x"EC68",
			x"0000" when x"EC69",
			x"0000" when x"EC6A",
			x"0000" when x"EC6B",
			x"0000" when x"EC6C",
			x"0000" when x"EC6D",
			x"0000" when x"EC6E",
			x"0000" when x"EC6F",
			x"0000" when x"EC70",
			x"0000" when x"EC71",
			x"0000" when x"EC72",
			x"0000" when x"EC73",
			x"0000" when x"EC74",
			x"0000" when x"EC75",
			x"0000" when x"EC76",
			x"0000" when x"EC77",
			x"0000" when x"EC78",
			x"0000" when x"EC79",
			x"0000" when x"EC7A",
			x"0000" when x"EC7B",
			x"0000" when x"EC7C",
			x"0000" when x"EC7D",
			x"0000" when x"EC7E",
			x"0000" when x"EC7F",
			x"0000" when x"EC80",
			x"0000" when x"EC81",
			x"0000" when x"EC82",
			x"0000" when x"EC83",
			x"0000" when x"EC84",
			x"0000" when x"EC85",
			x"0000" when x"EC86",
			x"0000" when x"EC87",
			x"0000" when x"EC88",
			x"0000" when x"EC89",
			x"0000" when x"EC8A",
			x"0000" when x"EC8B",
			x"0000" when x"EC8C",
			x"0000" when x"EC8D",
			x"0000" when x"EC8E",
			x"0000" when x"EC8F",
			x"0000" when x"EC90",
			x"0000" when x"EC91",
			x"0000" when x"EC92",
			x"0000" when x"EC93",
			x"0000" when x"EC94",
			x"0000" when x"EC95",
			x"0000" when x"EC96",
			x"0000" when x"EC97",
			x"0000" when x"EC98",
			x"0000" when x"EC99",
			x"0000" when x"EC9A",
			x"0000" when x"EC9B",
			x"0000" when x"EC9C",
			x"0000" when x"EC9D",
			x"0000" when x"EC9E",
			x"0000" when x"EC9F",
			x"0000" when x"ECA0",
			x"0000" when x"ECA1",
			x"0000" when x"ECA2",
			x"0000" when x"ECA3",
			x"0000" when x"ECA4",
			x"0000" when x"ECA5",
			x"0000" when x"ECA6",
			x"0000" when x"ECA7",
			x"0000" when x"ECA8",
			x"0000" when x"ECA9",
			x"0000" when x"ECAA",
			x"0000" when x"ECAB",
			x"0000" when x"ECAC",
			x"0000" when x"ECAD",
			x"0000" when x"ECAE",
			x"0000" when x"ECAF",
			x"0000" when x"ECB0",
			x"0000" when x"ECB1",
			x"0000" when x"ECB2",
			x"0000" when x"ECB3",
			x"0000" when x"ECB4",
			x"0000" when x"ECB5",
			x"0000" when x"ECB6",
			x"0000" when x"ECB7",
			x"0000" when x"ECB8",
			x"0000" when x"ECB9",
			x"0000" when x"ECBA",
			x"0000" when x"ECBB",
			x"0000" when x"ECBC",
			x"0000" when x"ECBD",
			x"0000" when x"ECBE",
			x"0000" when x"ECBF",
			x"0000" when x"ECC0",
			x"0000" when x"ECC1",
			x"0000" when x"ECC2",
			x"0000" when x"ECC3",
			x"0000" when x"ECC4",
			x"0000" when x"ECC5",
			x"0000" when x"ECC6",
			x"0000" when x"ECC7",
			x"0000" when x"ECC8",
			x"0000" when x"ECC9",
			x"0000" when x"ECCA",
			x"0000" when x"ECCB",
			x"0000" when x"ECCC",
			x"0000" when x"ECCD",
			x"0000" when x"ECCE",
			x"0000" when x"ECCF",
			x"0000" when x"ECD0",
			x"0000" when x"ECD1",
			x"0000" when x"ECD2",
			x"0000" when x"ECD3",
			x"0000" when x"ECD4",
			x"0000" when x"ECD5",
			x"0000" when x"ECD6",
			x"0000" when x"ECD7",
			x"0000" when x"ECD8",
			x"0000" when x"ECD9",
			x"0000" when x"ECDA",
			x"0000" when x"ECDB",
			x"0000" when x"ECDC",
			x"0000" when x"ECDD",
			x"0000" when x"ECDE",
			x"0000" when x"ECDF",
			x"0000" when x"ECE0",
			x"0000" when x"ECE1",
			x"0000" when x"ECE2",
			x"0000" when x"ECE3",
			x"0000" when x"ECE4",
			x"0000" when x"ECE5",
			x"0000" when x"ECE6",
			x"0000" when x"ECE7",
			x"0000" when x"ECE8",
			x"0000" when x"ECE9",
			x"0000" when x"ECEA",
			x"0000" when x"ECEB",
			x"0000" when x"ECEC",
			x"0000" when x"ECED",
			x"0000" when x"ECEE",
			x"0000" when x"ECEF",
			x"0000" when x"ECF0",
			x"0000" when x"ECF1",
			x"0000" when x"ECF2",
			x"0000" when x"ECF3",
			x"0000" when x"ECF4",
			x"0000" when x"ECF5",
			x"0000" when x"ECF6",
			x"0000" when x"ECF7",
			x"0000" when x"ECF8",
			x"0000" when x"ECF9",
			x"0000" when x"ECFA",
			x"0000" when x"ECFB",
			x"0000" when x"ECFC",
			x"0000" when x"ECFD",
			x"0000" when x"ECFE",
			x"0000" when x"ECFF",
			x"0000" when x"ED00",
			x"0000" when x"ED01",
			x"0000" when x"ED02",
			x"0000" when x"ED03",
			x"0000" when x"ED04",
			x"0000" when x"ED05",
			x"0000" when x"ED06",
			x"0000" when x"ED07",
			x"0000" when x"ED08",
			x"0000" when x"ED09",
			x"0000" when x"ED0A",
			x"0000" when x"ED0B",
			x"0000" when x"ED0C",
			x"0000" when x"ED0D",
			x"0000" when x"ED0E",
			x"0000" when x"ED0F",
			x"0000" when x"ED10",
			x"0000" when x"ED11",
			x"0000" when x"ED12",
			x"0000" when x"ED13",
			x"0000" when x"ED14",
			x"0000" when x"ED15",
			x"0000" when x"ED16",
			x"0000" when x"ED17",
			x"0000" when x"ED18",
			x"0000" when x"ED19",
			x"0000" when x"ED1A",
			x"0000" when x"ED1B",
			x"0000" when x"ED1C",
			x"0000" when x"ED1D",
			x"0000" when x"ED1E",
			x"0000" when x"ED1F",
			x"0000" when x"ED20",
			x"0000" when x"ED21",
			x"0000" when x"ED22",
			x"0000" when x"ED23",
			x"0000" when x"ED24",
			x"0000" when x"ED25",
			x"0000" when x"ED26",
			x"0000" when x"ED27",
			x"0000" when x"ED28",
			x"0000" when x"ED29",
			x"0000" when x"ED2A",
			x"0000" when x"ED2B",
			x"0000" when x"ED2C",
			x"0000" when x"ED2D",
			x"0000" when x"ED2E",
			x"0000" when x"ED2F",
			x"0000" when x"ED30",
			x"0000" when x"ED31",
			x"0000" when x"ED32",
			x"0000" when x"ED33",
			x"0000" when x"ED34",
			x"0000" when x"ED35",
			x"0000" when x"ED36",
			x"0000" when x"ED37",
			x"0000" when x"ED38",
			x"0000" when x"ED39",
			x"0000" when x"ED3A",
			x"0000" when x"ED3B",
			x"0000" when x"ED3C",
			x"0000" when x"ED3D",
			x"0000" when x"ED3E",
			x"0000" when x"ED3F",
			x"0000" when x"ED40",
			x"0000" when x"ED41",
			x"0000" when x"ED42",
			x"0000" when x"ED43",
			x"0000" when x"ED44",
			x"0000" when x"ED45",
			x"0000" when x"ED46",
			x"0000" when x"ED47",
			x"0000" when x"ED48",
			x"0000" when x"ED49",
			x"0000" when x"ED4A",
			x"0000" when x"ED4B",
			x"0000" when x"ED4C",
			x"0000" when x"ED4D",
			x"0000" when x"ED4E",
			x"0000" when x"ED4F",
			x"0000" when x"ED50",
			x"0000" when x"ED51",
			x"0000" when x"ED52",
			x"0000" when x"ED53",
			x"0000" when x"ED54",
			x"0000" when x"ED55",
			x"0000" when x"ED56",
			x"0000" when x"ED57",
			x"0000" when x"ED58",
			x"0000" when x"ED59",
			x"0000" when x"ED5A",
			x"0000" when x"ED5B",
			x"0000" when x"ED5C",
			x"0000" when x"ED5D",
			x"0000" when x"ED5E",
			x"0000" when x"ED5F",
			x"0000" when x"ED60",
			x"0000" when x"ED61",
			x"0000" when x"ED62",
			x"0000" when x"ED63",
			x"0000" when x"ED64",
			x"0000" when x"ED65",
			x"0000" when x"ED66",
			x"0000" when x"ED67",
			x"0000" when x"ED68",
			x"0000" when x"ED69",
			x"0000" when x"ED6A",
			x"0000" when x"ED6B",
			x"0000" when x"ED6C",
			x"0000" when x"ED6D",
			x"0000" when x"ED6E",
			x"0000" when x"ED6F",
			x"0000" when x"ED70",
			x"0000" when x"ED71",
			x"0000" when x"ED72",
			x"0000" when x"ED73",
			x"0000" when x"ED74",
			x"0000" when x"ED75",
			x"0000" when x"ED76",
			x"0000" when x"ED77",
			x"0000" when x"ED78",
			x"0000" when x"ED79",
			x"0000" when x"ED7A",
			x"0000" when x"ED7B",
			x"0000" when x"ED7C",
			x"0000" when x"ED7D",
			x"0000" when x"ED7E",
			x"0000" when x"ED7F",
			x"0000" when x"ED80",
			x"0000" when x"ED81",
			x"0000" when x"ED82",
			x"0000" when x"ED83",
			x"0000" when x"ED84",
			x"0000" when x"ED85",
			x"0000" when x"ED86",
			x"0000" when x"ED87",
			x"0000" when x"ED88",
			x"0000" when x"ED89",
			x"0000" when x"ED8A",
			x"0000" when x"ED8B",
			x"0000" when x"ED8C",
			x"0000" when x"ED8D",
			x"0000" when x"ED8E",
			x"0000" when x"ED8F",
			x"0000" when x"ED90",
			x"0000" when x"ED91",
			x"0000" when x"ED92",
			x"0000" when x"ED93",
			x"0000" when x"ED94",
			x"0000" when x"ED95",
			x"0000" when x"ED96",
			x"0000" when x"ED97",
			x"0000" when x"ED98",
			x"0000" when x"ED99",
			x"0000" when x"ED9A",
			x"0000" when x"ED9B",
			x"0000" when x"ED9C",
			x"0000" when x"ED9D",
			x"0000" when x"ED9E",
			x"0000" when x"ED9F",
			x"0000" when x"EDA0",
			x"0000" when x"EDA1",
			x"0000" when x"EDA2",
			x"0000" when x"EDA3",
			x"0000" when x"EDA4",
			x"0000" when x"EDA5",
			x"0000" when x"EDA6",
			x"0000" when x"EDA7",
			x"0000" when x"EDA8",
			x"0000" when x"EDA9",
			x"0000" when x"EDAA",
			x"0000" when x"EDAB",
			x"0000" when x"EDAC",
			x"0000" when x"EDAD",
			x"0000" when x"EDAE",
			x"0000" when x"EDAF",
			x"0000" when x"EDB0",
			x"0000" when x"EDB1",
			x"0000" when x"EDB2",
			x"0000" when x"EDB3",
			x"0000" when x"EDB4",
			x"0000" when x"EDB5",
			x"0000" when x"EDB6",
			x"0000" when x"EDB7",
			x"0000" when x"EDB8",
			x"0000" when x"EDB9",
			x"0000" when x"EDBA",
			x"0000" when x"EDBB",
			x"0000" when x"EDBC",
			x"0000" when x"EDBD",
			x"0000" when x"EDBE",
			x"0000" when x"EDBF",
			x"0000" when x"EDC0",
			x"0000" when x"EDC1",
			x"0000" when x"EDC2",
			x"0000" when x"EDC3",
			x"0000" when x"EDC4",
			x"0000" when x"EDC5",
			x"0000" when x"EDC6",
			x"0000" when x"EDC7",
			x"0000" when x"EDC8",
			x"0000" when x"EDC9",
			x"0000" when x"EDCA",
			x"0000" when x"EDCB",
			x"0000" when x"EDCC",
			x"0000" when x"EDCD",
			x"0000" when x"EDCE",
			x"0000" when x"EDCF",
			x"0000" when x"EDD0",
			x"0000" when x"EDD1",
			x"0000" when x"EDD2",
			x"0000" when x"EDD3",
			x"0000" when x"EDD4",
			x"0000" when x"EDD5",
			x"0000" when x"EDD6",
			x"0000" when x"EDD7",
			x"0000" when x"EDD8",
			x"0000" when x"EDD9",
			x"0000" when x"EDDA",
			x"0000" when x"EDDB",
			x"0000" when x"EDDC",
			x"0000" when x"EDDD",
			x"0000" when x"EDDE",
			x"0000" when x"EDDF",
			x"0000" when x"EDE0",
			x"0000" when x"EDE1",
			x"0000" when x"EDE2",
			x"0000" when x"EDE3",
			x"0000" when x"EDE4",
			x"0000" when x"EDE5",
			x"0000" when x"EDE6",
			x"0000" when x"EDE7",
			x"0000" when x"EDE8",
			x"0000" when x"EDE9",
			x"0000" when x"EDEA",
			x"0000" when x"EDEB",
			x"0000" when x"EDEC",
			x"0000" when x"EDED",
			x"0000" when x"EDEE",
			x"0000" when x"EDEF",
			x"0000" when x"EDF0",
			x"0000" when x"EDF1",
			x"0000" when x"EDF2",
			x"0000" when x"EDF3",
			x"0000" when x"EDF4",
			x"0000" when x"EDF5",
			x"0000" when x"EDF6",
			x"0000" when x"EDF7",
			x"0000" when x"EDF8",
			x"0000" when x"EDF9",
			x"0000" when x"EDFA",
			x"0000" when x"EDFB",
			x"0000" when x"EDFC",
			x"0000" when x"EDFD",
			x"0000" when x"EDFE",
			x"0000" when x"EDFF",
			x"0000" when x"EE00",
			x"0000" when x"EE01",
			x"0000" when x"EE02",
			x"0000" when x"EE03",
			x"0000" when x"EE04",
			x"0000" when x"EE05",
			x"0000" when x"EE06",
			x"0000" when x"EE07",
			x"0000" when x"EE08",
			x"0000" when x"EE09",
			x"0000" when x"EE0A",
			x"0000" when x"EE0B",
			x"0000" when x"EE0C",
			x"0000" when x"EE0D",
			x"0000" when x"EE0E",
			x"0000" when x"EE0F",
			x"0000" when x"EE10",
			x"0000" when x"EE11",
			x"0000" when x"EE12",
			x"0000" when x"EE13",
			x"0000" when x"EE14",
			x"0000" when x"EE15",
			x"0000" when x"EE16",
			x"0000" when x"EE17",
			x"0000" when x"EE18",
			x"0000" when x"EE19",
			x"0000" when x"EE1A",
			x"0000" when x"EE1B",
			x"0000" when x"EE1C",
			x"0000" when x"EE1D",
			x"0000" when x"EE1E",
			x"0000" when x"EE1F",
			x"0000" when x"EE20",
			x"0000" when x"EE21",
			x"0000" when x"EE22",
			x"0000" when x"EE23",
			x"0000" when x"EE24",
			x"0000" when x"EE25",
			x"0000" when x"EE26",
			x"0000" when x"EE27",
			x"0000" when x"EE28",
			x"0000" when x"EE29",
			x"0000" when x"EE2A",
			x"0000" when x"EE2B",
			x"0000" when x"EE2C",
			x"0000" when x"EE2D",
			x"0000" when x"EE2E",
			x"0000" when x"EE2F",
			x"0000" when x"EE30",
			x"0000" when x"EE31",
			x"0000" when x"EE32",
			x"0000" when x"EE33",
			x"0000" when x"EE34",
			x"0000" when x"EE35",
			x"0000" when x"EE36",
			x"0000" when x"EE37",
			x"0000" when x"EE38",
			x"0000" when x"EE39",
			x"0000" when x"EE3A",
			x"0000" when x"EE3B",
			x"0000" when x"EE3C",
			x"0000" when x"EE3D",
			x"0000" when x"EE3E",
			x"0000" when x"EE3F",
			x"0000" when x"EE40",
			x"0000" when x"EE41",
			x"0000" when x"EE42",
			x"0000" when x"EE43",
			x"0000" when x"EE44",
			x"0000" when x"EE45",
			x"0000" when x"EE46",
			x"0000" when x"EE47",
			x"0000" when x"EE48",
			x"0000" when x"EE49",
			x"0000" when x"EE4A",
			x"0000" when x"EE4B",
			x"0000" when x"EE4C",
			x"0000" when x"EE4D",
			x"0000" when x"EE4E",
			x"0000" when x"EE4F",
			x"0000" when x"EE50",
			x"0000" when x"EE51",
			x"0000" when x"EE52",
			x"0000" when x"EE53",
			x"0000" when x"EE54",
			x"0000" when x"EE55",
			x"0000" when x"EE56",
			x"0000" when x"EE57",
			x"0000" when x"EE58",
			x"0000" when x"EE59",
			x"0000" when x"EE5A",
			x"0000" when x"EE5B",
			x"0000" when x"EE5C",
			x"0000" when x"EE5D",
			x"0000" when x"EE5E",
			x"0000" when x"EE5F",
			x"0000" when x"EE60",
			x"0000" when x"EE61",
			x"0000" when x"EE62",
			x"0000" when x"EE63",
			x"0000" when x"EE64",
			x"0000" when x"EE65",
			x"0000" when x"EE66",
			x"0000" when x"EE67",
			x"0000" when x"EE68",
			x"0000" when x"EE69",
			x"0000" when x"EE6A",
			x"0000" when x"EE6B",
			x"0000" when x"EE6C",
			x"0000" when x"EE6D",
			x"0000" when x"EE6E",
			x"0000" when x"EE6F",
			x"0000" when x"EE70",
			x"0000" when x"EE71",
			x"0000" when x"EE72",
			x"0000" when x"EE73",
			x"0000" when x"EE74",
			x"0000" when x"EE75",
			x"0000" when x"EE76",
			x"0000" when x"EE77",
			x"0000" when x"EE78",
			x"0000" when x"EE79",
			x"0000" when x"EE7A",
			x"0000" when x"EE7B",
			x"0000" when x"EE7C",
			x"0000" when x"EE7D",
			x"0000" when x"EE7E",
			x"0000" when x"EE7F",
			x"0000" when x"EE80",
			x"0000" when x"EE81",
			x"0000" when x"EE82",
			x"0000" when x"EE83",
			x"0000" when x"EE84",
			x"0000" when x"EE85",
			x"0000" when x"EE86",
			x"0000" when x"EE87",
			x"0000" when x"EE88",
			x"0000" when x"EE89",
			x"0000" when x"EE8A",
			x"0000" when x"EE8B",
			x"0000" when x"EE8C",
			x"0000" when x"EE8D",
			x"0000" when x"EE8E",
			x"0000" when x"EE8F",
			x"0000" when x"EE90",
			x"0000" when x"EE91",
			x"0000" when x"EE92",
			x"0000" when x"EE93",
			x"0000" when x"EE94",
			x"0000" when x"EE95",
			x"0000" when x"EE96",
			x"0000" when x"EE97",
			x"0000" when x"EE98",
			x"0000" when x"EE99",
			x"0000" when x"EE9A",
			x"0000" when x"EE9B",
			x"0000" when x"EE9C",
			x"0000" when x"EE9D",
			x"0000" when x"EE9E",
			x"0000" when x"EE9F",
			x"0000" when x"EEA0",
			x"0000" when x"EEA1",
			x"0000" when x"EEA2",
			x"0000" when x"EEA3",
			x"0000" when x"EEA4",
			x"0000" when x"EEA5",
			x"0000" when x"EEA6",
			x"0000" when x"EEA7",
			x"0000" when x"EEA8",
			x"0000" when x"EEA9",
			x"0000" when x"EEAA",
			x"0000" when x"EEAB",
			x"0000" when x"EEAC",
			x"0000" when x"EEAD",
			x"0000" when x"EEAE",
			x"0000" when x"EEAF",
			x"0000" when x"EEB0",
			x"0000" when x"EEB1",
			x"0000" when x"EEB2",
			x"0000" when x"EEB3",
			x"0000" when x"EEB4",
			x"0000" when x"EEB5",
			x"0000" when x"EEB6",
			x"0000" when x"EEB7",
			x"0000" when x"EEB8",
			x"0000" when x"EEB9",
			x"0000" when x"EEBA",
			x"0000" when x"EEBB",
			x"0000" when x"EEBC",
			x"0000" when x"EEBD",
			x"0000" when x"EEBE",
			x"0000" when x"EEBF",
			x"0000" when x"EEC0",
			x"0000" when x"EEC1",
			x"0000" when x"EEC2",
			x"0000" when x"EEC3",
			x"0000" when x"EEC4",
			x"0000" when x"EEC5",
			x"0000" when x"EEC6",
			x"0000" when x"EEC7",
			x"0000" when x"EEC8",
			x"0000" when x"EEC9",
			x"0000" when x"EECA",
			x"0000" when x"EECB",
			x"0000" when x"EECC",
			x"0000" when x"EECD",
			x"0000" when x"EECE",
			x"0000" when x"EECF",
			x"0000" when x"EED0",
			x"0000" when x"EED1",
			x"0000" when x"EED2",
			x"0000" when x"EED3",
			x"0000" when x"EED4",
			x"0000" when x"EED5",
			x"0000" when x"EED6",
			x"0000" when x"EED7",
			x"0000" when x"EED8",
			x"0000" when x"EED9",
			x"0000" when x"EEDA",
			x"0000" when x"EEDB",
			x"0000" when x"EEDC",
			x"0000" when x"EEDD",
			x"0000" when x"EEDE",
			x"0000" when x"EEDF",
			x"0000" when x"EEE0",
			x"0000" when x"EEE1",
			x"0000" when x"EEE2",
			x"0000" when x"EEE3",
			x"0000" when x"EEE4",
			x"0000" when x"EEE5",
			x"0000" when x"EEE6",
			x"0000" when x"EEE7",
			x"0000" when x"EEE8",
			x"0000" when x"EEE9",
			x"0000" when x"EEEA",
			x"0000" when x"EEEB",
			x"0000" when x"EEEC",
			x"0000" when x"EEED",
			x"0000" when x"EEEE",
			x"0000" when x"EEEF",
			x"0000" when x"EEF0",
			x"0000" when x"EEF1",
			x"0000" when x"EEF2",
			x"0000" when x"EEF3",
			x"0000" when x"EEF4",
			x"0000" when x"EEF5",
			x"0000" when x"EEF6",
			x"0000" when x"EEF7",
			x"0000" when x"EEF8",
			x"0000" when x"EEF9",
			x"0000" when x"EEFA",
			x"0000" when x"EEFB",
			x"0000" when x"EEFC",
			x"0000" when x"EEFD",
			x"0000" when x"EEFE",
			x"0000" when x"EEFF",
			x"0000" when x"EF00",
			x"0000" when x"EF01",
			x"0000" when x"EF02",
			x"0000" when x"EF03",
			x"0000" when x"EF04",
			x"0000" when x"EF05",
			x"0000" when x"EF06",
			x"0000" when x"EF07",
			x"0000" when x"EF08",
			x"0000" when x"EF09",
			x"0000" when x"EF0A",
			x"0000" when x"EF0B",
			x"0000" when x"EF0C",
			x"0000" when x"EF0D",
			x"0000" when x"EF0E",
			x"0000" when x"EF0F",
			x"0000" when x"EF10",
			x"0000" when x"EF11",
			x"0000" when x"EF12",
			x"0000" when x"EF13",
			x"0000" when x"EF14",
			x"0000" when x"EF15",
			x"0000" when x"EF16",
			x"0000" when x"EF17",
			x"0000" when x"EF18",
			x"0000" when x"EF19",
			x"0000" when x"EF1A",
			x"0000" when x"EF1B",
			x"0000" when x"EF1C",
			x"0000" when x"EF1D",
			x"0000" when x"EF1E",
			x"0000" when x"EF1F",
			x"0000" when x"EF20",
			x"0000" when x"EF21",
			x"0000" when x"EF22",
			x"0000" when x"EF23",
			x"0000" when x"EF24",
			x"0000" when x"EF25",
			x"0000" when x"EF26",
			x"0000" when x"EF27",
			x"0000" when x"EF28",
			x"0000" when x"EF29",
			x"0000" when x"EF2A",
			x"0000" when x"EF2B",
			x"0000" when x"EF2C",
			x"0000" when x"EF2D",
			x"0000" when x"EF2E",
			x"0000" when x"EF2F",
			x"0000" when x"EF30",
			x"0000" when x"EF31",
			x"0000" when x"EF32",
			x"0000" when x"EF33",
			x"0000" when x"EF34",
			x"0000" when x"EF35",
			x"0000" when x"EF36",
			x"0000" when x"EF37",
			x"0000" when x"EF38",
			x"0000" when x"EF39",
			x"0000" when x"EF3A",
			x"0000" when x"EF3B",
			x"0000" when x"EF3C",
			x"0000" when x"EF3D",
			x"0000" when x"EF3E",
			x"0000" when x"EF3F",
			x"0000" when x"EF40",
			x"0000" when x"EF41",
			x"0000" when x"EF42",
			x"0000" when x"EF43",
			x"0000" when x"EF44",
			x"0000" when x"EF45",
			x"0000" when x"EF46",
			x"0000" when x"EF47",
			x"0000" when x"EF48",
			x"0000" when x"EF49",
			x"0000" when x"EF4A",
			x"0000" when x"EF4B",
			x"0000" when x"EF4C",
			x"0000" when x"EF4D",
			x"0000" when x"EF4E",
			x"0000" when x"EF4F",
			x"0000" when x"EF50",
			x"0000" when x"EF51",
			x"0000" when x"EF52",
			x"0000" when x"EF53",
			x"0000" when x"EF54",
			x"0000" when x"EF55",
			x"0000" when x"EF56",
			x"0000" when x"EF57",
			x"0000" when x"EF58",
			x"0000" when x"EF59",
			x"0000" when x"EF5A",
			x"0000" when x"EF5B",
			x"0000" when x"EF5C",
			x"0000" when x"EF5D",
			x"0000" when x"EF5E",
			x"0000" when x"EF5F",
			x"0000" when x"EF60",
			x"0000" when x"EF61",
			x"0000" when x"EF62",
			x"0000" when x"EF63",
			x"0000" when x"EF64",
			x"0000" when x"EF65",
			x"0000" when x"EF66",
			x"0000" when x"EF67",
			x"0000" when x"EF68",
			x"0000" when x"EF69",
			x"0000" when x"EF6A",
			x"0000" when x"EF6B",
			x"0000" when x"EF6C",
			x"0000" when x"EF6D",
			x"0000" when x"EF6E",
			x"0000" when x"EF6F",
			x"0000" when x"EF70",
			x"0000" when x"EF71",
			x"0000" when x"EF72",
			x"0000" when x"EF73",
			x"0000" when x"EF74",
			x"0000" when x"EF75",
			x"0000" when x"EF76",
			x"0000" when x"EF77",
			x"0000" when x"EF78",
			x"0000" when x"EF79",
			x"0000" when x"EF7A",
			x"0000" when x"EF7B",
			x"0000" when x"EF7C",
			x"0000" when x"EF7D",
			x"0000" when x"EF7E",
			x"0000" when x"EF7F",
			x"0000" when x"EF80",
			x"0000" when x"EF81",
			x"0000" when x"EF82",
			x"0000" when x"EF83",
			x"0000" when x"EF84",
			x"0000" when x"EF85",
			x"0000" when x"EF86",
			x"0000" when x"EF87",
			x"0000" when x"EF88",
			x"0000" when x"EF89",
			x"0000" when x"EF8A",
			x"0000" when x"EF8B",
			x"0000" when x"EF8C",
			x"0000" when x"EF8D",
			x"0000" when x"EF8E",
			x"0000" when x"EF8F",
			x"0000" when x"EF90",
			x"0000" when x"EF91",
			x"0000" when x"EF92",
			x"0000" when x"EF93",
			x"0000" when x"EF94",
			x"0000" when x"EF95",
			x"0000" when x"EF96",
			x"0000" when x"EF97",
			x"0000" when x"EF98",
			x"0000" when x"EF99",
			x"0000" when x"EF9A",
			x"0000" when x"EF9B",
			x"0000" when x"EF9C",
			x"0000" when x"EF9D",
			x"0000" when x"EF9E",
			x"0000" when x"EF9F",
			x"0000" when x"EFA0",
			x"0000" when x"EFA1",
			x"0000" when x"EFA2",
			x"0000" when x"EFA3",
			x"0000" when x"EFA4",
			x"0000" when x"EFA5",
			x"0000" when x"EFA6",
			x"0000" when x"EFA7",
			x"0000" when x"EFA8",
			x"0000" when x"EFA9",
			x"0000" when x"EFAA",
			x"0000" when x"EFAB",
			x"0000" when x"EFAC",
			x"0000" when x"EFAD",
			x"0000" when x"EFAE",
			x"0000" when x"EFAF",
			x"0000" when x"EFB0",
			x"0000" when x"EFB1",
			x"0000" when x"EFB2",
			x"0000" when x"EFB3",
			x"0000" when x"EFB4",
			x"0000" when x"EFB5",
			x"0000" when x"EFB6",
			x"0000" when x"EFB7",
			x"0000" when x"EFB8",
			x"0000" when x"EFB9",
			x"0000" when x"EFBA",
			x"0000" when x"EFBB",
			x"0000" when x"EFBC",
			x"0000" when x"EFBD",
			x"0000" when x"EFBE",
			x"0000" when x"EFBF",
			x"0000" when x"EFC0",
			x"0000" when x"EFC1",
			x"0000" when x"EFC2",
			x"0000" when x"EFC3",
			x"0000" when x"EFC4",
			x"0000" when x"EFC5",
			x"0000" when x"EFC6",
			x"0000" when x"EFC7",
			x"0000" when x"EFC8",
			x"0000" when x"EFC9",
			x"0000" when x"EFCA",
			x"0000" when x"EFCB",
			x"0000" when x"EFCC",
			x"0000" when x"EFCD",
			x"0000" when x"EFCE",
			x"0000" when x"EFCF",
			x"0000" when x"EFD0",
			x"0000" when x"EFD1",
			x"0000" when x"EFD2",
			x"0000" when x"EFD3",
			x"0000" when x"EFD4",
			x"0000" when x"EFD5",
			x"0000" when x"EFD6",
			x"0000" when x"EFD7",
			x"0000" when x"EFD8",
			x"0000" when x"EFD9",
			x"0000" when x"EFDA",
			x"0000" when x"EFDB",
			x"0000" when x"EFDC",
			x"0000" when x"EFDD",
			x"0000" when x"EFDE",
			x"0000" when x"EFDF",
			x"0000" when x"EFE0",
			x"0000" when x"EFE1",
			x"0000" when x"EFE2",
			x"0000" when x"EFE3",
			x"0000" when x"EFE4",
			x"0000" when x"EFE5",
			x"0000" when x"EFE6",
			x"0000" when x"EFE7",
			x"0000" when x"EFE8",
			x"0000" when x"EFE9",
			x"0000" when x"EFEA",
			x"0000" when x"EFEB",
			x"0000" when x"EFEC",
			x"0000" when x"EFED",
			x"0000" when x"EFEE",
			x"0000" when x"EFEF",
			x"0000" when x"EFF0",
			x"0000" when x"EFF1",
			x"0000" when x"EFF2",
			x"0000" when x"EFF3",
			x"0000" when x"EFF4",
			x"0000" when x"EFF5",
			x"0000" when x"EFF6",
			x"0000" when x"EFF7",
			x"0000" when x"EFF8",
			x"0000" when x"EFF9",
			x"0000" when x"EFFA",
			x"0000" when x"EFFB",
			x"0000" when x"EFFC",
			x"0000" when x"EFFD",
			x"0000" when x"EFFE",
			x"0000" when x"EFFF",
			x"0000" when x"F000",
			x"0000" when x"F001",
			x"0000" when x"F002",
			x"0000" when x"F003",
			x"0000" when x"F004",
			x"0000" when x"F005",
			x"0000" when x"F006",
			x"0000" when x"F007",
			x"0000" when x"F008",
			x"0000" when x"F009",
			x"0000" when x"F00A",
			x"0000" when x"F00B",
			x"0000" when x"F00C",
			x"0000" when x"F00D",
			x"0000" when x"F00E",
			x"0000" when x"F00F",
			x"0000" when x"F010",
			x"0000" when x"F011",
			x"0000" when x"F012",
			x"0000" when x"F013",
			x"0000" when x"F014",
			x"0000" when x"F015",
			x"0000" when x"F016",
			x"0000" when x"F017",
			x"0000" when x"F018",
			x"0000" when x"F019",
			x"0000" when x"F01A",
			x"0000" when x"F01B",
			x"0000" when x"F01C",
			x"0000" when x"F01D",
			x"0000" when x"F01E",
			x"0000" when x"F01F",
			x"0000" when x"F020",
			x"0000" when x"F021",
			x"0000" when x"F022",
			x"0000" when x"F023",
			x"0000" when x"F024",
			x"0000" when x"F025",
			x"0000" when x"F026",
			x"0000" when x"F027",
			x"0000" when x"F028",
			x"0000" when x"F029",
			x"0000" when x"F02A",
			x"0000" when x"F02B",
			x"0000" when x"F02C",
			x"0000" when x"F02D",
			x"0000" when x"F02E",
			x"0000" when x"F02F",
			x"0000" when x"F030",
			x"0000" when x"F031",
			x"0000" when x"F032",
			x"0000" when x"F033",
			x"0000" when x"F034",
			x"0000" when x"F035",
			x"0000" when x"F036",
			x"0000" when x"F037",
			x"0000" when x"F038",
			x"0000" when x"F039",
			x"0000" when x"F03A",
			x"0000" when x"F03B",
			x"0000" when x"F03C",
			x"0000" when x"F03D",
			x"0000" when x"F03E",
			x"0000" when x"F03F",
			x"0000" when x"F040",
			x"0000" when x"F041",
			x"0000" when x"F042",
			x"0000" when x"F043",
			x"0000" when x"F044",
			x"0000" when x"F045",
			x"0000" when x"F046",
			x"0000" when x"F047",
			x"0000" when x"F048",
			x"0000" when x"F049",
			x"0000" when x"F04A",
			x"0000" when x"F04B",
			x"0000" when x"F04C",
			x"0000" when x"F04D",
			x"0000" when x"F04E",
			x"0000" when x"F04F",
			x"0000" when x"F050",
			x"0000" when x"F051",
			x"0000" when x"F052",
			x"0000" when x"F053",
			x"0000" when x"F054",
			x"0000" when x"F055",
			x"0000" when x"F056",
			x"0000" when x"F057",
			x"0000" when x"F058",
			x"0000" when x"F059",
			x"0000" when x"F05A",
			x"0000" when x"F05B",
			x"0000" when x"F05C",
			x"0000" when x"F05D",
			x"0000" when x"F05E",
			x"0000" when x"F05F",
			x"0000" when x"F060",
			x"0000" when x"F061",
			x"0000" when x"F062",
			x"0000" when x"F063",
			x"0000" when x"F064",
			x"0000" when x"F065",
			x"0000" when x"F066",
			x"0000" when x"F067",
			x"0000" when x"F068",
			x"0000" when x"F069",
			x"0000" when x"F06A",
			x"0000" when x"F06B",
			x"0000" when x"F06C",
			x"0000" when x"F06D",
			x"0000" when x"F06E",
			x"0000" when x"F06F",
			x"0000" when x"F070",
			x"0000" when x"F071",
			x"0000" when x"F072",
			x"0000" when x"F073",
			x"0000" when x"F074",
			x"0000" when x"F075",
			x"0000" when x"F076",
			x"0000" when x"F077",
			x"0000" when x"F078",
			x"0000" when x"F079",
			x"0000" when x"F07A",
			x"0000" when x"F07B",
			x"0000" when x"F07C",
			x"0000" when x"F07D",
			x"0000" when x"F07E",
			x"0000" when x"F07F",
			x"0000" when x"F080",
			x"0000" when x"F081",
			x"0000" when x"F082",
			x"0000" when x"F083",
			x"0000" when x"F084",
			x"0000" when x"F085",
			x"0000" when x"F086",
			x"0000" when x"F087",
			x"0000" when x"F088",
			x"0000" when x"F089",
			x"0000" when x"F08A",
			x"0000" when x"F08B",
			x"0000" when x"F08C",
			x"0000" when x"F08D",
			x"0000" when x"F08E",
			x"0000" when x"F08F",
			x"0000" when x"F090",
			x"0000" when x"F091",
			x"0000" when x"F092",
			x"0000" when x"F093",
			x"0000" when x"F094",
			x"0000" when x"F095",
			x"0000" when x"F096",
			x"0000" when x"F097",
			x"0000" when x"F098",
			x"0000" when x"F099",
			x"0000" when x"F09A",
			x"0000" when x"F09B",
			x"0000" when x"F09C",
			x"0000" when x"F09D",
			x"0000" when x"F09E",
			x"0000" when x"F09F",
			x"0000" when x"F0A0",
			x"0000" when x"F0A1",
			x"0000" when x"F0A2",
			x"0000" when x"F0A3",
			x"0000" when x"F0A4",
			x"0000" when x"F0A5",
			x"0000" when x"F0A6",
			x"0000" when x"F0A7",
			x"0000" when x"F0A8",
			x"0000" when x"F0A9",
			x"0000" when x"F0AA",
			x"0000" when x"F0AB",
			x"0000" when x"F0AC",
			x"0000" when x"F0AD",
			x"0000" when x"F0AE",
			x"0000" when x"F0AF",
			x"0000" when x"F0B0",
			x"0000" when x"F0B1",
			x"0000" when x"F0B2",
			x"0000" when x"F0B3",
			x"0000" when x"F0B4",
			x"0000" when x"F0B5",
			x"0000" when x"F0B6",
			x"0000" when x"F0B7",
			x"0000" when x"F0B8",
			x"0000" when x"F0B9",
			x"0000" when x"F0BA",
			x"0000" when x"F0BB",
			x"0000" when x"F0BC",
			x"0000" when x"F0BD",
			x"0000" when x"F0BE",
			x"0000" when x"F0BF",
			x"0000" when x"F0C0",
			x"0000" when x"F0C1",
			x"0000" when x"F0C2",
			x"0000" when x"F0C3",
			x"0000" when x"F0C4",
			x"0000" when x"F0C5",
			x"0000" when x"F0C6",
			x"0000" when x"F0C7",
			x"0000" when x"F0C8",
			x"0000" when x"F0C9",
			x"0000" when x"F0CA",
			x"0000" when x"F0CB",
			x"0000" when x"F0CC",
			x"0000" when x"F0CD",
			x"0000" when x"F0CE",
			x"0000" when x"F0CF",
			x"0000" when x"F0D0",
			x"0000" when x"F0D1",
			x"0000" when x"F0D2",
			x"0000" when x"F0D3",
			x"0000" when x"F0D4",
			x"0000" when x"F0D5",
			x"0000" when x"F0D6",
			x"0000" when x"F0D7",
			x"0000" when x"F0D8",
			x"0000" when x"F0D9",
			x"0000" when x"F0DA",
			x"0000" when x"F0DB",
			x"0000" when x"F0DC",
			x"0000" when x"F0DD",
			x"0000" when x"F0DE",
			x"0000" when x"F0DF",
			x"0000" when x"F0E0",
			x"0000" when x"F0E1",
			x"0000" when x"F0E2",
			x"0000" when x"F0E3",
			x"0000" when x"F0E4",
			x"0000" when x"F0E5",
			x"0000" when x"F0E6",
			x"0000" when x"F0E7",
			x"0000" when x"F0E8",
			x"0000" when x"F0E9",
			x"0000" when x"F0EA",
			x"0000" when x"F0EB",
			x"0000" when x"F0EC",
			x"0000" when x"F0ED",
			x"0000" when x"F0EE",
			x"0000" when x"F0EF",
			x"0000" when x"F0F0",
			x"0000" when x"F0F1",
			x"0000" when x"F0F2",
			x"0000" when x"F0F3",
			x"0000" when x"F0F4",
			x"0000" when x"F0F5",
			x"0000" when x"F0F6",
			x"0000" when x"F0F7",
			x"0000" when x"F0F8",
			x"0000" when x"F0F9",
			x"0000" when x"F0FA",
			x"0000" when x"F0FB",
			x"0000" when x"F0FC",
			x"0000" when x"F0FD",
			x"0000" when x"F0FE",
			x"0000" when x"F0FF",
			x"0000" when x"F100",
			x"0000" when x"F101",
			x"0000" when x"F102",
			x"0000" when x"F103",
			x"0000" when x"F104",
			x"0000" when x"F105",
			x"0000" when x"F106",
			x"0000" when x"F107",
			x"0000" when x"F108",
			x"0000" when x"F109",
			x"0000" when x"F10A",
			x"0000" when x"F10B",
			x"0000" when x"F10C",
			x"0000" when x"F10D",
			x"0000" when x"F10E",
			x"0000" when x"F10F",
			x"0000" when x"F110",
			x"0000" when x"F111",
			x"0000" when x"F112",
			x"0000" when x"F113",
			x"0000" when x"F114",
			x"0000" when x"F115",
			x"0000" when x"F116",
			x"0000" when x"F117",
			x"0000" when x"F118",
			x"0000" when x"F119",
			x"0000" when x"F11A",
			x"0000" when x"F11B",
			x"0000" when x"F11C",
			x"0000" when x"F11D",
			x"0000" when x"F11E",
			x"0000" when x"F11F",
			x"0000" when x"F120",
			x"0000" when x"F121",
			x"0000" when x"F122",
			x"0000" when x"F123",
			x"0000" when x"F124",
			x"0000" when x"F125",
			x"0000" when x"F126",
			x"0000" when x"F127",
			x"0000" when x"F128",
			x"0000" when x"F129",
			x"0000" when x"F12A",
			x"0000" when x"F12B",
			x"0000" when x"F12C",
			x"0000" when x"F12D",
			x"0000" when x"F12E",
			x"0000" when x"F12F",
			x"0000" when x"F130",
			x"0000" when x"F131",
			x"0000" when x"F132",
			x"0000" when x"F133",
			x"0000" when x"F134",
			x"0000" when x"F135",
			x"0000" when x"F136",
			x"0000" when x"F137",
			x"0000" when x"F138",
			x"0000" when x"F139",
			x"0000" when x"F13A",
			x"0000" when x"F13B",
			x"0000" when x"F13C",
			x"0000" when x"F13D",
			x"0000" when x"F13E",
			x"0000" when x"F13F",
			x"0000" when x"F140",
			x"0000" when x"F141",
			x"0000" when x"F142",
			x"0000" when x"F143",
			x"0000" when x"F144",
			x"0000" when x"F145",
			x"0000" when x"F146",
			x"0000" when x"F147",
			x"0000" when x"F148",
			x"0000" when x"F149",
			x"0000" when x"F14A",
			x"0000" when x"F14B",
			x"0000" when x"F14C",
			x"0000" when x"F14D",
			x"0000" when x"F14E",
			x"0000" when x"F14F",
			x"0000" when x"F150",
			x"0000" when x"F151",
			x"0000" when x"F152",
			x"0000" when x"F153",
			x"0000" when x"F154",
			x"0000" when x"F155",
			x"0000" when x"F156",
			x"0000" when x"F157",
			x"0000" when x"F158",
			x"0000" when x"F159",
			x"0000" when x"F15A",
			x"0000" when x"F15B",
			x"0000" when x"F15C",
			x"0000" when x"F15D",
			x"0000" when x"F15E",
			x"0000" when x"F15F",
			x"0000" when x"F160",
			x"0000" when x"F161",
			x"0000" when x"F162",
			x"0000" when x"F163",
			x"0000" when x"F164",
			x"0000" when x"F165",
			x"0000" when x"F166",
			x"0000" when x"F167",
			x"0000" when x"F168",
			x"0000" when x"F169",
			x"0000" when x"F16A",
			x"0000" when x"F16B",
			x"0000" when x"F16C",
			x"0000" when x"F16D",
			x"0000" when x"F16E",
			x"0000" when x"F16F",
			x"0000" when x"F170",
			x"0000" when x"F171",
			x"0000" when x"F172",
			x"0000" when x"F173",
			x"0000" when x"F174",
			x"0000" when x"F175",
			x"0000" when x"F176",
			x"0000" when x"F177",
			x"0000" when x"F178",
			x"0000" when x"F179",
			x"0000" when x"F17A",
			x"0000" when x"F17B",
			x"0000" when x"F17C",
			x"0000" when x"F17D",
			x"0000" when x"F17E",
			x"0000" when x"F17F",
			x"0000" when x"F180",
			x"0000" when x"F181",
			x"0000" when x"F182",
			x"0000" when x"F183",
			x"0000" when x"F184",
			x"0000" when x"F185",
			x"0000" when x"F186",
			x"0000" when x"F187",
			x"0000" when x"F188",
			x"0000" when x"F189",
			x"0000" when x"F18A",
			x"0000" when x"F18B",
			x"0000" when x"F18C",
			x"0000" when x"F18D",
			x"0000" when x"F18E",
			x"0000" when x"F18F",
			x"0000" when x"F190",
			x"0000" when x"F191",
			x"0000" when x"F192",
			x"0000" when x"F193",
			x"0000" when x"F194",
			x"0000" when x"F195",
			x"0000" when x"F196",
			x"0000" when x"F197",
			x"0000" when x"F198",
			x"0000" when x"F199",
			x"0000" when x"F19A",
			x"0000" when x"F19B",
			x"0000" when x"F19C",
			x"0000" when x"F19D",
			x"0000" when x"F19E",
			x"0000" when x"F19F",
			x"0000" when x"F1A0",
			x"0000" when x"F1A1",
			x"0000" when x"F1A2",
			x"0000" when x"F1A3",
			x"0000" when x"F1A4",
			x"0000" when x"F1A5",
			x"0000" when x"F1A6",
			x"0000" when x"F1A7",
			x"0000" when x"F1A8",
			x"0000" when x"F1A9",
			x"0000" when x"F1AA",
			x"0000" when x"F1AB",
			x"0000" when x"F1AC",
			x"0000" when x"F1AD",
			x"0000" when x"F1AE",
			x"0000" when x"F1AF",
			x"0000" when x"F1B0",
			x"0000" when x"F1B1",
			x"0000" when x"F1B2",
			x"0000" when x"F1B3",
			x"0000" when x"F1B4",
			x"0000" when x"F1B5",
			x"0000" when x"F1B6",
			x"0000" when x"F1B7",
			x"0000" when x"F1B8",
			x"0000" when x"F1B9",
			x"0000" when x"F1BA",
			x"0000" when x"F1BB",
			x"0000" when x"F1BC",
			x"0000" when x"F1BD",
			x"0000" when x"F1BE",
			x"0000" when x"F1BF",
			x"0000" when x"F1C0",
			x"0000" when x"F1C1",
			x"0000" when x"F1C2",
			x"0000" when x"F1C3",
			x"0000" when x"F1C4",
			x"0000" when x"F1C5",
			x"0000" when x"F1C6",
			x"0000" when x"F1C7",
			x"0000" when x"F1C8",
			x"0000" when x"F1C9",
			x"0000" when x"F1CA",
			x"0000" when x"F1CB",
			x"0000" when x"F1CC",
			x"0000" when x"F1CD",
			x"0000" when x"F1CE",
			x"0000" when x"F1CF",
			x"0000" when x"F1D0",
			x"0000" when x"F1D1",
			x"0000" when x"F1D2",
			x"0000" when x"F1D3",
			x"0000" when x"F1D4",
			x"0000" when x"F1D5",
			x"0000" when x"F1D6",
			x"0000" when x"F1D7",
			x"0000" when x"F1D8",
			x"0000" when x"F1D9",
			x"0000" when x"F1DA",
			x"0000" when x"F1DB",
			x"0000" when x"F1DC",
			x"0000" when x"F1DD",
			x"0000" when x"F1DE",
			x"0000" when x"F1DF",
			x"0000" when x"F1E0",
			x"0000" when x"F1E1",
			x"0000" when x"F1E2",
			x"0000" when x"F1E3",
			x"0000" when x"F1E4",
			x"0000" when x"F1E5",
			x"0000" when x"F1E6",
			x"0000" when x"F1E7",
			x"0000" when x"F1E8",
			x"0000" when x"F1E9",
			x"0000" when x"F1EA",
			x"0000" when x"F1EB",
			x"0000" when x"F1EC",
			x"0000" when x"F1ED",
			x"0000" when x"F1EE",
			x"0000" when x"F1EF",
			x"0000" when x"F1F0",
			x"0000" when x"F1F1",
			x"0000" when x"F1F2",
			x"0000" when x"F1F3",
			x"0000" when x"F1F4",
			x"0000" when x"F1F5",
			x"0000" when x"F1F6",
			x"0000" when x"F1F7",
			x"0000" when x"F1F8",
			x"0000" when x"F1F9",
			x"0000" when x"F1FA",
			x"0000" when x"F1FB",
			x"0000" when x"F1FC",
			x"0000" when x"F1FD",
			x"0000" when x"F1FE",
			x"0000" when x"F1FF",
			x"0000" when x"F200",
			x"0000" when x"F201",
			x"0000" when x"F202",
			x"0000" when x"F203",
			x"0000" when x"F204",
			x"0000" when x"F205",
			x"0000" when x"F206",
			x"0000" when x"F207",
			x"0000" when x"F208",
			x"0000" when x"F209",
			x"0000" when x"F20A",
			x"0000" when x"F20B",
			x"0000" when x"F20C",
			x"0000" when x"F20D",
			x"0000" when x"F20E",
			x"0000" when x"F20F",
			x"0000" when x"F210",
			x"0000" when x"F211",
			x"0000" when x"F212",
			x"0000" when x"F213",
			x"0000" when x"F214",
			x"0000" when x"F215",
			x"0000" when x"F216",
			x"0000" when x"F217",
			x"0000" when x"F218",
			x"0000" when x"F219",
			x"0000" when x"F21A",
			x"0000" when x"F21B",
			x"0000" when x"F21C",
			x"0000" when x"F21D",
			x"0000" when x"F21E",
			x"0000" when x"F21F",
			x"0000" when x"F220",
			x"0000" when x"F221",
			x"0000" when x"F222",
			x"0000" when x"F223",
			x"0000" when x"F224",
			x"0000" when x"F225",
			x"0000" when x"F226",
			x"0000" when x"F227",
			x"0000" when x"F228",
			x"0000" when x"F229",
			x"0000" when x"F22A",
			x"0000" when x"F22B",
			x"0000" when x"F22C",
			x"0000" when x"F22D",
			x"0000" when x"F22E",
			x"0000" when x"F22F",
			x"0000" when x"F230",
			x"0000" when x"F231",
			x"0000" when x"F232",
			x"0000" when x"F233",
			x"0000" when x"F234",
			x"0000" when x"F235",
			x"0000" when x"F236",
			x"0000" when x"F237",
			x"0000" when x"F238",
			x"0000" when x"F239",
			x"0000" when x"F23A",
			x"0000" when x"F23B",
			x"0000" when x"F23C",
			x"0000" when x"F23D",
			x"0000" when x"F23E",
			x"0000" when x"F23F",
			x"0000" when x"F240",
			x"0000" when x"F241",
			x"0000" when x"F242",
			x"0000" when x"F243",
			x"0000" when x"F244",
			x"0000" when x"F245",
			x"0000" when x"F246",
			x"0000" when x"F247",
			x"0000" when x"F248",
			x"0000" when x"F249",
			x"0000" when x"F24A",
			x"0000" when x"F24B",
			x"0000" when x"F24C",
			x"0000" when x"F24D",
			x"0000" when x"F24E",
			x"0000" when x"F24F",
			x"0000" when x"F250",
			x"0000" when x"F251",
			x"0000" when x"F252",
			x"0000" when x"F253",
			x"0000" when x"F254",
			x"0000" when x"F255",
			x"0000" when x"F256",
			x"0000" when x"F257",
			x"0000" when x"F258",
			x"0000" when x"F259",
			x"0000" when x"F25A",
			x"0000" when x"F25B",
			x"0000" when x"F25C",
			x"0000" when x"F25D",
			x"0000" when x"F25E",
			x"0000" when x"F25F",
			x"0000" when x"F260",
			x"0000" when x"F261",
			x"0000" when x"F262",
			x"0000" when x"F263",
			x"0000" when x"F264",
			x"0000" when x"F265",
			x"0000" when x"F266",
			x"0000" when x"F267",
			x"0000" when x"F268",
			x"0000" when x"F269",
			x"0000" when x"F26A",
			x"0000" when x"F26B",
			x"0000" when x"F26C",
			x"0000" when x"F26D",
			x"0000" when x"F26E",
			x"0000" when x"F26F",
			x"0000" when x"F270",
			x"0000" when x"F271",
			x"0000" when x"F272",
			x"0000" when x"F273",
			x"0000" when x"F274",
			x"0000" when x"F275",
			x"0000" when x"F276",
			x"0000" when x"F277",
			x"0000" when x"F278",
			x"0000" when x"F279",
			x"0000" when x"F27A",
			x"0000" when x"F27B",
			x"0000" when x"F27C",
			x"0000" when x"F27D",
			x"0000" when x"F27E",
			x"0000" when x"F27F",
			x"0000" when x"F280",
			x"0000" when x"F281",
			x"0000" when x"F282",
			x"0000" when x"F283",
			x"0000" when x"F284",
			x"0000" when x"F285",
			x"0000" when x"F286",
			x"0000" when x"F287",
			x"0000" when x"F288",
			x"0000" when x"F289",
			x"0000" when x"F28A",
			x"0000" when x"F28B",
			x"0000" when x"F28C",
			x"0000" when x"F28D",
			x"0000" when x"F28E",
			x"0000" when x"F28F",
			x"0000" when x"F290",
			x"0000" when x"F291",
			x"0000" when x"F292",
			x"0000" when x"F293",
			x"0000" when x"F294",
			x"0000" when x"F295",
			x"0000" when x"F296",
			x"0000" when x"F297",
			x"0000" when x"F298",
			x"0000" when x"F299",
			x"0000" when x"F29A",
			x"0000" when x"F29B",
			x"0000" when x"F29C",
			x"0000" when x"F29D",
			x"0000" when x"F29E",
			x"0000" when x"F29F",
			x"0000" when x"F2A0",
			x"0000" when x"F2A1",
			x"0000" when x"F2A2",
			x"0000" when x"F2A3",
			x"0000" when x"F2A4",
			x"0000" when x"F2A5",
			x"0000" when x"F2A6",
			x"0000" when x"F2A7",
			x"0000" when x"F2A8",
			x"0000" when x"F2A9",
			x"0000" when x"F2AA",
			x"0000" when x"F2AB",
			x"0000" when x"F2AC",
			x"0000" when x"F2AD",
			x"0000" when x"F2AE",
			x"0000" when x"F2AF",
			x"0000" when x"F2B0",
			x"0000" when x"F2B1",
			x"0000" when x"F2B2",
			x"0000" when x"F2B3",
			x"0000" when x"F2B4",
			x"0000" when x"F2B5",
			x"0000" when x"F2B6",
			x"0000" when x"F2B7",
			x"0000" when x"F2B8",
			x"0000" when x"F2B9",
			x"0000" when x"F2BA",
			x"0000" when x"F2BB",
			x"0000" when x"F2BC",
			x"0000" when x"F2BD",
			x"0000" when x"F2BE",
			x"0000" when x"F2BF",
			x"0000" when x"F2C0",
			x"0000" when x"F2C1",
			x"0000" when x"F2C2",
			x"0000" when x"F2C3",
			x"0000" when x"F2C4",
			x"0000" when x"F2C5",
			x"0000" when x"F2C6",
			x"0000" when x"F2C7",
			x"0000" when x"F2C8",
			x"0000" when x"F2C9",
			x"0000" when x"F2CA",
			x"0000" when x"F2CB",
			x"0000" when x"F2CC",
			x"0000" when x"F2CD",
			x"0000" when x"F2CE",
			x"0000" when x"F2CF",
			x"0000" when x"F2D0",
			x"0000" when x"F2D1",
			x"0000" when x"F2D2",
			x"0000" when x"F2D3",
			x"0000" when x"F2D4",
			x"0000" when x"F2D5",
			x"0000" when x"F2D6",
			x"0000" when x"F2D7",
			x"0000" when x"F2D8",
			x"0000" when x"F2D9",
			x"0000" when x"F2DA",
			x"0000" when x"F2DB",
			x"0000" when x"F2DC",
			x"0000" when x"F2DD",
			x"0000" when x"F2DE",
			x"0000" when x"F2DF",
			x"0000" when x"F2E0",
			x"0000" when x"F2E1",
			x"0000" when x"F2E2",
			x"0000" when x"F2E3",
			x"0000" when x"F2E4",
			x"0000" when x"F2E5",
			x"0000" when x"F2E6",
			x"0000" when x"F2E7",
			x"0000" when x"F2E8",
			x"0000" when x"F2E9",
			x"0000" when x"F2EA",
			x"0000" when x"F2EB",
			x"0000" when x"F2EC",
			x"0000" when x"F2ED",
			x"0000" when x"F2EE",
			x"0000" when x"F2EF",
			x"0000" when x"F2F0",
			x"0000" when x"F2F1",
			x"0000" when x"F2F2",
			x"0000" when x"F2F3",
			x"0000" when x"F2F4",
			x"0000" when x"F2F5",
			x"0000" when x"F2F6",
			x"0000" when x"F2F7",
			x"0000" when x"F2F8",
			x"0000" when x"F2F9",
			x"0000" when x"F2FA",
			x"0000" when x"F2FB",
			x"0000" when x"F2FC",
			x"0000" when x"F2FD",
			x"0000" when x"F2FE",
			x"0000" when x"F2FF",
			x"0000" when x"F300",
			x"0000" when x"F301",
			x"0000" when x"F302",
			x"0000" when x"F303",
			x"0000" when x"F304",
			x"0000" when x"F305",
			x"0000" when x"F306",
			x"0000" when x"F307",
			x"0000" when x"F308",
			x"0000" when x"F309",
			x"0000" when x"F30A",
			x"0000" when x"F30B",
			x"0000" when x"F30C",
			x"0000" when x"F30D",
			x"0000" when x"F30E",
			x"0000" when x"F30F",
			x"0000" when x"F310",
			x"0000" when x"F311",
			x"0000" when x"F312",
			x"0000" when x"F313",
			x"0000" when x"F314",
			x"0000" when x"F315",
			x"0000" when x"F316",
			x"0000" when x"F317",
			x"0000" when x"F318",
			x"0000" when x"F319",
			x"0000" when x"F31A",
			x"0000" when x"F31B",
			x"0000" when x"F31C",
			x"0000" when x"F31D",
			x"0000" when x"F31E",
			x"0000" when x"F31F",
			x"0000" when x"F320",
			x"0000" when x"F321",
			x"0000" when x"F322",
			x"0000" when x"F323",
			x"0000" when x"F324",
			x"0000" when x"F325",
			x"0000" when x"F326",
			x"0000" when x"F327",
			x"0000" when x"F328",
			x"0000" when x"F329",
			x"0000" when x"F32A",
			x"0000" when x"F32B",
			x"0000" when x"F32C",
			x"0000" when x"F32D",
			x"0000" when x"F32E",
			x"0000" when x"F32F",
			x"0000" when x"F330",
			x"0000" when x"F331",
			x"0000" when x"F332",
			x"0000" when x"F333",
			x"0000" when x"F334",
			x"0000" when x"F335",
			x"0000" when x"F336",
			x"0000" when x"F337",
			x"0000" when x"F338",
			x"0000" when x"F339",
			x"0000" when x"F33A",
			x"0000" when x"F33B",
			x"0000" when x"F33C",
			x"0000" when x"F33D",
			x"0000" when x"F33E",
			x"0000" when x"F33F",
			x"0000" when x"F340",
			x"0000" when x"F341",
			x"0000" when x"F342",
			x"0000" when x"F343",
			x"0000" when x"F344",
			x"0000" when x"F345",
			x"0000" when x"F346",
			x"0000" when x"F347",
			x"0000" when x"F348",
			x"0000" when x"F349",
			x"0000" when x"F34A",
			x"0000" when x"F34B",
			x"0000" when x"F34C",
			x"0000" when x"F34D",
			x"0000" when x"F34E",
			x"0000" when x"F34F",
			x"0000" when x"F350",
			x"0000" when x"F351",
			x"0000" when x"F352",
			x"0000" when x"F353",
			x"0000" when x"F354",
			x"0000" when x"F355",
			x"0000" when x"F356",
			x"0000" when x"F357",
			x"0000" when x"F358",
			x"0000" when x"F359",
			x"0000" when x"F35A",
			x"0000" when x"F35B",
			x"0000" when x"F35C",
			x"0000" when x"F35D",
			x"0000" when x"F35E",
			x"0000" when x"F35F",
			x"0000" when x"F360",
			x"0000" when x"F361",
			x"0000" when x"F362",
			x"0000" when x"F363",
			x"0000" when x"F364",
			x"0000" when x"F365",
			x"0000" when x"F366",
			x"0000" when x"F367",
			x"0000" when x"F368",
			x"0000" when x"F369",
			x"0000" when x"F36A",
			x"0000" when x"F36B",
			x"0000" when x"F36C",
			x"0000" when x"F36D",
			x"0000" when x"F36E",
			x"0000" when x"F36F",
			x"0000" when x"F370",
			x"0000" when x"F371",
			x"0000" when x"F372",
			x"0000" when x"F373",
			x"0000" when x"F374",
			x"0000" when x"F375",
			x"0000" when x"F376",
			x"0000" when x"F377",
			x"0000" when x"F378",
			x"0000" when x"F379",
			x"0000" when x"F37A",
			x"0000" when x"F37B",
			x"0000" when x"F37C",
			x"0000" when x"F37D",
			x"0000" when x"F37E",
			x"0000" when x"F37F",
			x"0000" when x"F380",
			x"0000" when x"F381",
			x"0000" when x"F382",
			x"0000" when x"F383",
			x"0000" when x"F384",
			x"0000" when x"F385",
			x"0000" when x"F386",
			x"0000" when x"F387",
			x"0000" when x"F388",
			x"0000" when x"F389",
			x"0000" when x"F38A",
			x"0000" when x"F38B",
			x"0000" when x"F38C",
			x"0000" when x"F38D",
			x"0000" when x"F38E",
			x"0000" when x"F38F",
			x"0000" when x"F390",
			x"0000" when x"F391",
			x"0000" when x"F392",
			x"0000" when x"F393",
			x"0000" when x"F394",
			x"0000" when x"F395",
			x"0000" when x"F396",
			x"0000" when x"F397",
			x"0000" when x"F398",
			x"0000" when x"F399",
			x"0000" when x"F39A",
			x"0000" when x"F39B",
			x"0000" when x"F39C",
			x"0000" when x"F39D",
			x"0000" when x"F39E",
			x"0000" when x"F39F",
			x"0000" when x"F3A0",
			x"0000" when x"F3A1",
			x"0000" when x"F3A2",
			x"0000" when x"F3A3",
			x"0000" when x"F3A4",
			x"0000" when x"F3A5",
			x"0000" when x"F3A6",
			x"0000" when x"F3A7",
			x"0000" when x"F3A8",
			x"0000" when x"F3A9",
			x"0000" when x"F3AA",
			x"0000" when x"F3AB",
			x"0000" when x"F3AC",
			x"0000" when x"F3AD",
			x"0000" when x"F3AE",
			x"0000" when x"F3AF",
			x"0000" when x"F3B0",
			x"0000" when x"F3B1",
			x"0000" when x"F3B2",
			x"0000" when x"F3B3",
			x"0000" when x"F3B4",
			x"0000" when x"F3B5",
			x"0000" when x"F3B6",
			x"0000" when x"F3B7",
			x"0000" when x"F3B8",
			x"0000" when x"F3B9",
			x"0000" when x"F3BA",
			x"0000" when x"F3BB",
			x"0000" when x"F3BC",
			x"0000" when x"F3BD",
			x"0000" when x"F3BE",
			x"0000" when x"F3BF",
			x"0000" when x"F3C0",
			x"0000" when x"F3C1",
			x"0000" when x"F3C2",
			x"0000" when x"F3C3",
			x"0000" when x"F3C4",
			x"0000" when x"F3C5",
			x"0000" when x"F3C6",
			x"0000" when x"F3C7",
			x"0000" when x"F3C8",
			x"0000" when x"F3C9",
			x"0000" when x"F3CA",
			x"0000" when x"F3CB",
			x"0000" when x"F3CC",
			x"0000" when x"F3CD",
			x"0000" when x"F3CE",
			x"0000" when x"F3CF",
			x"0000" when x"F3D0",
			x"0000" when x"F3D1",
			x"0000" when x"F3D2",
			x"0000" when x"F3D3",
			x"0000" when x"F3D4",
			x"0000" when x"F3D5",
			x"0000" when x"F3D6",
			x"0000" when x"F3D7",
			x"0000" when x"F3D8",
			x"0000" when x"F3D9",
			x"0000" when x"F3DA",
			x"0000" when x"F3DB",
			x"0000" when x"F3DC",
			x"0000" when x"F3DD",
			x"0000" when x"F3DE",
			x"0000" when x"F3DF",
			x"0000" when x"F3E0",
			x"0000" when x"F3E1",
			x"0000" when x"F3E2",
			x"0000" when x"F3E3",
			x"0000" when x"F3E4",
			x"0000" when x"F3E5",
			x"0000" when x"F3E6",
			x"0000" when x"F3E7",
			x"0000" when x"F3E8",
			x"0000" when x"F3E9",
			x"0000" when x"F3EA",
			x"0000" when x"F3EB",
			x"0000" when x"F3EC",
			x"0000" when x"F3ED",
			x"0000" when x"F3EE",
			x"0000" when x"F3EF",
			x"0000" when x"F3F0",
			x"0000" when x"F3F1",
			x"0000" when x"F3F2",
			x"0000" when x"F3F3",
			x"0000" when x"F3F4",
			x"0000" when x"F3F5",
			x"0000" when x"F3F6",
			x"0000" when x"F3F7",
			x"0000" when x"F3F8",
			x"0000" when x"F3F9",
			x"0000" when x"F3FA",
			x"0000" when x"F3FB",
			x"0000" when x"F3FC",
			x"0000" when x"F3FD",
			x"0000" when x"F3FE",
			x"0000" when x"F3FF",
			x"0000" when x"F400",
			x"0000" when x"F401",
			x"0000" when x"F402",
			x"0000" when x"F403",
			x"0000" when x"F404",
			x"0000" when x"F405",
			x"0000" when x"F406",
			x"0000" when x"F407",
			x"0000" when x"F408",
			x"0000" when x"F409",
			x"0000" when x"F40A",
			x"0000" when x"F40B",
			x"0000" when x"F40C",
			x"0000" when x"F40D",
			x"0000" when x"F40E",
			x"0000" when x"F40F",
			x"0000" when x"F410",
			x"0000" when x"F411",
			x"0000" when x"F412",
			x"0000" when x"F413",
			x"0000" when x"F414",
			x"0000" when x"F415",
			x"0000" when x"F416",
			x"0000" when x"F417",
			x"0000" when x"F418",
			x"0000" when x"F419",
			x"0000" when x"F41A",
			x"0000" when x"F41B",
			x"0000" when x"F41C",
			x"0000" when x"F41D",
			x"0000" when x"F41E",
			x"0000" when x"F41F",
			x"0000" when x"F420",
			x"0000" when x"F421",
			x"0000" when x"F422",
			x"0000" when x"F423",
			x"0000" when x"F424",
			x"0000" when x"F425",
			x"0000" when x"F426",
			x"0000" when x"F427",
			x"0000" when x"F428",
			x"0000" when x"F429",
			x"0000" when x"F42A",
			x"0000" when x"F42B",
			x"0000" when x"F42C",
			x"0000" when x"F42D",
			x"0000" when x"F42E",
			x"0000" when x"F42F",
			x"0000" when x"F430",
			x"0000" when x"F431",
			x"0000" when x"F432",
			x"0000" when x"F433",
			x"0000" when x"F434",
			x"0000" when x"F435",
			x"0000" when x"F436",
			x"0000" when x"F437",
			x"0000" when x"F438",
			x"0000" when x"F439",
			x"0000" when x"F43A",
			x"0000" when x"F43B",
			x"0000" when x"F43C",
			x"0000" when x"F43D",
			x"0000" when x"F43E",
			x"0000" when x"F43F",
			x"0000" when x"F440",
			x"0000" when x"F441",
			x"0000" when x"F442",
			x"0000" when x"F443",
			x"0000" when x"F444",
			x"0000" when x"F445",
			x"0000" when x"F446",
			x"0000" when x"F447",
			x"0000" when x"F448",
			x"0000" when x"F449",
			x"0000" when x"F44A",
			x"0000" when x"F44B",
			x"0000" when x"F44C",
			x"0000" when x"F44D",
			x"0000" when x"F44E",
			x"0000" when x"F44F",
			x"0000" when x"F450",
			x"0000" when x"F451",
			x"0000" when x"F452",
			x"0000" when x"F453",
			x"0000" when x"F454",
			x"0000" when x"F455",
			x"0000" when x"F456",
			x"0000" when x"F457",
			x"0000" when x"F458",
			x"0000" when x"F459",
			x"0000" when x"F45A",
			x"0000" when x"F45B",
			x"0000" when x"F45C",
			x"0000" when x"F45D",
			x"0000" when x"F45E",
			x"0000" when x"F45F",
			x"0000" when x"F460",
			x"0000" when x"F461",
			x"0000" when x"F462",
			x"0000" when x"F463",
			x"0000" when x"F464",
			x"0000" when x"F465",
			x"0000" when x"F466",
			x"0000" when x"F467",
			x"0000" when x"F468",
			x"0000" when x"F469",
			x"0000" when x"F46A",
			x"0000" when x"F46B",
			x"0000" when x"F46C",
			x"0000" when x"F46D",
			x"0000" when x"F46E",
			x"0000" when x"F46F",
			x"0000" when x"F470",
			x"0000" when x"F471",
			x"0000" when x"F472",
			x"0000" when x"F473",
			x"0000" when x"F474",
			x"0000" when x"F475",
			x"0000" when x"F476",
			x"0000" when x"F477",
			x"0000" when x"F478",
			x"0000" when x"F479",
			x"0000" when x"F47A",
			x"0000" when x"F47B",
			x"0000" when x"F47C",
			x"0000" when x"F47D",
			x"0000" when x"F47E",
			x"0000" when x"F47F",
			x"0000" when x"F480",
			x"0000" when x"F481",
			x"0000" when x"F482",
			x"0000" when x"F483",
			x"0000" when x"F484",
			x"0000" when x"F485",
			x"0000" when x"F486",
			x"0000" when x"F487",
			x"0000" when x"F488",
			x"0000" when x"F489",
			x"0000" when x"F48A",
			x"0000" when x"F48B",
			x"0000" when x"F48C",
			x"0000" when x"F48D",
			x"0000" when x"F48E",
			x"0000" when x"F48F",
			x"0000" when x"F490",
			x"0000" when x"F491",
			x"0000" when x"F492",
			x"0000" when x"F493",
			x"0000" when x"F494",
			x"0000" when x"F495",
			x"0000" when x"F496",
			x"0000" when x"F497",
			x"0000" when x"F498",
			x"0000" when x"F499",
			x"0000" when x"F49A",
			x"0000" when x"F49B",
			x"0000" when x"F49C",
			x"0000" when x"F49D",
			x"0000" when x"F49E",
			x"0000" when x"F49F",
			x"0000" when x"F4A0",
			x"0000" when x"F4A1",
			x"0000" when x"F4A2",
			x"0000" when x"F4A3",
			x"0000" when x"F4A4",
			x"0000" when x"F4A5",
			x"0000" when x"F4A6",
			x"0000" when x"F4A7",
			x"0000" when x"F4A8",
			x"0000" when x"F4A9",
			x"0000" when x"F4AA",
			x"0000" when x"F4AB",
			x"0000" when x"F4AC",
			x"0000" when x"F4AD",
			x"0000" when x"F4AE",
			x"0000" when x"F4AF",
			x"0000" when x"F4B0",
			x"0000" when x"F4B1",
			x"0000" when x"F4B2",
			x"0000" when x"F4B3",
			x"0000" when x"F4B4",
			x"0000" when x"F4B5",
			x"0000" when x"F4B6",
			x"0000" when x"F4B7",
			x"0000" when x"F4B8",
			x"0000" when x"F4B9",
			x"0000" when x"F4BA",
			x"0000" when x"F4BB",
			x"0000" when x"F4BC",
			x"0000" when x"F4BD",
			x"0000" when x"F4BE",
			x"0000" when x"F4BF",
			x"0000" when x"F4C0",
			x"0000" when x"F4C1",
			x"0000" when x"F4C2",
			x"0000" when x"F4C3",
			x"0000" when x"F4C4",
			x"0000" when x"F4C5",
			x"0000" when x"F4C6",
			x"0000" when x"F4C7",
			x"0000" when x"F4C8",
			x"0000" when x"F4C9",
			x"0000" when x"F4CA",
			x"0000" when x"F4CB",
			x"0000" when x"F4CC",
			x"0000" when x"F4CD",
			x"0000" when x"F4CE",
			x"0000" when x"F4CF",
			x"0000" when x"F4D0",
			x"0000" when x"F4D1",
			x"0000" when x"F4D2",
			x"0000" when x"F4D3",
			x"0000" when x"F4D4",
			x"0000" when x"F4D5",
			x"0000" when x"F4D6",
			x"0000" when x"F4D7",
			x"0000" when x"F4D8",
			x"0000" when x"F4D9",
			x"0000" when x"F4DA",
			x"0000" when x"F4DB",
			x"0000" when x"F4DC",
			x"0000" when x"F4DD",
			x"0000" when x"F4DE",
			x"0000" when x"F4DF",
			x"0000" when x"F4E0",
			x"0000" when x"F4E1",
			x"0000" when x"F4E2",
			x"0000" when x"F4E3",
			x"0000" when x"F4E4",
			x"0000" when x"F4E5",
			x"0000" when x"F4E6",
			x"0000" when x"F4E7",
			x"0000" when x"F4E8",
			x"0000" when x"F4E9",
			x"0000" when x"F4EA",
			x"0000" when x"F4EB",
			x"0000" when x"F4EC",
			x"0000" when x"F4ED",
			x"0000" when x"F4EE",
			x"0000" when x"F4EF",
			x"0000" when x"F4F0",
			x"0000" when x"F4F1",
			x"0000" when x"F4F2",
			x"0000" when x"F4F3",
			x"0000" when x"F4F4",
			x"0000" when x"F4F5",
			x"0000" when x"F4F6",
			x"0000" when x"F4F7",
			x"0000" when x"F4F8",
			x"0000" when x"F4F9",
			x"0000" when x"F4FA",
			x"0000" when x"F4FB",
			x"0000" when x"F4FC",
			x"0000" when x"F4FD",
			x"0000" when x"F4FE",
			x"0000" when x"F4FF",
			x"0000" when x"F500",
			x"0000" when x"F501",
			x"0000" when x"F502",
			x"0000" when x"F503",
			x"0000" when x"F504",
			x"0000" when x"F505",
			x"0000" when x"F506",
			x"0000" when x"F507",
			x"0000" when x"F508",
			x"0000" when x"F509",
			x"0000" when x"F50A",
			x"0000" when x"F50B",
			x"0000" when x"F50C",
			x"0000" when x"F50D",
			x"0000" when x"F50E",
			x"0000" when x"F50F",
			x"0000" when x"F510",
			x"0000" when x"F511",
			x"0000" when x"F512",
			x"0000" when x"F513",
			x"0000" when x"F514",
			x"0000" when x"F515",
			x"0000" when x"F516",
			x"0000" when x"F517",
			x"0000" when x"F518",
			x"0000" when x"F519",
			x"0000" when x"F51A",
			x"0000" when x"F51B",
			x"0000" when x"F51C",
			x"0000" when x"F51D",
			x"0000" when x"F51E",
			x"0000" when x"F51F",
			x"0000" when x"F520",
			x"0000" when x"F521",
			x"0000" when x"F522",
			x"0000" when x"F523",
			x"0000" when x"F524",
			x"0000" when x"F525",
			x"0000" when x"F526",
			x"0000" when x"F527",
			x"0000" when x"F528",
			x"0000" when x"F529",
			x"0000" when x"F52A",
			x"0000" when x"F52B",
			x"0000" when x"F52C",
			x"0000" when x"F52D",
			x"0000" when x"F52E",
			x"0000" when x"F52F",
			x"0000" when x"F530",
			x"0000" when x"F531",
			x"0000" when x"F532",
			x"0000" when x"F533",
			x"0000" when x"F534",
			x"0000" when x"F535",
			x"0000" when x"F536",
			x"0000" when x"F537",
			x"0000" when x"F538",
			x"0000" when x"F539",
			x"0000" when x"F53A",
			x"0000" when x"F53B",
			x"0000" when x"F53C",
			x"0000" when x"F53D",
			x"0000" when x"F53E",
			x"0000" when x"F53F",
			x"0000" when x"F540",
			x"0000" when x"F541",
			x"0000" when x"F542",
			x"0000" when x"F543",
			x"0000" when x"F544",
			x"0000" when x"F545",
			x"0000" when x"F546",
			x"0000" when x"F547",
			x"0000" when x"F548",
			x"0000" when x"F549",
			x"0000" when x"F54A",
			x"0000" when x"F54B",
			x"0000" when x"F54C",
			x"0000" when x"F54D",
			x"0000" when x"F54E",
			x"0000" when x"F54F",
			x"0000" when x"F550",
			x"0000" when x"F551",
			x"0000" when x"F552",
			x"0000" when x"F553",
			x"0000" when x"F554",
			x"0000" when x"F555",
			x"0000" when x"F556",
			x"0000" when x"F557",
			x"0000" when x"F558",
			x"0000" when x"F559",
			x"0000" when x"F55A",
			x"0000" when x"F55B",
			x"0000" when x"F55C",
			x"0000" when x"F55D",
			x"0000" when x"F55E",
			x"0000" when x"F55F",
			x"0000" when x"F560",
			x"0000" when x"F561",
			x"0000" when x"F562",
			x"0000" when x"F563",
			x"0000" when x"F564",
			x"0000" when x"F565",
			x"0000" when x"F566",
			x"0000" when x"F567",
			x"0000" when x"F568",
			x"0000" when x"F569",
			x"0000" when x"F56A",
			x"0000" when x"F56B",
			x"0000" when x"F56C",
			x"0000" when x"F56D",
			x"0000" when x"F56E",
			x"0000" when x"F56F",
			x"0000" when x"F570",
			x"0000" when x"F571",
			x"0000" when x"F572",
			x"0000" when x"F573",
			x"0000" when x"F574",
			x"0000" when x"F575",
			x"0000" when x"F576",
			x"0000" when x"F577",
			x"0000" when x"F578",
			x"0000" when x"F579",
			x"0000" when x"F57A",
			x"0000" when x"F57B",
			x"0000" when x"F57C",
			x"0000" when x"F57D",
			x"0000" when x"F57E",
			x"0000" when x"F57F",
			x"0000" when x"F580",
			x"0000" when x"F581",
			x"0000" when x"F582",
			x"0000" when x"F583",
			x"0000" when x"F584",
			x"0000" when x"F585",
			x"0000" when x"F586",
			x"0000" when x"F587",
			x"0000" when x"F588",
			x"0000" when x"F589",
			x"0000" when x"F58A",
			x"0000" when x"F58B",
			x"0000" when x"F58C",
			x"0000" when x"F58D",
			x"0000" when x"F58E",
			x"0000" when x"F58F",
			x"0000" when x"F590",
			x"0000" when x"F591",
			x"0000" when x"F592",
			x"0000" when x"F593",
			x"0000" when x"F594",
			x"0000" when x"F595",
			x"0000" when x"F596",
			x"0000" when x"F597",
			x"0000" when x"F598",
			x"0000" when x"F599",
			x"0000" when x"F59A",
			x"0000" when x"F59B",
			x"0000" when x"F59C",
			x"0000" when x"F59D",
			x"0000" when x"F59E",
			x"0000" when x"F59F",
			x"0000" when x"F5A0",
			x"0000" when x"F5A1",
			x"0000" when x"F5A2",
			x"0000" when x"F5A3",
			x"0000" when x"F5A4",
			x"0000" when x"F5A5",
			x"0000" when x"F5A6",
			x"0000" when x"F5A7",
			x"0000" when x"F5A8",
			x"0000" when x"F5A9",
			x"0000" when x"F5AA",
			x"0000" when x"F5AB",
			x"0000" when x"F5AC",
			x"0000" when x"F5AD",
			x"0000" when x"F5AE",
			x"0000" when x"F5AF",
			x"0000" when x"F5B0",
			x"0000" when x"F5B1",
			x"0000" when x"F5B2",
			x"0000" when x"F5B3",
			x"0000" when x"F5B4",
			x"0000" when x"F5B5",
			x"0000" when x"F5B6",
			x"0000" when x"F5B7",
			x"0000" when x"F5B8",
			x"0000" when x"F5B9",
			x"0000" when x"F5BA",
			x"0000" when x"F5BB",
			x"0000" when x"F5BC",
			x"0000" when x"F5BD",
			x"0000" when x"F5BE",
			x"0000" when x"F5BF",
			x"0000" when x"F5C0",
			x"0000" when x"F5C1",
			x"0000" when x"F5C2",
			x"0000" when x"F5C3",
			x"0000" when x"F5C4",
			x"0000" when x"F5C5",
			x"0000" when x"F5C6",
			x"0000" when x"F5C7",
			x"0000" when x"F5C8",
			x"0000" when x"F5C9",
			x"0000" when x"F5CA",
			x"0000" when x"F5CB",
			x"0000" when x"F5CC",
			x"0000" when x"F5CD",
			x"0000" when x"F5CE",
			x"0000" when x"F5CF",
			x"0000" when x"F5D0",
			x"0000" when x"F5D1",
			x"0000" when x"F5D2",
			x"0000" when x"F5D3",
			x"0000" when x"F5D4",
			x"0000" when x"F5D5",
			x"0000" when x"F5D6",
			x"0000" when x"F5D7",
			x"0000" when x"F5D8",
			x"0000" when x"F5D9",
			x"0000" when x"F5DA",
			x"0000" when x"F5DB",
			x"0000" when x"F5DC",
			x"0000" when x"F5DD",
			x"0000" when x"F5DE",
			x"0000" when x"F5DF",
			x"0000" when x"F5E0",
			x"0000" when x"F5E1",
			x"0000" when x"F5E2",
			x"0000" when x"F5E3",
			x"0000" when x"F5E4",
			x"0000" when x"F5E5",
			x"0000" when x"F5E6",
			x"0000" when x"F5E7",
			x"0000" when x"F5E8",
			x"0000" when x"F5E9",
			x"0000" when x"F5EA",
			x"0000" when x"F5EB",
			x"0000" when x"F5EC",
			x"0000" when x"F5ED",
			x"0000" when x"F5EE",
			x"0000" when x"F5EF",
			x"0000" when x"F5F0",
			x"0000" when x"F5F1",
			x"0000" when x"F5F2",
			x"0000" when x"F5F3",
			x"0000" when x"F5F4",
			x"0000" when x"F5F5",
			x"0000" when x"F5F6",
			x"0000" when x"F5F7",
			x"0000" when x"F5F8",
			x"0000" when x"F5F9",
			x"0000" when x"F5FA",
			x"0000" when x"F5FB",
			x"0000" when x"F5FC",
			x"0000" when x"F5FD",
			x"0000" when x"F5FE",
			x"0000" when x"F5FF",
			x"0000" when x"F600",
			x"0000" when x"F601",
			x"0000" when x"F602",
			x"0000" when x"F603",
			x"0000" when x"F604",
			x"0000" when x"F605",
			x"0000" when x"F606",
			x"0000" when x"F607",
			x"0000" when x"F608",
			x"0000" when x"F609",
			x"0000" when x"F60A",
			x"0000" when x"F60B",
			x"0000" when x"F60C",
			x"0000" when x"F60D",
			x"0000" when x"F60E",
			x"0000" when x"F60F",
			x"0000" when x"F610",
			x"0000" when x"F611",
			x"0000" when x"F612",
			x"0000" when x"F613",
			x"0000" when x"F614",
			x"0000" when x"F615",
			x"0000" when x"F616",
			x"0000" when x"F617",
			x"0000" when x"F618",
			x"0000" when x"F619",
			x"0000" when x"F61A",
			x"0000" when x"F61B",
			x"0000" when x"F61C",
			x"0000" when x"F61D",
			x"0000" when x"F61E",
			x"0000" when x"F61F",
			x"0000" when x"F620",
			x"0000" when x"F621",
			x"0000" when x"F622",
			x"0000" when x"F623",
			x"0000" when x"F624",
			x"0000" when x"F625",
			x"0000" when x"F626",
			x"0000" when x"F627",
			x"0000" when x"F628",
			x"0000" when x"F629",
			x"0000" when x"F62A",
			x"0000" when x"F62B",
			x"0000" when x"F62C",
			x"0000" when x"F62D",
			x"0000" when x"F62E",
			x"0000" when x"F62F",
			x"0000" when x"F630",
			x"0000" when x"F631",
			x"0000" when x"F632",
			x"0000" when x"F633",
			x"0000" when x"F634",
			x"0000" when x"F635",
			x"0000" when x"F636",
			x"0000" when x"F637",
			x"0000" when x"F638",
			x"0000" when x"F639",
			x"0000" when x"F63A",
			x"0000" when x"F63B",
			x"0000" when x"F63C",
			x"0000" when x"F63D",
			x"0000" when x"F63E",
			x"0000" when x"F63F",
			x"0000" when x"F640",
			x"0000" when x"F641",
			x"0000" when x"F642",
			x"0000" when x"F643",
			x"0000" when x"F644",
			x"0000" when x"F645",
			x"0000" when x"F646",
			x"0000" when x"F647",
			x"0000" when x"F648",
			x"0000" when x"F649",
			x"0000" when x"F64A",
			x"0000" when x"F64B",
			x"0000" when x"F64C",
			x"0000" when x"F64D",
			x"0000" when x"F64E",
			x"0000" when x"F64F",
			x"0000" when x"F650",
			x"0000" when x"F651",
			x"0000" when x"F652",
			x"0000" when x"F653",
			x"0000" when x"F654",
			x"0000" when x"F655",
			x"0000" when x"F656",
			x"0000" when x"F657",
			x"0000" when x"F658",
			x"0000" when x"F659",
			x"0000" when x"F65A",
			x"0000" when x"F65B",
			x"0000" when x"F65C",
			x"0000" when x"F65D",
			x"0000" when x"F65E",
			x"0000" when x"F65F",
			x"0000" when x"F660",
			x"0000" when x"F661",
			x"0000" when x"F662",
			x"0000" when x"F663",
			x"0000" when x"F664",
			x"0000" when x"F665",
			x"0000" when x"F666",
			x"0000" when x"F667",
			x"0000" when x"F668",
			x"0000" when x"F669",
			x"0000" when x"F66A",
			x"0000" when x"F66B",
			x"0000" when x"F66C",
			x"0000" when x"F66D",
			x"0000" when x"F66E",
			x"0000" when x"F66F",
			x"0000" when x"F670",
			x"0000" when x"F671",
			x"0000" when x"F672",
			x"0000" when x"F673",
			x"0000" when x"F674",
			x"0000" when x"F675",
			x"0000" when x"F676",
			x"0000" when x"F677",
			x"0000" when x"F678",
			x"0000" when x"F679",
			x"0000" when x"F67A",
			x"0000" when x"F67B",
			x"0000" when x"F67C",
			x"0000" when x"F67D",
			x"0000" when x"F67E",
			x"0000" when x"F67F",
			x"0000" when x"F680",
			x"0000" when x"F681",
			x"0000" when x"F682",
			x"0000" when x"F683",
			x"0000" when x"F684",
			x"0000" when x"F685",
			x"0000" when x"F686",
			x"0000" when x"F687",
			x"0000" when x"F688",
			x"0000" when x"F689",
			x"0000" when x"F68A",
			x"0000" when x"F68B",
			x"0000" when x"F68C",
			x"0000" when x"F68D",
			x"0000" when x"F68E",
			x"0000" when x"F68F",
			x"0000" when x"F690",
			x"0000" when x"F691",
			x"0000" when x"F692",
			x"0000" when x"F693",
			x"0000" when x"F694",
			x"0000" when x"F695",
			x"0000" when x"F696",
			x"0000" when x"F697",
			x"0000" when x"F698",
			x"0000" when x"F699",
			x"0000" when x"F69A",
			x"0000" when x"F69B",
			x"0000" when x"F69C",
			x"0000" when x"F69D",
			x"0000" when x"F69E",
			x"0000" when x"F69F",
			x"0000" when x"F6A0",
			x"0000" when x"F6A1",
			x"0000" when x"F6A2",
			x"0000" when x"F6A3",
			x"0000" when x"F6A4",
			x"0000" when x"F6A5",
			x"0000" when x"F6A6",
			x"0000" when x"F6A7",
			x"0000" when x"F6A8",
			x"0000" when x"F6A9",
			x"0000" when x"F6AA",
			x"0000" when x"F6AB",
			x"0000" when x"F6AC",
			x"0000" when x"F6AD",
			x"0000" when x"F6AE",
			x"0000" when x"F6AF",
			x"0000" when x"F6B0",
			x"0000" when x"F6B1",
			x"0000" when x"F6B2",
			x"0000" when x"F6B3",
			x"0000" when x"F6B4",
			x"0000" when x"F6B5",
			x"0000" when x"F6B6",
			x"0000" when x"F6B7",
			x"0000" when x"F6B8",
			x"0000" when x"F6B9",
			x"0000" when x"F6BA",
			x"0000" when x"F6BB",
			x"0000" when x"F6BC",
			x"0000" when x"F6BD",
			x"0000" when x"F6BE",
			x"0000" when x"F6BF",
			x"0000" when x"F6C0",
			x"0000" when x"F6C1",
			x"0000" when x"F6C2",
			x"0000" when x"F6C3",
			x"0000" when x"F6C4",
			x"0000" when x"F6C5",
			x"0000" when x"F6C6",
			x"0000" when x"F6C7",
			x"0000" when x"F6C8",
			x"0000" when x"F6C9",
			x"0000" when x"F6CA",
			x"0000" when x"F6CB",
			x"0000" when x"F6CC",
			x"0000" when x"F6CD",
			x"0000" when x"F6CE",
			x"0000" when x"F6CF",
			x"0000" when x"F6D0",
			x"0000" when x"F6D1",
			x"0000" when x"F6D2",
			x"0000" when x"F6D3",
			x"0000" when x"F6D4",
			x"0000" when x"F6D5",
			x"0000" when x"F6D6",
			x"0000" when x"F6D7",
			x"0000" when x"F6D8",
			x"0000" when x"F6D9",
			x"0000" when x"F6DA",
			x"0000" when x"F6DB",
			x"0000" when x"F6DC",
			x"0000" when x"F6DD",
			x"0000" when x"F6DE",
			x"0000" when x"F6DF",
			x"0000" when x"F6E0",
			x"0000" when x"F6E1",
			x"0000" when x"F6E2",
			x"0000" when x"F6E3",
			x"0000" when x"F6E4",
			x"0000" when x"F6E5",
			x"0000" when x"F6E6",
			x"0000" when x"F6E7",
			x"0000" when x"F6E8",
			x"0000" when x"F6E9",
			x"0000" when x"F6EA",
			x"0000" when x"F6EB",
			x"0000" when x"F6EC",
			x"0000" when x"F6ED",
			x"0000" when x"F6EE",
			x"0000" when x"F6EF",
			x"0000" when x"F6F0",
			x"0000" when x"F6F1",
			x"0000" when x"F6F2",
			x"0000" when x"F6F3",
			x"0000" when x"F6F4",
			x"0000" when x"F6F5",
			x"0000" when x"F6F6",
			x"0000" when x"F6F7",
			x"0000" when x"F6F8",
			x"0000" when x"F6F9",
			x"0000" when x"F6FA",
			x"0000" when x"F6FB",
			x"0000" when x"F6FC",
			x"0000" when x"F6FD",
			x"0000" when x"F6FE",
			x"0000" when x"F6FF",
			x"0000" when x"F700",
			x"0000" when x"F701",
			x"0000" when x"F702",
			x"0000" when x"F703",
			x"0000" when x"F704",
			x"0000" when x"F705",
			x"0000" when x"F706",
			x"0000" when x"F707",
			x"0000" when x"F708",
			x"0000" when x"F709",
			x"0000" when x"F70A",
			x"0000" when x"F70B",
			x"0000" when x"F70C",
			x"0000" when x"F70D",
			x"0000" when x"F70E",
			x"0000" when x"F70F",
			x"0000" when x"F710",
			x"0000" when x"F711",
			x"0000" when x"F712",
			x"0000" when x"F713",
			x"0000" when x"F714",
			x"0000" when x"F715",
			x"0000" when x"F716",
			x"0000" when x"F717",
			x"0000" when x"F718",
			x"0000" when x"F719",
			x"0000" when x"F71A",
			x"0000" when x"F71B",
			x"0000" when x"F71C",
			x"0000" when x"F71D",
			x"0000" when x"F71E",
			x"0000" when x"F71F",
			x"0000" when x"F720",
			x"0000" when x"F721",
			x"0000" when x"F722",
			x"0000" when x"F723",
			x"0000" when x"F724",
			x"0000" when x"F725",
			x"0000" when x"F726",
			x"0000" when x"F727",
			x"0000" when x"F728",
			x"0000" when x"F729",
			x"0000" when x"F72A",
			x"0000" when x"F72B",
			x"0000" when x"F72C",
			x"0000" when x"F72D",
			x"0000" when x"F72E",
			x"0000" when x"F72F",
			x"0000" when x"F730",
			x"0000" when x"F731",
			x"0000" when x"F732",
			x"0000" when x"F733",
			x"0000" when x"F734",
			x"0000" when x"F735",
			x"0000" when x"F736",
			x"0000" when x"F737",
			x"0000" when x"F738",
			x"0000" when x"F739",
			x"0000" when x"F73A",
			x"0000" when x"F73B",
			x"0000" when x"F73C",
			x"0000" when x"F73D",
			x"0000" when x"F73E",
			x"0000" when x"F73F",
			x"0000" when x"F740",
			x"0000" when x"F741",
			x"0000" when x"F742",
			x"0000" when x"F743",
			x"0000" when x"F744",
			x"0000" when x"F745",
			x"0000" when x"F746",
			x"0000" when x"F747",
			x"0000" when x"F748",
			x"0000" when x"F749",
			x"0000" when x"F74A",
			x"0000" when x"F74B",
			x"0000" when x"F74C",
			x"0000" when x"F74D",
			x"0000" when x"F74E",
			x"0000" when x"F74F",
			x"0000" when x"F750",
			x"0000" when x"F751",
			x"0000" when x"F752",
			x"0000" when x"F753",
			x"0000" when x"F754",
			x"0000" when x"F755",
			x"0000" when x"F756",
			x"0000" when x"F757",
			x"0000" when x"F758",
			x"0000" when x"F759",
			x"0000" when x"F75A",
			x"0000" when x"F75B",
			x"0000" when x"F75C",
			x"0000" when x"F75D",
			x"0000" when x"F75E",
			x"0000" when x"F75F",
			x"0000" when x"F760",
			x"0000" when x"F761",
			x"0000" when x"F762",
			x"0000" when x"F763",
			x"0000" when x"F764",
			x"0000" when x"F765",
			x"0000" when x"F766",
			x"0000" when x"F767",
			x"0000" when x"F768",
			x"0000" when x"F769",
			x"0000" when x"F76A",
			x"0000" when x"F76B",
			x"0000" when x"F76C",
			x"0000" when x"F76D",
			x"0000" when x"F76E",
			x"0000" when x"F76F",
			x"0000" when x"F770",
			x"0000" when x"F771",
			x"0000" when x"F772",
			x"0000" when x"F773",
			x"0000" when x"F774",
			x"0000" when x"F775",
			x"0000" when x"F776",
			x"0000" when x"F777",
			x"0000" when x"F778",
			x"0000" when x"F779",
			x"0000" when x"F77A",
			x"0000" when x"F77B",
			x"0000" when x"F77C",
			x"0000" when x"F77D",
			x"0000" when x"F77E",
			x"0000" when x"F77F",
			x"0000" when x"F780",
			x"0000" when x"F781",
			x"0000" when x"F782",
			x"0000" when x"F783",
			x"0000" when x"F784",
			x"0000" when x"F785",
			x"0000" when x"F786",
			x"0000" when x"F787",
			x"0000" when x"F788",
			x"0000" when x"F789",
			x"0000" when x"F78A",
			x"0000" when x"F78B",
			x"0000" when x"F78C",
			x"0000" when x"F78D",
			x"0000" when x"F78E",
			x"0000" when x"F78F",
			x"0000" when x"F790",
			x"0000" when x"F791",
			x"0000" when x"F792",
			x"0000" when x"F793",
			x"0000" when x"F794",
			x"0000" when x"F795",
			x"0000" when x"F796",
			x"0000" when x"F797",
			x"0000" when x"F798",
			x"0000" when x"F799",
			x"0000" when x"F79A",
			x"0000" when x"F79B",
			x"0000" when x"F79C",
			x"0000" when x"F79D",
			x"0000" when x"F79E",
			x"0000" when x"F79F",
			x"0000" when x"F7A0",
			x"0000" when x"F7A1",
			x"0000" when x"F7A2",
			x"0000" when x"F7A3",
			x"0000" when x"F7A4",
			x"0000" when x"F7A5",
			x"0000" when x"F7A6",
			x"0000" when x"F7A7",
			x"0000" when x"F7A8",
			x"0000" when x"F7A9",
			x"0000" when x"F7AA",
			x"0000" when x"F7AB",
			x"0000" when x"F7AC",
			x"0000" when x"F7AD",
			x"0000" when x"F7AE",
			x"0000" when x"F7AF",
			x"0000" when x"F7B0",
			x"0000" when x"F7B1",
			x"0000" when x"F7B2",
			x"0000" when x"F7B3",
			x"0000" when x"F7B4",
			x"0000" when x"F7B5",
			x"0000" when x"F7B6",
			x"0000" when x"F7B7",
			x"0000" when x"F7B8",
			x"0000" when x"F7B9",
			x"0000" when x"F7BA",
			x"0000" when x"F7BB",
			x"0000" when x"F7BC",
			x"0000" when x"F7BD",
			x"0000" when x"F7BE",
			x"0000" when x"F7BF",
			x"0000" when x"F7C0",
			x"0000" when x"F7C1",
			x"0000" when x"F7C2",
			x"0000" when x"F7C3",
			x"0000" when x"F7C4",
			x"0000" when x"F7C5",
			x"0000" when x"F7C6",
			x"0000" when x"F7C7",
			x"0000" when x"F7C8",
			x"0000" when x"F7C9",
			x"0000" when x"F7CA",
			x"0000" when x"F7CB",
			x"0000" when x"F7CC",
			x"0000" when x"F7CD",
			x"0000" when x"F7CE",
			x"0000" when x"F7CF",
			x"0000" when x"F7D0",
			x"0000" when x"F7D1",
			x"0000" when x"F7D2",
			x"0000" when x"F7D3",
			x"0000" when x"F7D4",
			x"0000" when x"F7D5",
			x"0000" when x"F7D6",
			x"0000" when x"F7D7",
			x"0000" when x"F7D8",
			x"0000" when x"F7D9",
			x"0000" when x"F7DA",
			x"0000" when x"F7DB",
			x"0000" when x"F7DC",
			x"0000" when x"F7DD",
			x"0000" when x"F7DE",
			x"0000" when x"F7DF",
			x"0000" when x"F7E0",
			x"0000" when x"F7E1",
			x"0000" when x"F7E2",
			x"0000" when x"F7E3",
			x"0000" when x"F7E4",
			x"0000" when x"F7E5",
			x"0000" when x"F7E6",
			x"0000" when x"F7E7",
			x"0000" when x"F7E8",
			x"0000" when x"F7E9",
			x"0000" when x"F7EA",
			x"0000" when x"F7EB",
			x"0000" when x"F7EC",
			x"0000" when x"F7ED",
			x"0000" when x"F7EE",
			x"0000" when x"F7EF",
			x"0000" when x"F7F0",
			x"0000" when x"F7F1",
			x"0000" when x"F7F2",
			x"0000" when x"F7F3",
			x"0000" when x"F7F4",
			x"0000" when x"F7F5",
			x"0000" when x"F7F6",
			x"0000" when x"F7F7",
			x"0000" when x"F7F8",
			x"0000" when x"F7F9",
			x"0000" when x"F7FA",
			x"0000" when x"F7FB",
			x"0000" when x"F7FC",
			x"0000" when x"F7FD",
			x"0000" when x"F7FE",
			x"0000" when x"F7FF",
			x"0000" when x"F800",
			x"0000" when x"F801",
			x"0000" when x"F802",
			x"0000" when x"F803",
			x"0000" when x"F804",
			x"0000" when x"F805",
			x"0000" when x"F806",
			x"0000" when x"F807",
			x"0000" when x"F808",
			x"0000" when x"F809",
			x"0000" when x"F80A",
			x"0000" when x"F80B",
			x"0000" when x"F80C",
			x"0000" when x"F80D",
			x"0000" when x"F80E",
			x"0000" when x"F80F",
			x"0000" when x"F810",
			x"0000" when x"F811",
			x"0000" when x"F812",
			x"0000" when x"F813",
			x"0000" when x"F814",
			x"0000" when x"F815",
			x"0000" when x"F816",
			x"0000" when x"F817",
			x"0000" when x"F818",
			x"0000" when x"F819",
			x"0000" when x"F81A",
			x"0000" when x"F81B",
			x"0000" when x"F81C",
			x"0000" when x"F81D",
			x"0000" when x"F81E",
			x"0000" when x"F81F",
			x"0000" when x"F820",
			x"0000" when x"F821",
			x"0000" when x"F822",
			x"0000" when x"F823",
			x"0000" when x"F824",
			x"0000" when x"F825",
			x"0000" when x"F826",
			x"0000" when x"F827",
			x"0000" when x"F828",
			x"0000" when x"F829",
			x"0000" when x"F82A",
			x"0000" when x"F82B",
			x"0000" when x"F82C",
			x"0000" when x"F82D",
			x"0000" when x"F82E",
			x"0000" when x"F82F",
			x"0000" when x"F830",
			x"0000" when x"F831",
			x"0000" when x"F832",
			x"0000" when x"F833",
			x"0000" when x"F834",
			x"0000" when x"F835",
			x"0000" when x"F836",
			x"0000" when x"F837",
			x"0000" when x"F838",
			x"0000" when x"F839",
			x"0000" when x"F83A",
			x"0000" when x"F83B",
			x"0000" when x"F83C",
			x"0000" when x"F83D",
			x"0000" when x"F83E",
			x"0000" when x"F83F",
			x"0000" when x"F840",
			x"0000" when x"F841",
			x"0000" when x"F842",
			x"0000" when x"F843",
			x"0000" when x"F844",
			x"0000" when x"F845",
			x"0000" when x"F846",
			x"0000" when x"F847",
			x"0000" when x"F848",
			x"0000" when x"F849",
			x"0000" when x"F84A",
			x"0000" when x"F84B",
			x"0000" when x"F84C",
			x"0000" when x"F84D",
			x"0000" when x"F84E",
			x"0000" when x"F84F",
			x"0000" when x"F850",
			x"0000" when x"F851",
			x"0000" when x"F852",
			x"0000" when x"F853",
			x"0000" when x"F854",
			x"0000" when x"F855",
			x"0000" when x"F856",
			x"0000" when x"F857",
			x"0000" when x"F858",
			x"0000" when x"F859",
			x"0000" when x"F85A",
			x"0000" when x"F85B",
			x"0000" when x"F85C",
			x"0000" when x"F85D",
			x"0000" when x"F85E",
			x"0000" when x"F85F",
			x"0000" when x"F860",
			x"0000" when x"F861",
			x"0000" when x"F862",
			x"0000" when x"F863",
			x"0000" when x"F864",
			x"0000" when x"F865",
			x"0000" when x"F866",
			x"0000" when x"F867",
			x"0000" when x"F868",
			x"0000" when x"F869",
			x"0000" when x"F86A",
			x"0000" when x"F86B",
			x"0000" when x"F86C",
			x"0000" when x"F86D",
			x"0000" when x"F86E",
			x"0000" when x"F86F",
			x"0000" when x"F870",
			x"0000" when x"F871",
			x"0000" when x"F872",
			x"0000" when x"F873",
			x"0000" when x"F874",
			x"0000" when x"F875",
			x"0000" when x"F876",
			x"0000" when x"F877",
			x"0000" when x"F878",
			x"0000" when x"F879",
			x"0000" when x"F87A",
			x"0000" when x"F87B",
			x"0000" when x"F87C",
			x"0000" when x"F87D",
			x"0000" when x"F87E",
			x"0000" when x"F87F",
			x"0000" when x"F880",
			x"0000" when x"F881",
			x"0000" when x"F882",
			x"0000" when x"F883",
			x"0000" when x"F884",
			x"0000" when x"F885",
			x"0000" when x"F886",
			x"0000" when x"F887",
			x"0000" when x"F888",
			x"0000" when x"F889",
			x"0000" when x"F88A",
			x"0000" when x"F88B",
			x"0000" when x"F88C",
			x"0000" when x"F88D",
			x"0000" when x"F88E",
			x"0000" when x"F88F",
			x"0000" when x"F890",
			x"0000" when x"F891",
			x"0000" when x"F892",
			x"0000" when x"F893",
			x"0000" when x"F894",
			x"0000" when x"F895",
			x"0000" when x"F896",
			x"0000" when x"F897",
			x"0000" when x"F898",
			x"0000" when x"F899",
			x"0000" when x"F89A",
			x"0000" when x"F89B",
			x"0000" when x"F89C",
			x"0000" when x"F89D",
			x"0000" when x"F89E",
			x"0000" when x"F89F",
			x"0000" when x"F8A0",
			x"0000" when x"F8A1",
			x"0000" when x"F8A2",
			x"0000" when x"F8A3",
			x"0000" when x"F8A4",
			x"0000" when x"F8A5",
			x"0000" when x"F8A6",
			x"0000" when x"F8A7",
			x"0000" when x"F8A8",
			x"0000" when x"F8A9",
			x"0000" when x"F8AA",
			x"0000" when x"F8AB",
			x"0000" when x"F8AC",
			x"0000" when x"F8AD",
			x"0000" when x"F8AE",
			x"0000" when x"F8AF",
			x"0000" when x"F8B0",
			x"0000" when x"F8B1",
			x"0000" when x"F8B2",
			x"0000" when x"F8B3",
			x"0000" when x"F8B4",
			x"0000" when x"F8B5",
			x"0000" when x"F8B6",
			x"0000" when x"F8B7",
			x"0000" when x"F8B8",
			x"0000" when x"F8B9",
			x"0000" when x"F8BA",
			x"0000" when x"F8BB",
			x"0000" when x"F8BC",
			x"0000" when x"F8BD",
			x"0000" when x"F8BE",
			x"0000" when x"F8BF",
			x"0000" when x"F8C0",
			x"0000" when x"F8C1",
			x"0000" when x"F8C2",
			x"0000" when x"F8C3",
			x"0000" when x"F8C4",
			x"0000" when x"F8C5",
			x"0000" when x"F8C6",
			x"0000" when x"F8C7",
			x"0000" when x"F8C8",
			x"0000" when x"F8C9",
			x"0000" when x"F8CA",
			x"0000" when x"F8CB",
			x"0000" when x"F8CC",
			x"0000" when x"F8CD",
			x"0000" when x"F8CE",
			x"0000" when x"F8CF",
			x"0000" when x"F8D0",
			x"0000" when x"F8D1",
			x"0000" when x"F8D2",
			x"0000" when x"F8D3",
			x"0000" when x"F8D4",
			x"0000" when x"F8D5",
			x"0000" when x"F8D6",
			x"0000" when x"F8D7",
			x"0000" when x"F8D8",
			x"0000" when x"F8D9",
			x"0000" when x"F8DA",
			x"0000" when x"F8DB",
			x"0000" when x"F8DC",
			x"0000" when x"F8DD",
			x"0000" when x"F8DE",
			x"0000" when x"F8DF",
			x"0000" when x"F8E0",
			x"0000" when x"F8E1",
			x"0000" when x"F8E2",
			x"0000" when x"F8E3",
			x"0000" when x"F8E4",
			x"0000" when x"F8E5",
			x"0000" when x"F8E6",
			x"0000" when x"F8E7",
			x"0000" when x"F8E8",
			x"0000" when x"F8E9",
			x"0000" when x"F8EA",
			x"0000" when x"F8EB",
			x"0000" when x"F8EC",
			x"0000" when x"F8ED",
			x"0000" when x"F8EE",
			x"0000" when x"F8EF",
			x"0000" when x"F8F0",
			x"0000" when x"F8F1",
			x"0000" when x"F8F2",
			x"0000" when x"F8F3",
			x"0000" when x"F8F4",
			x"0000" when x"F8F5",
			x"0000" when x"F8F6",
			x"0000" when x"F8F7",
			x"0000" when x"F8F8",
			x"0000" when x"F8F9",
			x"0000" when x"F8FA",
			x"0000" when x"F8FB",
			x"0000" when x"F8FC",
			x"0000" when x"F8FD",
			x"0000" when x"F8FE",
			x"0000" when x"F8FF",
			x"0000" when x"F900",
			x"0000" when x"F901",
			x"0000" when x"F902",
			x"0000" when x"F903",
			x"0000" when x"F904",
			x"0000" when x"F905",
			x"0000" when x"F906",
			x"0000" when x"F907",
			x"0000" when x"F908",
			x"0000" when x"F909",
			x"0000" when x"F90A",
			x"0000" when x"F90B",
			x"0000" when x"F90C",
			x"0000" when x"F90D",
			x"0000" when x"F90E",
			x"0000" when x"F90F",
			x"0000" when x"F910",
			x"0000" when x"F911",
			x"0000" when x"F912",
			x"0000" when x"F913",
			x"0000" when x"F914",
			x"0000" when x"F915",
			x"0000" when x"F916",
			x"0000" when x"F917",
			x"0000" when x"F918",
			x"0000" when x"F919",
			x"0000" when x"F91A",
			x"0000" when x"F91B",
			x"0000" when x"F91C",
			x"0000" when x"F91D",
			x"0000" when x"F91E",
			x"0000" when x"F91F",
			x"0000" when x"F920",
			x"0000" when x"F921",
			x"0000" when x"F922",
			x"0000" when x"F923",
			x"0000" when x"F924",
			x"0000" when x"F925",
			x"0000" when x"F926",
			x"0000" when x"F927",
			x"0000" when x"F928",
			x"0000" when x"F929",
			x"0000" when x"F92A",
			x"0000" when x"F92B",
			x"0000" when x"F92C",
			x"0000" when x"F92D",
			x"0000" when x"F92E",
			x"0000" when x"F92F",
			x"0000" when x"F930",
			x"0000" when x"F931",
			x"0000" when x"F932",
			x"0000" when x"F933",
			x"0000" when x"F934",
			x"0000" when x"F935",
			x"0000" when x"F936",
			x"0000" when x"F937",
			x"0000" when x"F938",
			x"0000" when x"F939",
			x"0000" when x"F93A",
			x"0000" when x"F93B",
			x"0000" when x"F93C",
			x"0000" when x"F93D",
			x"0000" when x"F93E",
			x"0000" when x"F93F",
			x"0000" when x"F940",
			x"0000" when x"F941",
			x"0000" when x"F942",
			x"0000" when x"F943",
			x"0000" when x"F944",
			x"0000" when x"F945",
			x"0000" when x"F946",
			x"0000" when x"F947",
			x"0000" when x"F948",
			x"0000" when x"F949",
			x"0000" when x"F94A",
			x"0000" when x"F94B",
			x"0000" when x"F94C",
			x"0000" when x"F94D",
			x"0000" when x"F94E",
			x"0000" when x"F94F",
			x"0000" when x"F950",
			x"0000" when x"F951",
			x"0000" when x"F952",
			x"0000" when x"F953",
			x"0000" when x"F954",
			x"0000" when x"F955",
			x"0000" when x"F956",
			x"0000" when x"F957",
			x"0000" when x"F958",
			x"0000" when x"F959",
			x"0000" when x"F95A",
			x"0000" when x"F95B",
			x"0000" when x"F95C",
			x"0000" when x"F95D",
			x"0000" when x"F95E",
			x"0000" when x"F95F",
			x"0000" when x"F960",
			x"0000" when x"F961",
			x"0000" when x"F962",
			x"0000" when x"F963",
			x"0000" when x"F964",
			x"0000" when x"F965",
			x"0000" when x"F966",
			x"0000" when x"F967",
			x"0000" when x"F968",
			x"0000" when x"F969",
			x"0000" when x"F96A",
			x"0000" when x"F96B",
			x"0000" when x"F96C",
			x"0000" when x"F96D",
			x"0000" when x"F96E",
			x"0000" when x"F96F",
			x"0000" when x"F970",
			x"0000" when x"F971",
			x"0000" when x"F972",
			x"0000" when x"F973",
			x"0000" when x"F974",
			x"0000" when x"F975",
			x"0000" when x"F976",
			x"0000" when x"F977",
			x"0000" when x"F978",
			x"0000" when x"F979",
			x"0000" when x"F97A",
			x"0000" when x"F97B",
			x"0000" when x"F97C",
			x"0000" when x"F97D",
			x"0000" when x"F97E",
			x"0000" when x"F97F",
			x"0000" when x"F980",
			x"0000" when x"F981",
			x"0000" when x"F982",
			x"0000" when x"F983",
			x"0000" when x"F984",
			x"0000" when x"F985",
			x"0000" when x"F986",
			x"0000" when x"F987",
			x"0000" when x"F988",
			x"0000" when x"F989",
			x"0000" when x"F98A",
			x"0000" when x"F98B",
			x"0000" when x"F98C",
			x"0000" when x"F98D",
			x"0000" when x"F98E",
			x"0000" when x"F98F",
			x"0000" when x"F990",
			x"0000" when x"F991",
			x"0000" when x"F992",
			x"0000" when x"F993",
			x"0000" when x"F994",
			x"0000" when x"F995",
			x"0000" when x"F996",
			x"0000" when x"F997",
			x"0000" when x"F998",
			x"0000" when x"F999",
			x"0000" when x"F99A",
			x"0000" when x"F99B",
			x"0000" when x"F99C",
			x"0000" when x"F99D",
			x"0000" when x"F99E",
			x"0000" when x"F99F",
			x"0000" when x"F9A0",
			x"0000" when x"F9A1",
			x"0000" when x"F9A2",
			x"0000" when x"F9A3",
			x"0000" when x"F9A4",
			x"0000" when x"F9A5",
			x"0000" when x"F9A6",
			x"0000" when x"F9A7",
			x"0000" when x"F9A8",
			x"0000" when x"F9A9",
			x"0000" when x"F9AA",
			x"0000" when x"F9AB",
			x"0000" when x"F9AC",
			x"0000" when x"F9AD",
			x"0000" when x"F9AE",
			x"0000" when x"F9AF",
			x"0000" when x"F9B0",
			x"0000" when x"F9B1",
			x"0000" when x"F9B2",
			x"0000" when x"F9B3",
			x"0000" when x"F9B4",
			x"0000" when x"F9B5",
			x"0000" when x"F9B6",
			x"0000" when x"F9B7",
			x"0000" when x"F9B8",
			x"0000" when x"F9B9",
			x"0000" when x"F9BA",
			x"0000" when x"F9BB",
			x"0000" when x"F9BC",
			x"0000" when x"F9BD",
			x"0000" when x"F9BE",
			x"0000" when x"F9BF",
			x"0000" when x"F9C0",
			x"0000" when x"F9C1",
			x"0000" when x"F9C2",
			x"0000" when x"F9C3",
			x"0000" when x"F9C4",
			x"0000" when x"F9C5",
			x"0000" when x"F9C6",
			x"0000" when x"F9C7",
			x"0000" when x"F9C8",
			x"0000" when x"F9C9",
			x"0000" when x"F9CA",
			x"0000" when x"F9CB",
			x"0000" when x"F9CC",
			x"0000" when x"F9CD",
			x"0000" when x"F9CE",
			x"0000" when x"F9CF",
			x"0000" when x"F9D0",
			x"0000" when x"F9D1",
			x"0000" when x"F9D2",
			x"0000" when x"F9D3",
			x"0000" when x"F9D4",
			x"0000" when x"F9D5",
			x"0000" when x"F9D6",
			x"0000" when x"F9D7",
			x"0000" when x"F9D8",
			x"0000" when x"F9D9",
			x"0000" when x"F9DA",
			x"0000" when x"F9DB",
			x"0000" when x"F9DC",
			x"0000" when x"F9DD",
			x"0000" when x"F9DE",
			x"0000" when x"F9DF",
			x"0000" when x"F9E0",
			x"0000" when x"F9E1",
			x"0000" when x"F9E2",
			x"0000" when x"F9E3",
			x"0000" when x"F9E4",
			x"0000" when x"F9E5",
			x"0000" when x"F9E6",
			x"0000" when x"F9E7",
			x"0000" when x"F9E8",
			x"0000" when x"F9E9",
			x"0000" when x"F9EA",
			x"0000" when x"F9EB",
			x"0000" when x"F9EC",
			x"0000" when x"F9ED",
			x"0000" when x"F9EE",
			x"0000" when x"F9EF",
			x"0000" when x"F9F0",
			x"0000" when x"F9F1",
			x"0000" when x"F9F2",
			x"0000" when x"F9F3",
			x"0000" when x"F9F4",
			x"0000" when x"F9F5",
			x"0000" when x"F9F6",
			x"0000" when x"F9F7",
			x"0000" when x"F9F8",
			x"0000" when x"F9F9",
			x"0000" when x"F9FA",
			x"0000" when x"F9FB",
			x"0000" when x"F9FC",
			x"0000" when x"F9FD",
			x"0000" when x"F9FE",
			x"0000" when x"F9FF",
			x"0000" when x"FA00",
			x"0000" when x"FA01",
			x"0000" when x"FA02",
			x"0000" when x"FA03",
			x"0000" when x"FA04",
			x"0000" when x"FA05",
			x"0000" when x"FA06",
			x"0000" when x"FA07",
			x"0000" when x"FA08",
			x"0000" when x"FA09",
			x"0000" when x"FA0A",
			x"0000" when x"FA0B",
			x"0000" when x"FA0C",
			x"0000" when x"FA0D",
			x"0000" when x"FA0E",
			x"0000" when x"FA0F",
			x"0000" when x"FA10",
			x"0000" when x"FA11",
			x"0000" when x"FA12",
			x"0000" when x"FA13",
			x"0000" when x"FA14",
			x"0000" when x"FA15",
			x"0000" when x"FA16",
			x"0000" when x"FA17",
			x"0000" when x"FA18",
			x"0000" when x"FA19",
			x"0000" when x"FA1A",
			x"0000" when x"FA1B",
			x"0000" when x"FA1C",
			x"0000" when x"FA1D",
			x"0000" when x"FA1E",
			x"0000" when x"FA1F",
			x"0000" when x"FA20",
			x"0000" when x"FA21",
			x"0000" when x"FA22",
			x"0000" when x"FA23",
			x"0000" when x"FA24",
			x"0000" when x"FA25",
			x"0000" when x"FA26",
			x"0000" when x"FA27",
			x"0000" when x"FA28",
			x"0000" when x"FA29",
			x"0000" when x"FA2A",
			x"0000" when x"FA2B",
			x"0000" when x"FA2C",
			x"0000" when x"FA2D",
			x"0000" when x"FA2E",
			x"0000" when x"FA2F",
			x"0000" when x"FA30",
			x"0000" when x"FA31",
			x"0000" when x"FA32",
			x"0000" when x"FA33",
			x"0000" when x"FA34",
			x"0000" when x"FA35",
			x"0000" when x"FA36",
			x"0000" when x"FA37",
			x"0000" when x"FA38",
			x"0000" when x"FA39",
			x"0000" when x"FA3A",
			x"0000" when x"FA3B",
			x"0000" when x"FA3C",
			x"0000" when x"FA3D",
			x"0000" when x"FA3E",
			x"0000" when x"FA3F",
			x"0000" when x"FA40",
			x"0000" when x"FA41",
			x"0000" when x"FA42",
			x"0000" when x"FA43",
			x"0000" when x"FA44",
			x"0000" when x"FA45",
			x"0000" when x"FA46",
			x"0000" when x"FA47",
			x"0000" when x"FA48",
			x"0000" when x"FA49",
			x"0000" when x"FA4A",
			x"0000" when x"FA4B",
			x"0000" when x"FA4C",
			x"0000" when x"FA4D",
			x"0000" when x"FA4E",
			x"0000" when x"FA4F",
			x"0000" when x"FA50",
			x"0000" when x"FA51",
			x"0000" when x"FA52",
			x"0000" when x"FA53",
			x"0000" when x"FA54",
			x"0000" when x"FA55",
			x"0000" when x"FA56",
			x"0000" when x"FA57",
			x"0000" when x"FA58",
			x"0000" when x"FA59",
			x"0000" when x"FA5A",
			x"0000" when x"FA5B",
			x"0000" when x"FA5C",
			x"0000" when x"FA5D",
			x"0000" when x"FA5E",
			x"0000" when x"FA5F",
			x"0000" when x"FA60",
			x"0000" when x"FA61",
			x"0000" when x"FA62",
			x"0000" when x"FA63",
			x"0000" when x"FA64",
			x"0000" when x"FA65",
			x"0000" when x"FA66",
			x"0000" when x"FA67",
			x"0000" when x"FA68",
			x"0000" when x"FA69",
			x"0000" when x"FA6A",
			x"0000" when x"FA6B",
			x"0000" when x"FA6C",
			x"0000" when x"FA6D",
			x"0000" when x"FA6E",
			x"0000" when x"FA6F",
			x"0000" when x"FA70",
			x"0000" when x"FA71",
			x"0000" when x"FA72",
			x"0000" when x"FA73",
			x"0000" when x"FA74",
			x"0000" when x"FA75",
			x"0000" when x"FA76",
			x"0000" when x"FA77",
			x"0000" when x"FA78",
			x"0000" when x"FA79",
			x"0000" when x"FA7A",
			x"0000" when x"FA7B",
			x"0000" when x"FA7C",
			x"0000" when x"FA7D",
			x"0000" when x"FA7E",
			x"0000" when x"FA7F",
			x"0000" when x"FA80",
			x"0000" when x"FA81",
			x"0000" when x"FA82",
			x"0000" when x"FA83",
			x"0000" when x"FA84",
			x"0000" when x"FA85",
			x"0000" when x"FA86",
			x"0000" when x"FA87",
			x"0000" when x"FA88",
			x"0000" when x"FA89",
			x"0000" when x"FA8A",
			x"0000" when x"FA8B",
			x"0000" when x"FA8C",
			x"0000" when x"FA8D",
			x"0000" when x"FA8E",
			x"0000" when x"FA8F",
			x"0000" when x"FA90",
			x"0000" when x"FA91",
			x"0000" when x"FA92",
			x"0000" when x"FA93",
			x"0000" when x"FA94",
			x"0000" when x"FA95",
			x"0000" when x"FA96",
			x"0000" when x"FA97",
			x"0000" when x"FA98",
			x"0000" when x"FA99",
			x"0000" when x"FA9A",
			x"0000" when x"FA9B",
			x"0000" when x"FA9C",
			x"0000" when x"FA9D",
			x"0000" when x"FA9E",
			x"0000" when x"FA9F",
			x"0000" when x"FAA0",
			x"0000" when x"FAA1",
			x"0000" when x"FAA2",
			x"0000" when x"FAA3",
			x"0000" when x"FAA4",
			x"0000" when x"FAA5",
			x"0000" when x"FAA6",
			x"0000" when x"FAA7",
			x"0000" when x"FAA8",
			x"0000" when x"FAA9",
			x"0000" when x"FAAA",
			x"0000" when x"FAAB",
			x"0000" when x"FAAC",
			x"0000" when x"FAAD",
			x"0000" when x"FAAE",
			x"0000" when x"FAAF",
			x"0000" when x"FAB0",
			x"0000" when x"FAB1",
			x"0000" when x"FAB2",
			x"0000" when x"FAB3",
			x"0000" when x"FAB4",
			x"0000" when x"FAB5",
			x"0000" when x"FAB6",
			x"0000" when x"FAB7",
			x"0000" when x"FAB8",
			x"0000" when x"FAB9",
			x"0000" when x"FABA",
			x"0000" when x"FABB",
			x"0000" when x"FABC",
			x"0000" when x"FABD",
			x"0000" when x"FABE",
			x"0000" when x"FABF",
			x"0000" when x"FAC0",
			x"0000" when x"FAC1",
			x"0000" when x"FAC2",
			x"0000" when x"FAC3",
			x"0000" when x"FAC4",
			x"0000" when x"FAC5",
			x"0000" when x"FAC6",
			x"0000" when x"FAC7",
			x"0000" when x"FAC8",
			x"0000" when x"FAC9",
			x"0000" when x"FACA",
			x"0000" when x"FACB",
			x"0000" when x"FACC",
			x"0000" when x"FACD",
			x"0000" when x"FACE",
			x"0000" when x"FACF",
			x"0000" when x"FAD0",
			x"0000" when x"FAD1",
			x"0000" when x"FAD2",
			x"0000" when x"FAD3",
			x"0000" when x"FAD4",
			x"0000" when x"FAD5",
			x"0000" when x"FAD6",
			x"0000" when x"FAD7",
			x"0000" when x"FAD8",
			x"0000" when x"FAD9",
			x"0000" when x"FADA",
			x"0000" when x"FADB",
			x"0000" when x"FADC",
			x"0000" when x"FADD",
			x"0000" when x"FADE",
			x"0000" when x"FADF",
			x"0000" when x"FAE0",
			x"0000" when x"FAE1",
			x"0000" when x"FAE2",
			x"0000" when x"FAE3",
			x"0000" when x"FAE4",
			x"0000" when x"FAE5",
			x"0000" when x"FAE6",
			x"0000" when x"FAE7",
			x"0000" when x"FAE8",
			x"0000" when x"FAE9",
			x"0000" when x"FAEA",
			x"0000" when x"FAEB",
			x"0000" when x"FAEC",
			x"0000" when x"FAED",
			x"0000" when x"FAEE",
			x"0000" when x"FAEF",
			x"0000" when x"FAF0",
			x"0000" when x"FAF1",
			x"0000" when x"FAF2",
			x"0000" when x"FAF3",
			x"0000" when x"FAF4",
			x"0000" when x"FAF5",
			x"0000" when x"FAF6",
			x"0000" when x"FAF7",
			x"0000" when x"FAF8",
			x"0000" when x"FAF9",
			x"0000" when x"FAFA",
			x"0000" when x"FAFB",
			x"0000" when x"FAFC",
			x"0000" when x"FAFD",
			x"0000" when x"FAFE",
			x"0000" when x"FAFF",
			x"0000" when x"FB00",
			x"0000" when x"FB01",
			x"0000" when x"FB02",
			x"0000" when x"FB03",
			x"0000" when x"FB04",
			x"0000" when x"FB05",
			x"0000" when x"FB06",
			x"0000" when x"FB07",
			x"0000" when x"FB08",
			x"0000" when x"FB09",
			x"0000" when x"FB0A",
			x"0000" when x"FB0B",
			x"0000" when x"FB0C",
			x"0000" when x"FB0D",
			x"0000" when x"FB0E",
			x"0000" when x"FB0F",
			x"0000" when x"FB10",
			x"0000" when x"FB11",
			x"0000" when x"FB12",
			x"0000" when x"FB13",
			x"0000" when x"FB14",
			x"0000" when x"FB15",
			x"0000" when x"FB16",
			x"0000" when x"FB17",
			x"0000" when x"FB18",
			x"0000" when x"FB19",
			x"0000" when x"FB1A",
			x"0000" when x"FB1B",
			x"0000" when x"FB1C",
			x"0000" when x"FB1D",
			x"0000" when x"FB1E",
			x"0000" when x"FB1F",
			x"0000" when x"FB20",
			x"0000" when x"FB21",
			x"0000" when x"FB22",
			x"0000" when x"FB23",
			x"0000" when x"FB24",
			x"0000" when x"FB25",
			x"0000" when x"FB26",
			x"0000" when x"FB27",
			x"0000" when x"FB28",
			x"0000" when x"FB29",
			x"0000" when x"FB2A",
			x"0000" when x"FB2B",
			x"0000" when x"FB2C",
			x"0000" when x"FB2D",
			x"0000" when x"FB2E",
			x"0000" when x"FB2F",
			x"0000" when x"FB30",
			x"0000" when x"FB31",
			x"0000" when x"FB32",
			x"0000" when x"FB33",
			x"0000" when x"FB34",
			x"0000" when x"FB35",
			x"0000" when x"FB36",
			x"0000" when x"FB37",
			x"0000" when x"FB38",
			x"0000" when x"FB39",
			x"0000" when x"FB3A",
			x"0000" when x"FB3B",
			x"0000" when x"FB3C",
			x"0000" when x"FB3D",
			x"0000" when x"FB3E",
			x"0000" when x"FB3F",
			x"0000" when x"FB40",
			x"0000" when x"FB41",
			x"0000" when x"FB42",
			x"0000" when x"FB43",
			x"0000" when x"FB44",
			x"0000" when x"FB45",
			x"0000" when x"FB46",
			x"0000" when x"FB47",
			x"0000" when x"FB48",
			x"0000" when x"FB49",
			x"0000" when x"FB4A",
			x"0000" when x"FB4B",
			x"0000" when x"FB4C",
			x"0000" when x"FB4D",
			x"0000" when x"FB4E",
			x"0000" when x"FB4F",
			x"0000" when x"FB50",
			x"0000" when x"FB51",
			x"0000" when x"FB52",
			x"0000" when x"FB53",
			x"0000" when x"FB54",
			x"0000" when x"FB55",
			x"0000" when x"FB56",
			x"0000" when x"FB57",
			x"0000" when x"FB58",
			x"0000" when x"FB59",
			x"0000" when x"FB5A",
			x"0000" when x"FB5B",
			x"0000" when x"FB5C",
			x"0000" when x"FB5D",
			x"0000" when x"FB5E",
			x"0000" when x"FB5F",
			x"0000" when x"FB60",
			x"0000" when x"FB61",
			x"0000" when x"FB62",
			x"0000" when x"FB63",
			x"0000" when x"FB64",
			x"0000" when x"FB65",
			x"0000" when x"FB66",
			x"0000" when x"FB67",
			x"0000" when x"FB68",
			x"0000" when x"FB69",
			x"0000" when x"FB6A",
			x"0000" when x"FB6B",
			x"0000" when x"FB6C",
			x"0000" when x"FB6D",
			x"0000" when x"FB6E",
			x"0000" when x"FB6F",
			x"0000" when x"FB70",
			x"0000" when x"FB71",
			x"0000" when x"FB72",
			x"0000" when x"FB73",
			x"0000" when x"FB74",
			x"0000" when x"FB75",
			x"0000" when x"FB76",
			x"0000" when x"FB77",
			x"0000" when x"FB78",
			x"0000" when x"FB79",
			x"0000" when x"FB7A",
			x"0000" when x"FB7B",
			x"0000" when x"FB7C",
			x"0000" when x"FB7D",
			x"0000" when x"FB7E",
			x"0000" when x"FB7F",
			x"0000" when x"FB80",
			x"0000" when x"FB81",
			x"0000" when x"FB82",
			x"0000" when x"FB83",
			x"0000" when x"FB84",
			x"0000" when x"FB85",
			x"0000" when x"FB86",
			x"0000" when x"FB87",
			x"0000" when x"FB88",
			x"0000" when x"FB89",
			x"0000" when x"FB8A",
			x"0000" when x"FB8B",
			x"0000" when x"FB8C",
			x"0000" when x"FB8D",
			x"0000" when x"FB8E",
			x"0000" when x"FB8F",
			x"0000" when x"FB90",
			x"0000" when x"FB91",
			x"0000" when x"FB92",
			x"0000" when x"FB93",
			x"0000" when x"FB94",
			x"0000" when x"FB95",
			x"0000" when x"FB96",
			x"0000" when x"FB97",
			x"0000" when x"FB98",
			x"0000" when x"FB99",
			x"0000" when x"FB9A",
			x"0000" when x"FB9B",
			x"0000" when x"FB9C",
			x"0000" when x"FB9D",
			x"0000" when x"FB9E",
			x"0000" when x"FB9F",
			x"0000" when x"FBA0",
			x"0000" when x"FBA1",
			x"0000" when x"FBA2",
			x"0000" when x"FBA3",
			x"0000" when x"FBA4",
			x"0000" when x"FBA5",
			x"0000" when x"FBA6",
			x"0000" when x"FBA7",
			x"0000" when x"FBA8",
			x"0000" when x"FBA9",
			x"0000" when x"FBAA",
			x"0000" when x"FBAB",
			x"0000" when x"FBAC",
			x"0000" when x"FBAD",
			x"0000" when x"FBAE",
			x"0000" when x"FBAF",
			x"0000" when x"FBB0",
			x"0000" when x"FBB1",
			x"0000" when x"FBB2",
			x"0000" when x"FBB3",
			x"0000" when x"FBB4",
			x"0000" when x"FBB5",
			x"0000" when x"FBB6",
			x"0000" when x"FBB7",
			x"0000" when x"FBB8",
			x"0000" when x"FBB9",
			x"0000" when x"FBBA",
			x"0000" when x"FBBB",
			x"0000" when x"FBBC",
			x"0000" when x"FBBD",
			x"0000" when x"FBBE",
			x"0000" when x"FBBF",
			x"0000" when x"FBC0",
			x"0000" when x"FBC1",
			x"0000" when x"FBC2",
			x"0000" when x"FBC3",
			x"0000" when x"FBC4",
			x"0000" when x"FBC5",
			x"0000" when x"FBC6",
			x"0000" when x"FBC7",
			x"0000" when x"FBC8",
			x"0000" when x"FBC9",
			x"0000" when x"FBCA",
			x"0000" when x"FBCB",
			x"0000" when x"FBCC",
			x"0000" when x"FBCD",
			x"0000" when x"FBCE",
			x"0000" when x"FBCF",
			x"0000" when x"FBD0",
			x"0000" when x"FBD1",
			x"0000" when x"FBD2",
			x"0000" when x"FBD3",
			x"0000" when x"FBD4",
			x"0000" when x"FBD5",
			x"0000" when x"FBD6",
			x"0000" when x"FBD7",
			x"0000" when x"FBD8",
			x"0000" when x"FBD9",
			x"0000" when x"FBDA",
			x"0000" when x"FBDB",
			x"0000" when x"FBDC",
			x"0000" when x"FBDD",
			x"0000" when x"FBDE",
			x"0000" when x"FBDF",
			x"0000" when x"FBE0",
			x"0000" when x"FBE1",
			x"0000" when x"FBE2",
			x"0000" when x"FBE3",
			x"0000" when x"FBE4",
			x"0000" when x"FBE5",
			x"0000" when x"FBE6",
			x"0000" when x"FBE7",
			x"0000" when x"FBE8",
			x"0000" when x"FBE9",
			x"0000" when x"FBEA",
			x"0000" when x"FBEB",
			x"0000" when x"FBEC",
			x"0000" when x"FBED",
			x"0000" when x"FBEE",
			x"0000" when x"FBEF",
			x"0000" when x"FBF0",
			x"0000" when x"FBF1",
			x"0000" when x"FBF2",
			x"0000" when x"FBF3",
			x"0000" when x"FBF4",
			x"0000" when x"FBF5",
			x"0000" when x"FBF6",
			x"0000" when x"FBF7",
			x"0000" when x"FBF8",
			x"0000" when x"FBF9",
			x"0000" when x"FBFA",
			x"0000" when x"FBFB",
			x"0000" when x"FBFC",
			x"0000" when x"FBFD",
			x"0000" when x"FBFE",
			x"0000" when x"FBFF",
			x"0000" when x"FC00",
			x"0000" when x"FC01",
			x"0000" when x"FC02",
			x"0000" when x"FC03",
			x"0000" when x"FC04",
			x"0000" when x"FC05",
			x"0000" when x"FC06",
			x"0000" when x"FC07",
			x"0000" when x"FC08",
			x"0000" when x"FC09",
			x"0000" when x"FC0A",
			x"0000" when x"FC0B",
			x"0000" when x"FC0C",
			x"0000" when x"FC0D",
			x"0000" when x"FC0E",
			x"0000" when x"FC0F",
			x"0000" when x"FC10",
			x"0000" when x"FC11",
			x"0000" when x"FC12",
			x"0000" when x"FC13",
			x"0000" when x"FC14",
			x"0000" when x"FC15",
			x"0000" when x"FC16",
			x"0000" when x"FC17",
			x"0000" when x"FC18",
			x"0000" when x"FC19",
			x"0000" when x"FC1A",
			x"0000" when x"FC1B",
			x"0000" when x"FC1C",
			x"0000" when x"FC1D",
			x"0000" when x"FC1E",
			x"0000" when x"FC1F",
			x"0000" when x"FC20",
			x"0000" when x"FC21",
			x"0000" when x"FC22",
			x"0000" when x"FC23",
			x"0000" when x"FC24",
			x"0000" when x"FC25",
			x"0000" when x"FC26",
			x"0000" when x"FC27",
			x"0000" when x"FC28",
			x"0000" when x"FC29",
			x"0000" when x"FC2A",
			x"0000" when x"FC2B",
			x"0000" when x"FC2C",
			x"0000" when x"FC2D",
			x"0000" when x"FC2E",
			x"0000" when x"FC2F",
			x"0000" when x"FC30",
			x"0000" when x"FC31",
			x"0000" when x"FC32",
			x"0000" when x"FC33",
			x"0000" when x"FC34",
			x"0000" when x"FC35",
			x"0000" when x"FC36",
			x"0000" when x"FC37",
			x"0000" when x"FC38",
			x"0000" when x"FC39",
			x"0000" when x"FC3A",
			x"0000" when x"FC3B",
			x"0000" when x"FC3C",
			x"0000" when x"FC3D",
			x"0000" when x"FC3E",
			x"0000" when x"FC3F",
			x"0000" when x"FC40",
			x"0000" when x"FC41",
			x"0000" when x"FC42",
			x"0000" when x"FC43",
			x"0000" when x"FC44",
			x"0000" when x"FC45",
			x"0000" when x"FC46",
			x"0000" when x"FC47",
			x"0000" when x"FC48",
			x"0000" when x"FC49",
			x"0000" when x"FC4A",
			x"0000" when x"FC4B",
			x"0000" when x"FC4C",
			x"0000" when x"FC4D",
			x"0000" when x"FC4E",
			x"0000" when x"FC4F",
			x"0000" when x"FC50",
			x"0000" when x"FC51",
			x"0000" when x"FC52",
			x"0000" when x"FC53",
			x"0000" when x"FC54",
			x"0000" when x"FC55",
			x"0000" when x"FC56",
			x"0000" when x"FC57",
			x"0000" when x"FC58",
			x"0000" when x"FC59",
			x"0000" when x"FC5A",
			x"0000" when x"FC5B",
			x"0000" when x"FC5C",
			x"0000" when x"FC5D",
			x"0000" when x"FC5E",
			x"0000" when x"FC5F",
			x"0000" when x"FC60",
			x"0000" when x"FC61",
			x"0000" when x"FC62",
			x"0000" when x"FC63",
			x"0000" when x"FC64",
			x"0000" when x"FC65",
			x"0000" when x"FC66",
			x"0000" when x"FC67",
			x"0000" when x"FC68",
			x"0000" when x"FC69",
			x"0000" when x"FC6A",
			x"0000" when x"FC6B",
			x"0000" when x"FC6C",
			x"0000" when x"FC6D",
			x"0000" when x"FC6E",
			x"0000" when x"FC6F",
			x"0000" when x"FC70",
			x"0000" when x"FC71",
			x"0000" when x"FC72",
			x"0000" when x"FC73",
			x"0000" when x"FC74",
			x"0000" when x"FC75",
			x"0000" when x"FC76",
			x"0000" when x"FC77",
			x"0000" when x"FC78",
			x"0000" when x"FC79",
			x"0000" when x"FC7A",
			x"0000" when x"FC7B",
			x"0000" when x"FC7C",
			x"0000" when x"FC7D",
			x"0000" when x"FC7E",
			x"0000" when x"FC7F",
			x"0000" when x"FC80",
			x"0000" when x"FC81",
			x"0000" when x"FC82",
			x"0000" when x"FC83",
			x"0000" when x"FC84",
			x"0000" when x"FC85",
			x"0000" when x"FC86",
			x"0000" when x"FC87",
			x"0000" when x"FC88",
			x"0000" when x"FC89",
			x"0000" when x"FC8A",
			x"0000" when x"FC8B",
			x"0000" when x"FC8C",
			x"0000" when x"FC8D",
			x"0000" when x"FC8E",
			x"0000" when x"FC8F",
			x"0000" when x"FC90",
			x"0000" when x"FC91",
			x"0000" when x"FC92",
			x"0000" when x"FC93",
			x"0000" when x"FC94",
			x"0000" when x"FC95",
			x"0000" when x"FC96",
			x"0000" when x"FC97",
			x"0000" when x"FC98",
			x"0000" when x"FC99",
			x"0000" when x"FC9A",
			x"0000" when x"FC9B",
			x"0000" when x"FC9C",
			x"0000" when x"FC9D",
			x"0000" when x"FC9E",
			x"0000" when x"FC9F",
			x"0000" when x"FCA0",
			x"0000" when x"FCA1",
			x"0000" when x"FCA2",
			x"0000" when x"FCA3",
			x"0000" when x"FCA4",
			x"0000" when x"FCA5",
			x"0000" when x"FCA6",
			x"0000" when x"FCA7",
			x"0000" when x"FCA8",
			x"0000" when x"FCA9",
			x"0000" when x"FCAA",
			x"0000" when x"FCAB",
			x"0000" when x"FCAC",
			x"0000" when x"FCAD",
			x"0000" when x"FCAE",
			x"0000" when x"FCAF",
			x"0000" when x"FCB0",
			x"0000" when x"FCB1",
			x"0000" when x"FCB2",
			x"0000" when x"FCB3",
			x"0000" when x"FCB4",
			x"0000" when x"FCB5",
			x"0000" when x"FCB6",
			x"0000" when x"FCB7",
			x"0000" when x"FCB8",
			x"0000" when x"FCB9",
			x"0000" when x"FCBA",
			x"0000" when x"FCBB",
			x"0000" when x"FCBC",
			x"0000" when x"FCBD",
			x"0000" when x"FCBE",
			x"0000" when x"FCBF",
			x"0000" when x"FCC0",
			x"0000" when x"FCC1",
			x"0000" when x"FCC2",
			x"0000" when x"FCC3",
			x"0000" when x"FCC4",
			x"0000" when x"FCC5",
			x"0000" when x"FCC6",
			x"0000" when x"FCC7",
			x"0000" when x"FCC8",
			x"0000" when x"FCC9",
			x"0000" when x"FCCA",
			x"0000" when x"FCCB",
			x"0000" when x"FCCC",
			x"0000" when x"FCCD",
			x"0000" when x"FCCE",
			x"0000" when x"FCCF",
			x"0000" when x"FCD0",
			x"0000" when x"FCD1",
			x"0000" when x"FCD2",
			x"0000" when x"FCD3",
			x"0000" when x"FCD4",
			x"0000" when x"FCD5",
			x"0000" when x"FCD6",
			x"0000" when x"FCD7",
			x"0000" when x"FCD8",
			x"0000" when x"FCD9",
			x"0000" when x"FCDA",
			x"0000" when x"FCDB",
			x"0000" when x"FCDC",
			x"0000" when x"FCDD",
			x"0000" when x"FCDE",
			x"0000" when x"FCDF",
			x"0000" when x"FCE0",
			x"0000" when x"FCE1",
			x"0000" when x"FCE2",
			x"0000" when x"FCE3",
			x"0000" when x"FCE4",
			x"0000" when x"FCE5",
			x"0000" when x"FCE6",
			x"0000" when x"FCE7",
			x"0000" when x"FCE8",
			x"0000" when x"FCE9",
			x"0000" when x"FCEA",
			x"0000" when x"FCEB",
			x"0000" when x"FCEC",
			x"0000" when x"FCED",
			x"0000" when x"FCEE",
			x"0000" when x"FCEF",
			x"0000" when x"FCF0",
			x"0000" when x"FCF1",
			x"0000" when x"FCF2",
			x"0000" when x"FCF3",
			x"0000" when x"FCF4",
			x"0000" when x"FCF5",
			x"0000" when x"FCF6",
			x"0000" when x"FCF7",
			x"0000" when x"FCF8",
			x"0000" when x"FCF9",
			x"0000" when x"FCFA",
			x"0000" when x"FCFB",
			x"0000" when x"FCFC",
			x"0000" when x"FCFD",
			x"0000" when x"FCFE",
			x"0000" when x"FCFF",
			x"0000" when x"FD00",
			x"0000" when x"FD01",
			x"0000" when x"FD02",
			x"0000" when x"FD03",
			x"0000" when x"FD04",
			x"0000" when x"FD05",
			x"0000" when x"FD06",
			x"0000" when x"FD07",
			x"0000" when x"FD08",
			x"0000" when x"FD09",
			x"0000" when x"FD0A",
			x"0000" when x"FD0B",
			x"0000" when x"FD0C",
			x"0000" when x"FD0D",
			x"0000" when x"FD0E",
			x"0000" when x"FD0F",
			x"0000" when x"FD10",
			x"0000" when x"FD11",
			x"0000" when x"FD12",
			x"0000" when x"FD13",
			x"0000" when x"FD14",
			x"0000" when x"FD15",
			x"0000" when x"FD16",
			x"0000" when x"FD17",
			x"0000" when x"FD18",
			x"0000" when x"FD19",
			x"0000" when x"FD1A",
			x"0000" when x"FD1B",
			x"0000" when x"FD1C",
			x"0000" when x"FD1D",
			x"0000" when x"FD1E",
			x"0000" when x"FD1F",
			x"0000" when x"FD20",
			x"0000" when x"FD21",
			x"0000" when x"FD22",
			x"0000" when x"FD23",
			x"0000" when x"FD24",
			x"0000" when x"FD25",
			x"0000" when x"FD26",
			x"0000" when x"FD27",
			x"0000" when x"FD28",
			x"0000" when x"FD29",
			x"0000" when x"FD2A",
			x"0000" when x"FD2B",
			x"0000" when x"FD2C",
			x"0000" when x"FD2D",
			x"0000" when x"FD2E",
			x"0000" when x"FD2F",
			x"0000" when x"FD30",
			x"0000" when x"FD31",
			x"0000" when x"FD32",
			x"0000" when x"FD33",
			x"0000" when x"FD34",
			x"0000" when x"FD35",
			x"0000" when x"FD36",
			x"0000" when x"FD37",
			x"0000" when x"FD38",
			x"0000" when x"FD39",
			x"0000" when x"FD3A",
			x"0000" when x"FD3B",
			x"0000" when x"FD3C",
			x"0000" when x"FD3D",
			x"0000" when x"FD3E",
			x"0000" when x"FD3F",
			x"0000" when x"FD40",
			x"0000" when x"FD41",
			x"0000" when x"FD42",
			x"0000" when x"FD43",
			x"0000" when x"FD44",
			x"0000" when x"FD45",
			x"0000" when x"FD46",
			x"0000" when x"FD47",
			x"0000" when x"FD48",
			x"0000" when x"FD49",
			x"0000" when x"FD4A",
			x"0000" when x"FD4B",
			x"0000" when x"FD4C",
			x"0000" when x"FD4D",
			x"0000" when x"FD4E",
			x"0000" when x"FD4F",
			x"0000" when x"FD50",
			x"0000" when x"FD51",
			x"0000" when x"FD52",
			x"0000" when x"FD53",
			x"0000" when x"FD54",
			x"0000" when x"FD55",
			x"0000" when x"FD56",
			x"0000" when x"FD57",
			x"0000" when x"FD58",
			x"0000" when x"FD59",
			x"0000" when x"FD5A",
			x"0000" when x"FD5B",
			x"0000" when x"FD5C",
			x"0000" when x"FD5D",
			x"0000" when x"FD5E",
			x"0000" when x"FD5F",
			x"0000" when x"FD60",
			x"0000" when x"FD61",
			x"0000" when x"FD62",
			x"0000" when x"FD63",
			x"0000" when x"FD64",
			x"0000" when x"FD65",
			x"0000" when x"FD66",
			x"0000" when x"FD67",
			x"0000" when x"FD68",
			x"0000" when x"FD69",
			x"0000" when x"FD6A",
			x"0000" when x"FD6B",
			x"0000" when x"FD6C",
			x"0000" when x"FD6D",
			x"0000" when x"FD6E",
			x"0000" when x"FD6F",
			x"0000" when x"FD70",
			x"0000" when x"FD71",
			x"0000" when x"FD72",
			x"0000" when x"FD73",
			x"0000" when x"FD74",
			x"0000" when x"FD75",
			x"0000" when x"FD76",
			x"0000" when x"FD77",
			x"0000" when x"FD78",
			x"0000" when x"FD79",
			x"0000" when x"FD7A",
			x"0000" when x"FD7B",
			x"0000" when x"FD7C",
			x"0000" when x"FD7D",
			x"0000" when x"FD7E",
			x"0000" when x"FD7F",
			x"0000" when x"FD80",
			x"0000" when x"FD81",
			x"0000" when x"FD82",
			x"0000" when x"FD83",
			x"0000" when x"FD84",
			x"0000" when x"FD85",
			x"0000" when x"FD86",
			x"0000" when x"FD87",
			x"0000" when x"FD88",
			x"0000" when x"FD89",
			x"0000" when x"FD8A",
			x"0000" when x"FD8B",
			x"0000" when x"FD8C",
			x"0000" when x"FD8D",
			x"0000" when x"FD8E",
			x"0000" when x"FD8F",
			x"0000" when x"FD90",
			x"0000" when x"FD91",
			x"0000" when x"FD92",
			x"0000" when x"FD93",
			x"0000" when x"FD94",
			x"0000" when x"FD95",
			x"0000" when x"FD96",
			x"0000" when x"FD97",
			x"0000" when x"FD98",
			x"0000" when x"FD99",
			x"0000" when x"FD9A",
			x"0000" when x"FD9B",
			x"0000" when x"FD9C",
			x"0000" when x"FD9D",
			x"0000" when x"FD9E",
			x"0000" when x"FD9F",
			x"0000" when x"FDA0",
			x"0000" when x"FDA1",
			x"0000" when x"FDA2",
			x"0000" when x"FDA3",
			x"0000" when x"FDA4",
			x"0000" when x"FDA5",
			x"0000" when x"FDA6",
			x"0000" when x"FDA7",
			x"0000" when x"FDA8",
			x"0000" when x"FDA9",
			x"0000" when x"FDAA",
			x"0000" when x"FDAB",
			x"0000" when x"FDAC",
			x"0000" when x"FDAD",
			x"0000" when x"FDAE",
			x"0000" when x"FDAF",
			x"0000" when x"FDB0",
			x"0000" when x"FDB1",
			x"0000" when x"FDB2",
			x"0000" when x"FDB3",
			x"0000" when x"FDB4",
			x"0000" when x"FDB5",
			x"0000" when x"FDB6",
			x"0000" when x"FDB7",
			x"0000" when x"FDB8",
			x"0000" when x"FDB9",
			x"0000" when x"FDBA",
			x"0000" when x"FDBB",
			x"0000" when x"FDBC",
			x"0000" when x"FDBD",
			x"0000" when x"FDBE",
			x"0000" when x"FDBF",
			x"0000" when x"FDC0",
			x"0000" when x"FDC1",
			x"0000" when x"FDC2",
			x"0000" when x"FDC3",
			x"0000" when x"FDC4",
			x"0000" when x"FDC5",
			x"0000" when x"FDC6",
			x"0000" when x"FDC7",
			x"0000" when x"FDC8",
			x"0000" when x"FDC9",
			x"0000" when x"FDCA",
			x"0000" when x"FDCB",
			x"0000" when x"FDCC",
			x"0000" when x"FDCD",
			x"0000" when x"FDCE",
			x"0000" when x"FDCF",
			x"0000" when x"FDD0",
			x"0000" when x"FDD1",
			x"0000" when x"FDD2",
			x"0000" when x"FDD3",
			x"0000" when x"FDD4",
			x"0000" when x"FDD5",
			x"0000" when x"FDD6",
			x"0000" when x"FDD7",
			x"0000" when x"FDD8",
			x"0000" when x"FDD9",
			x"0000" when x"FDDA",
			x"0000" when x"FDDB",
			x"0000" when x"FDDC",
			x"0000" when x"FDDD",
			x"0000" when x"FDDE",
			x"0000" when x"FDDF",
			x"0000" when x"FDE0",
			x"0000" when x"FDE1",
			x"0000" when x"FDE2",
			x"0000" when x"FDE3",
			x"0000" when x"FDE4",
			x"0000" when x"FDE5",
			x"0000" when x"FDE6",
			x"0000" when x"FDE7",
			x"0000" when x"FDE8",
			x"0000" when x"FDE9",
			x"0000" when x"FDEA",
			x"0000" when x"FDEB",
			x"0000" when x"FDEC",
			x"0000" when x"FDED",
			x"0000" when x"FDEE",
			x"0000" when x"FDEF",
			x"0000" when x"FDF0",
			x"0000" when x"FDF1",
			x"0000" when x"FDF2",
			x"0000" when x"FDF3",
			x"0000" when x"FDF4",
			x"0000" when x"FDF5",
			x"0000" when x"FDF6",
			x"0000" when x"FDF7",
			x"0000" when x"FDF8",
			x"0000" when x"FDF9",
			x"0000" when x"FDFA",
			x"0000" when x"FDFB",
			x"0000" when x"FDFC",
			x"0000" when x"FDFD",
			x"0000" when x"FDFE",
			x"0000" when x"FDFF",
			x"0000" when x"FE00",
			x"0000" when x"FE01",
			x"0000" when x"FE02",
			x"0000" when x"FE03",
			x"0000" when x"FE04",
			x"0000" when x"FE05",
			x"0000" when x"FE06",
			x"0000" when x"FE07",
			x"0000" when x"FE08",
			x"0000" when x"FE09",
			x"0000" when x"FE0A",
			x"0000" when x"FE0B",
			x"0000" when x"FE0C",
			x"0000" when x"FE0D",
			x"0000" when x"FE0E",
			x"0000" when x"FE0F",
			x"0000" when x"FE10",
			x"0000" when x"FE11",
			x"0000" when x"FE12",
			x"0000" when x"FE13",
			x"0000" when x"FE14",
			x"0000" when x"FE15",
			x"0000" when x"FE16",
			x"0000" when x"FE17",
			x"0000" when x"FE18",
			x"0000" when x"FE19",
			x"0000" when x"FE1A",
			x"0000" when x"FE1B",
			x"0000" when x"FE1C",
			x"0000" when x"FE1D",
			x"0000" when x"FE1E",
			x"0000" when x"FE1F",
			x"0000" when x"FE20",
			x"0000" when x"FE21",
			x"0000" when x"FE22",
			x"0000" when x"FE23",
			x"0000" when x"FE24",
			x"0000" when x"FE25",
			x"0000" when x"FE26",
			x"0000" when x"FE27",
			x"0000" when x"FE28",
			x"0000" when x"FE29",
			x"0000" when x"FE2A",
			x"0000" when x"FE2B",
			x"0000" when x"FE2C",
			x"0000" when x"FE2D",
			x"0000" when x"FE2E",
			x"0000" when x"FE2F",
			x"0000" when x"FE30",
			x"0000" when x"FE31",
			x"0000" when x"FE32",
			x"0000" when x"FE33",
			x"0000" when x"FE34",
			x"0000" when x"FE35",
			x"0000" when x"FE36",
			x"0000" when x"FE37",
			x"0000" when x"FE38",
			x"0000" when x"FE39",
			x"0000" when x"FE3A",
			x"0000" when x"FE3B",
			x"0000" when x"FE3C",
			x"0000" when x"FE3D",
			x"0000" when x"FE3E",
			x"0000" when x"FE3F",
			x"0000" when x"FE40",
			x"0000" when x"FE41",
			x"0000" when x"FE42",
			x"0000" when x"FE43",
			x"0000" when x"FE44",
			x"0000" when x"FE45",
			x"0000" when x"FE46",
			x"0000" when x"FE47",
			x"0000" when x"FE48",
			x"0000" when x"FE49",
			x"0000" when x"FE4A",
			x"0000" when x"FE4B",
			x"0000" when x"FE4C",
			x"0000" when x"FE4D",
			x"0000" when x"FE4E",
			x"0000" when x"FE4F",
			x"0000" when x"FE50",
			x"0000" when x"FE51",
			x"0000" when x"FE52",
			x"0000" when x"FE53",
			x"0000" when x"FE54",
			x"0000" when x"FE55",
			x"0000" when x"FE56",
			x"0000" when x"FE57",
			x"0000" when x"FE58",
			x"0000" when x"FE59",
			x"0000" when x"FE5A",
			x"0000" when x"FE5B",
			x"0000" when x"FE5C",
			x"0000" when x"FE5D",
			x"0000" when x"FE5E",
			x"0000" when x"FE5F",
			x"0000" when x"FE60",
			x"0000" when x"FE61",
			x"0000" when x"FE62",
			x"0000" when x"FE63",
			x"0000" when x"FE64",
			x"0000" when x"FE65",
			x"0000" when x"FE66",
			x"0000" when x"FE67",
			x"0000" when x"FE68",
			x"0000" when x"FE69",
			x"0000" when x"FE6A",
			x"0000" when x"FE6B",
			x"0000" when x"FE6C",
			x"0000" when x"FE6D",
			x"0000" when x"FE6E",
			x"0000" when x"FE6F",
			x"0000" when x"FE70",
			x"0000" when x"FE71",
			x"0000" when x"FE72",
			x"0000" when x"FE73",
			x"0000" when x"FE74",
			x"0000" when x"FE75",
			x"0000" when x"FE76",
			x"0000" when x"FE77",
			x"0000" when x"FE78",
			x"0000" when x"FE79",
			x"0000" when x"FE7A",
			x"0000" when x"FE7B",
			x"0000" when x"FE7C",
			x"0000" when x"FE7D",
			x"0000" when x"FE7E",
			x"0000" when x"FE7F",
			x"0000" when x"FE80",
			x"0000" when x"FE81",
			x"0000" when x"FE82",
			x"0000" when x"FE83",
			x"0000" when x"FE84",
			x"0000" when x"FE85",
			x"0000" when x"FE86",
			x"0000" when x"FE87",
			x"0000" when x"FE88",
			x"0000" when x"FE89",
			x"0000" when x"FE8A",
			x"0000" when x"FE8B",
			x"0000" when x"FE8C",
			x"0000" when x"FE8D",
			x"0000" when x"FE8E",
			x"0000" when x"FE8F",
			x"0000" when x"FE90",
			x"0000" when x"FE91",
			x"0000" when x"FE92",
			x"0000" when x"FE93",
			x"0000" when x"FE94",
			x"0000" when x"FE95",
			x"0000" when x"FE96",
			x"0000" when x"FE97",
			x"0000" when x"FE98",
			x"0000" when x"FE99",
			x"0000" when x"FE9A",
			x"0000" when x"FE9B",
			x"0000" when x"FE9C",
			x"0000" when x"FE9D",
			x"0000" when x"FE9E",
			x"0000" when x"FE9F",
			x"0000" when x"FEA0",
			x"0000" when x"FEA1",
			x"0000" when x"FEA2",
			x"0000" when x"FEA3",
			x"0000" when x"FEA4",
			x"0000" when x"FEA5",
			x"0000" when x"FEA6",
			x"0000" when x"FEA7",
			x"0000" when x"FEA8",
			x"0000" when x"FEA9",
			x"0000" when x"FEAA",
			x"0000" when x"FEAB",
			x"0000" when x"FEAC",
			x"0000" when x"FEAD",
			x"0000" when x"FEAE",
			x"0000" when x"FEAF",
			x"0000" when x"FEB0",
			x"0000" when x"FEB1",
			x"0000" when x"FEB2",
			x"0000" when x"FEB3",
			x"0000" when x"FEB4",
			x"0000" when x"FEB5",
			x"0000" when x"FEB6",
			x"0000" when x"FEB7",
			x"0000" when x"FEB8",
			x"0000" when x"FEB9",
			x"0000" when x"FEBA",
			x"0000" when x"FEBB",
			x"0000" when x"FEBC",
			x"0000" when x"FEBD",
			x"0000" when x"FEBE",
			x"0000" when x"FEBF",
			x"0000" when x"FEC0",
			x"0000" when x"FEC1",
			x"0000" when x"FEC2",
			x"0000" when x"FEC3",
			x"0000" when x"FEC4",
			x"0000" when x"FEC5",
			x"0000" when x"FEC6",
			x"0000" when x"FEC7",
			x"0000" when x"FEC8",
			x"0000" when x"FEC9",
			x"0000" when x"FECA",
			x"0000" when x"FECB",
			x"0000" when x"FECC",
			x"0000" when x"FECD",
			x"0000" when x"FECE",
			x"0000" when x"FECF",
			x"0000" when x"FED0",
			x"0000" when x"FED1",
			x"0000" when x"FED2",
			x"0000" when x"FED3",
			x"0000" when x"FED4",
			x"0000" when x"FED5",
			x"0000" when x"FED6",
			x"0000" when x"FED7",
			x"0000" when x"FED8",
			x"0000" when x"FED9",
			x"0000" when x"FEDA",
			x"0000" when x"FEDB",
			x"0000" when x"FEDC",
			x"0000" when x"FEDD",
			x"0000" when x"FEDE",
			x"0000" when x"FEDF",
			x"0000" when x"FEE0",
			x"0000" when x"FEE1",
			x"0000" when x"FEE2",
			x"0000" when x"FEE3",
			x"0000" when x"FEE4",
			x"0000" when x"FEE5",
			x"0000" when x"FEE6",
			x"0000" when x"FEE7",
			x"0000" when x"FEE8",
			x"0000" when x"FEE9",
			x"0000" when x"FEEA",
			x"0000" when x"FEEB",
			x"0000" when x"FEEC",
			x"0000" when x"FEED",
			x"0000" when x"FEEE",
			x"0000" when x"FEEF",
			x"0000" when x"FEF0",
			x"0000" when x"FEF1",
			x"0000" when x"FEF2",
			x"0000" when x"FEF3",
			x"0000" when x"FEF4",
			x"0000" when x"FEF5",
			x"0000" when x"FEF6",
			x"0000" when x"FEF7",
			x"0000" when x"FEF8",
			x"0000" when x"FEF9",
			x"0000" when x"FEFA",
			x"0000" when x"FEFB",
			x"0000" when x"FEFC",
			x"0000" when x"FEFD",
			x"0000" when x"FEFE",
			x"0000" when x"FEFF",
			x"0000" when x"FF00",
			x"0000" when x"FF01",
			x"0000" when x"FF02",
			x"0000" when x"FF03",
			x"0000" when x"FF04",
			x"0000" when x"FF05",
			x"0000" when x"FF06",
			x"0000" when x"FF07",
			x"0000" when x"FF08",
			x"0000" when x"FF09",
			x"0000" when x"FF0A",
			x"0000" when x"FF0B",
			x"0000" when x"FF0C",
			x"0000" when x"FF0D",
			x"0000" when x"FF0E",
			x"0000" when x"FF0F",
			x"0000" when x"FF10",
			x"0000" when x"FF11",
			x"0000" when x"FF12",
			x"0000" when x"FF13",
			x"0000" when x"FF14",
			x"0000" when x"FF15",
			x"0000" when x"FF16",
			x"0000" when x"FF17",
			x"0000" when x"FF18",
			x"0000" when x"FF19",
			x"0000" when x"FF1A",
			x"0000" when x"FF1B",
			x"0000" when x"FF1C",
			x"0000" when x"FF1D",
			x"0000" when x"FF1E",
			x"0000" when x"FF1F",
			x"0000" when x"FF20",
			x"0000" when x"FF21",
			x"0000" when x"FF22",
			x"0000" when x"FF23",
			x"0000" when x"FF24",
			x"0000" when x"FF25",
			x"0000" when x"FF26",
			x"0000" when x"FF27",
			x"0000" when x"FF28",
			x"0000" when x"FF29",
			x"0000" when x"FF2A",
			x"0000" when x"FF2B",
			x"0000" when x"FF2C",
			x"0000" when x"FF2D",
			x"0000" when x"FF2E",
			x"0000" when x"FF2F",
			x"0000" when x"FF30",
			x"0000" when x"FF31",
			x"0000" when x"FF32",
			x"0000" when x"FF33",
			x"0000" when x"FF34",
			x"0000" when x"FF35",
			x"0000" when x"FF36",
			x"0000" when x"FF37",
			x"0000" when x"FF38",
			x"0000" when x"FF39",
			x"0000" when x"FF3A",
			x"0000" when x"FF3B",
			x"0000" when x"FF3C",
			x"0000" when x"FF3D",
			x"0000" when x"FF3E",
			x"0000" when x"FF3F",
			x"0000" when x"FF40",
			x"0000" when x"FF41",
			x"0000" when x"FF42",
			x"0000" when x"FF43",
			x"0000" when x"FF44",
			x"0000" when x"FF45",
			x"0000" when x"FF46",
			x"0000" when x"FF47",
			x"0000" when x"FF48",
			x"0000" when x"FF49",
			x"0000" when x"FF4A",
			x"0000" when x"FF4B",
			x"0000" when x"FF4C",
			x"0000" when x"FF4D",
			x"0000" when x"FF4E",
			x"0000" when x"FF4F",
			x"0000" when x"FF50",
			x"0000" when x"FF51",
			x"0000" when x"FF52",
			x"0000" when x"FF53",
			x"0000" when x"FF54",
			x"0000" when x"FF55",
			x"0000" when x"FF56",
			x"0000" when x"FF57",
			x"0000" when x"FF58",
			x"0000" when x"FF59",
			x"0000" when x"FF5A",
			x"0000" when x"FF5B",
			x"0000" when x"FF5C",
			x"0000" when x"FF5D",
			x"0000" when x"FF5E",
			x"0000" when x"FF5F",
			x"0000" when x"FF60",
			x"0000" when x"FF61",
			x"0000" when x"FF62",
			x"0000" when x"FF63",
			x"0000" when x"FF64",
			x"0000" when x"FF65",
			x"0000" when x"FF66",
			x"0000" when x"FF67",
			x"0000" when x"FF68",
			x"0000" when x"FF69",
			x"0000" when x"FF6A",
			x"0000" when x"FF6B",
			x"0000" when x"FF6C",
			x"0000" when x"FF6D",
			x"0000" when x"FF6E",
			x"0000" when x"FF6F",
			x"0000" when x"FF70",
			x"0000" when x"FF71",
			x"0000" when x"FF72",
			x"0000" when x"FF73",
			x"0000" when x"FF74",
			x"0000" when x"FF75",
			x"0000" when x"FF76",
			x"0000" when x"FF77",
			x"0000" when x"FF78",
			x"0000" when x"FF79",
			x"0000" when x"FF7A",
			x"0000" when x"FF7B",
			x"0000" when x"FF7C",
			x"0000" when x"FF7D",
			x"0000" when x"FF7E",
			x"0000" when x"FF7F",
			x"0000" when x"FF80",
			x"0000" when x"FF81",
			x"0000" when x"FF82",
			x"0000" when x"FF83",
			x"0000" when x"FF84",
			x"0000" when x"FF85",
			x"0000" when x"FF86",
			x"0000" when x"FF87",
			x"0000" when x"FF88",
			x"0000" when x"FF89",
			x"0000" when x"FF8A",
			x"0000" when x"FF8B",
			x"0000" when x"FF8C",
			x"0000" when x"FF8D",
			x"0000" when x"FF8E",
			x"0000" when x"FF8F",
			x"0000" when x"FF90",
			x"0000" when x"FF91",
			x"0000" when x"FF92",
			x"0000" when x"FF93",
			x"0000" when x"FF94",
			x"0000" when x"FF95",
			x"0000" when x"FF96",
			x"0000" when x"FF97",
			x"0000" when x"FF98",
			x"0000" when x"FF99",
			x"0000" when x"FF9A",
			x"0000" when x"FF9B",
			x"0000" when x"FF9C",
			x"0000" when x"FF9D",
			x"0000" when x"FF9E",
			x"0000" when x"FF9F",
			x"0000" when x"FFA0",
			x"0000" when x"FFA1",
			x"0000" when x"FFA2",
			x"0000" when x"FFA3",
			x"0000" when x"FFA4",
			x"0000" when x"FFA5",
			x"0000" when x"FFA6",
			x"0000" when x"FFA7",
			x"0000" when x"FFA8",
			x"0000" when x"FFA9",
			x"0000" when x"FFAA",
			x"0000" when x"FFAB",
			x"0000" when x"FFAC",
			x"0000" when x"FFAD",
			x"0000" when x"FFAE",
			x"0000" when x"FFAF",
			x"0000" when x"FFB0",
			x"0000" when x"FFB1",
			x"0000" when x"FFB2",
			x"0000" when x"FFB3",
			x"0000" when x"FFB4",
			x"0000" when x"FFB5",
			x"0000" when x"FFB6",
			x"0000" when x"FFB7",
			x"0000" when x"FFB8",
			x"0000" when x"FFB9",
			x"0000" when x"FFBA",
			x"0000" when x"FFBB",
			x"0000" when x"FFBC",
			x"0000" when x"FFBD",
			x"0000" when x"FFBE",
			x"0000" when x"FFBF",
			x"0000" when x"FFC0",
			x"0000" when x"FFC1",
			x"0000" when x"FFC2",
			x"0000" when x"FFC3",
			x"0000" when x"FFC4",
			x"0000" when x"FFC5",
			x"0000" when x"FFC6",
			x"0000" when x"FFC7",
			x"0000" when x"FFC8",
			x"0000" when x"FFC9",
			x"0000" when x"FFCA",
			x"0000" when x"FFCB",
			x"0000" when x"FFCC",
			x"0000" when x"FFCD",
			x"0000" when x"FFCE",
			x"0000" when x"FFCF",
			x"0000" when x"FFD0",
			x"0000" when x"FFD1",
			x"0000" when x"FFD2",
			x"0000" when x"FFD3",
			x"0000" when x"FFD4",
			x"0000" when x"FFD5",
			x"0000" when x"FFD6",
			x"0000" when x"FFD7",
			x"0000" when x"FFD8",
			x"0000" when x"FFD9",
			x"0000" when x"FFDA",
			x"0000" when x"FFDB",
			x"0000" when x"FFDC",
			x"0000" when x"FFDD",
			x"0000" when x"FFDE",
			x"0000" when x"FFDF",
			x"0000" when x"FFE0",
			x"0000" when x"FFE1",
			x"0000" when x"FFE2",
			x"0000" when x"FFE3",
			x"0000" when x"FFE4",
			x"0000" when x"FFE5",
			x"0000" when x"FFE6",
			x"0000" when x"FFE7",
			x"0000" when x"FFE8",
			x"0000" when x"FFE9",
			x"0000" when x"FFEA",
			x"0000" when x"FFEB",
			x"0000" when x"FFEC",
			x"0000" when x"FFED",
			x"0000" when x"FFEE",
			x"0000" when x"FFEF",
			x"0000" when x"FFF0",
			x"0000" when x"FFF1",
			x"0000" when x"FFF2",
			x"0000" when x"FFF3",
			x"0000" when x"FFF4",
			x"0000" when x"FFF5",
			x"0000" when x"FFF6",
			x"0000" when x"FFF7",
			x"0000" when x"FFF8",
			x"0000" when x"FFF9",
			x"0000" when x"FFFA",
			x"0000" when x"FFFB",
			x"0000" when x"FFFC",
			x"0000" when x"FFFD",
			x"0000" when x"FFFE",
			x"0000" when x"FFFF";

end architecture;
