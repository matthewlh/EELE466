`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
DvYvlhLNE4Z5g/PdkH93s94O7DQWjXfApiLaWuzUtF3pkLENvNbvFLUfGKoSbNAW
isekdYisxWmbgLUZM1L1zqnRA9CzZxtbh0xz3Qef2w0ia6QNNS7Au/KyU7MKhVKt
2htTmnLslGN+JoxCxdCibcIEgvxbhepDnXdBj36dlm/Gsaw9NIzXKE3hdjguqr00
ux6zoREgeC+sctIoLq2y68w6xmTBF0qdybXC+gUGRj99YvboQiVf3edHLIaoZxeQ
KXg6crBk1NXgQqGlDzQNgQwuE1XOouB/4Ry9hKBg9Js4RDSaKi0ZKawKWgpUQMfY
1YZptsHFX11syhtaAhg0W+LLOHNJsH2KtRNJr+dyoWN50iYFC+eyfw1phcuWmaHB
bpqcW1xaXDziIu06mjNZtB1ElkQJ2C0GqFfLq6+vOgTPD3TKfG425QQpBDstUbRB
syTmKZecE8LaCrsCd4YguEYUH/rjNGCLgCdEjeN2HKAK6JrNzHgmKnEhKl39wjvp
2C7aKSQW3WoOAMlzwfrTY273DNLGpv0Tt2vgnmjBHucMJqIxU3GN7y9RfXoK9j/a
zgDsfMMGFfQZGCy3CSF1Vo83k354CuE0PxKvvRMdAVvmBGOjKAKMRHZ/RjeE1c0e
fb+f/+e7yfT+jpS18Rq8N6Zu7bsZaVQiDTIb3m8G6A0clYSJbEntr5FNLLQCR1E4
Q9Noj6Y2qAa1gOok4pn7zI7wpnxJds4EX+i8aFlNWfBQAp3hbJpbhsU6mm/vV/iH
T+T0WtQUD6k/SqRLjAuGOeGhT7y3Qb4vwDhXSmPMcbAK0bdHaxXRlKBL/+WN6ZUg
qoz4xaf8Jvw8VbHHKiE0H1LvQjsjsnTyq+5vJnE2rdD6s3RSj3DDfUVCPjrRSyTD
UhW6jKLPqKqz/LYXyfowLkSzy+LNfnu6OjoBPIra6H9JIa/G457gF7gGHhMLbSco
6ru+wRl4zv+GW5/15GJvD0Xqw5bmOoZcFrjk67gx7FoZ6Qxhks7xCKniM3n2DMif
nvsP98LE/V8N3TN6ExDbzCv4rJJwwpzdNXsRsPhGRK/CcGME2DD4EBckjVLr5EOv
9T2YtjlPPYalujE3ZWg2Wxbqfa8Zcnc3Lgi4Z7mvy+/Au5JFZx471R5nBPkocJQi
ml58L7oLvFrBqBrqcLfwYhVU4N6O6UigQkbQcP0X7DeAgxYHnh5kjJe8f/hrywDb
y5XCALKLZXurqLCr4uy6qXdMkQieJUveCl/JRgawmYU81tnzDFxU/r26hJG6Uvut
rAdtXPACZDNkyI743UCLNFew86Nq+OC1PEkfmUR+ENsdR9dtQ4HSzmDpWFP8jO8T
0RDbpliHlOGPJ3P4QVGQRhmcte6MewN7y0xAOaML2SpujVy3Dp0eU1+/gV2n5e6J
zksvgQ+9E45YpcBKGTIENmchdhdZpJUfgN0c9OW7vIp3A1yXVkJjt5l1yhsH7cWx
KMITvYIlntlesPSKB1GbujSe3LBi8GTXRTbz4fHN6DLQbYAyDVOxRDKGyH4Dtxsb
51ETwx8Q9070ebSf1u+3Gg==
`protect END_PROTECTED
