`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
vy2mBF1OURbVbItdcHZrcJgF0YWCvTrRPWCgJPzJt95+itIioeXMXHsNO6yEtaNC
7kaq/3g1ZAfGGB9Z4xrZqGM+DSXMmj3x8y9Z4YEe6iG0C/zyn1RW2KLOylxeliFr
hNPjXFdoRaNikkDD2knrTU92lO4bnVPFBxpn0yhRCWCZ6BezdlHu07cF7pG/qY9t
RoNxOWRAe1jM0dtjxjjex7F+ikF5DU/jWZhWqzEHNptFZTL6zCZEwNVbhYLgK3SM
OZCpB+gf/3TWmD4pJcoq1YbdIOBdrU0DknwFWDv1BLpkbTnEjlx3Kx+XZgBDFy8Z
Hl39EU5+nrA55Q59mxtGOrqK44aP8QHF1KeJOAxGcQKB/9lw6OcghI7ao6dsjFg5
7tBb5OEOJ7ZtJ7mz/jUaLiYcNGSUmZ497tQfN+LubEk1AP3U7N1ahSZ8B5FGp2LT
Foq1ADSA8a1qVbPn84yA2ATUvpKQ1U4oZqKG1DWtZSkUaTFBYD8PMeJ8iAdaeFSf
xS+EWtGow4FGKFbYHW0aMnKbONetAgup2IYnYbZLV26R3UlNdXQLikcAb7SsM+OJ
wkWYZOXmcanriovF4ay3cnySWg65qzrq+stSi153ESeOnYRPakQElP42dZ0oVn7p
pV8PMatARuUIBKe0tgwGBDgFUSUGyTC0NvYiiCyIoWEbBxmwzK2Gst5Dg2YJeOPk
3/AAd7j3OJjlrmUacmfvPbIj8S9YAJyZhYPANzgzGMdkzEZpwIN0d7Mg0P8JQJKn
l9F3YniWb0hnT63+jTnOA96mH1sMZdG9knV013Ph0nTDd2Ap8xv8Ye5tyexfDJSI
+ovser45WDX1+FV+arZaGO52j5PgCV0vWCvsl+bM7H4qa/0Gz/inqJaT5AmTx3Vm
YN4qtKQHa+24wZ/QpvUJu7HnrNB1UJqeQzOHj6ZJqOm1bZBKZmbIW5ZEkWuylaqX
RPBb5Kwzk46hW8epXB6s2rkf8SPBEm90Tpn/KOfEzdeZlnYOvwPculXa+YBxV06r
c+bc3VMRHFexm1B/uJ3CFnva5ELgYQAuGF/Y/unSXKJIigukH9PzCAnkVEj+f1Vn
git37bVMZzyU1tlDnFVcEIHIOSUsOXDs9rRQ70B57LHTz6hyJGpqfRwRztUouQDy
BogV+H4TBhRO31NAUS3aEjpdK7C68og8GV47azue8Pdl0PnVtDPAe0YQXQf3nPiH
48AUarghpzWTrC2DX/Fuhdz2HUIr1TmshmyFjFz83t7qsu4Hw7wosPZ/9saYQ9gZ
L0epT02YzwQYuE9+uhm9xoDe9lqxxdDT8h0NqFpvMegLfArbSSs4V5TnDBWGEx02
hHe6V6ryoFzBco5N6AqwWPUw9i513VfP+YbdGkscIR3kWqGYFGxF1+vRC/dtDur6
7WFHGGJew/cTxta5n1pzzxgtyEf686gxQRHqUl7D0WCzKEJBxXkkZUEWayWhXfmW
YkH8HmHnYQRnSGDd6CiDSr8EBXN8gjg/vSVTqKtQTYLdpiv+SoCb2SaRy3ducdJt
ra8ijOjctvlY01p9UTJjZA==
`protect END_PROTECTED
