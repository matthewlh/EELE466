`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
v/8DCYPTbcB4lW9R1hbzIm1MMbYXcXcHqaWTtQmQVnpFSlHL8C34KKksG/ElEv7A
OgJ1/VpVk6Ns39WIuehrFSd/8RoWhbqac1RDrp5cke0MS+fEPZORtfecDDdcyIvM
bpcwEQp+v801slc2KmarULbiXSWR0X28Ty8EpqFp4utew64l1GON8AjvXSYBUx1+
FhxN9fX+Tg/MldbMFpFuAc2Lp9tuLR9aDR41aSIs7v8qyzc2H+I0SUWj/QHuVO1w
svWEKp+K41DuYOuBfs8nRoFp1nrpTXH0tCVhsZeA0G8KJHSEvLsGmRy+st3LtiiM
YvMZ9JhcqA0NWv+ffHDJhh9uSG8XBUf4h2EXnFR+SSJv2R0blYiNBXi6aarufrZC
PqKR4nR4/E6UP2nioEba3MoEOn9GoYsURf6q+xnFrLqRg6GDHkPPbR1I4peI3uXc
e5mwFjtkLVWn5si+Dia/hwnGwmk2yoWFziHCwDmoSqVIeroXATJmcob7l7FlNLGZ
FCgvLI8ekInZy/AtqSnxCe22hwA671irjkYw2gOcpXwI3YFf3SlY4jYoe+8kwswE
1GFMc+rB6ogGpk6bjT3a3equHt6r2QuJoT4ci90NgB9UylcM6khc8jyzFQc2LO+p
+b9W9T4ZGf+exAICiau/ErG/fGXOwPsbYtjZGYUrGAYcS313yZGfd6f+5lCLRJLH
63IKPmrtUnASJq+avpi5h6r3odyyQzDSYEdPUUygStf+F8seib0t0vavlKTeAykE
6JNxK5/vG2A5X7JGmPCRuqWOfVxDiZX6zalKmXpjnx8n1DF+vqIQKgTw6J2Ywbz5
tI25lEl8el0GhDzeHh5X+R5KFy8ySxXoOSli78D7Sspan6ZOBLkFtWzGzJH45HpU
lOJo7wyMx8TAftpdnxkWsLRkNgFYmwO/Pwe5EiKE6dyilO2So03HYJSQwyAK0MiV
ZBDB0C5AKr9OpHm1JAGpIoD4evuv9g3Y8jd0FyXEcbCuw4zg1GlgnF2wBGnDUsGm
EGLaTo65RjT7Y2b/NcxS6x9l9BoBdbaj+zTK3PdSX/FbEdci02RDMKqqN1OL3U2x
F8MNwqk2LjndkSyglFG/H4vFJFLkRFMt+eLTDKJWFp9+/OFWNfOefpSqBNTLPF6T
Xjoc0VH3Dcx9+YerSy0OPq0q63H8qzmmoOLXr/zox6+/arlix9XjwcHw2Ndf61MK
KXVW8fPaiJQaKjP2y7yTGbxvXR6PGJRVDiCGJPdQaTxZZCfI1u4aW2diMuD2hqW+
tBLf6/p8pb8mi3fmAr165ZXY9IbWAQIpLCBY4KRXXP1MuGcUzDCHJvFmOc212h44
R7UyFYzqQfynjfCIla7U5iqdHWtRxOSnZ6d+sajZ3fXQ5D2eJ670o/CULzWek4sv
dnnMwJmo8Og75LanRWnBDlTjVUHBaKhC+4CnLShUmYOPGme8NoSkl0J8cvewILgI
RV0kMt04hXA8S5YwF+J+s6DQwlWcPZPZD8vraSXBsyJyFu1/uzpAO5p7wE3lgqka
ppMYmtddVAn2sW0j5S4aNGf0d/amdlAFGPQhQ3XEm7nC9H1tqWfFDURYTtn9mAmp
nsAFD3+0w4FJJr/zQ54g7c7EEx48pRsu0TW15fHVqG8GUeXlHZo0WMsWgcGiQJHq
lHaiWlXEz9BT/NBKholYigl5N1AzeyFXm/fVMaWUMEW/Dj6MJHkMXX9YYQPCZQdw
1gKnrIB3NIhSAMNEU+8/seediMCA78+l9mRdc4pRM2nzPYlw8xHjS8v1lnvDHmFr
`protect END_PROTECTED
