`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
GOtL+bizVD4lP/KYDjLFPAHbpF74hOTe5bcT3KLuEJJ1y9Vs3jIpEapc4BRLbNGd
BqMknuB/5tni+ywC8OhzvFl8GhUxcobn77mzF1PAKkhdfFhPZBXELGHFQU3rrAZl
JMW6D1134mRlvtbNcQPpYwV9UROE7jM+h3Wk+LnYnzaBIq5yJRVJqPw91tUj15lT
z7ul5YksDZ2j+0BWgKfUsW8lL/iLZ6FQnzaSF5DUzUt8WwDvRzmtMmij/pFc1YuG
jUmJP2ts5te1Y7uRvFqCjsEH9BBE1SFxAXNj4ml0ZsKgC+1OBVDwi3zPhWBjVIbl
IoxZe4M1mWZc2M8WqElwVJ/+Fg2PTwn+FXrm8rXHA7ycMvWOyCFf0qLTevBZ3Ikm
H+4Y+rZ9rDqAtq1ny0fmZfafPARIkHMLR/aVXVztl7G2/oRM6Az+45mnGZgctpSW
LYRbKoH/+ZL5i/JxcC08vlZ0XFAcnopcI7rrbA7xiS+tUNARYbac0d9J5faiFKS1
w7Lw9j/XCykYzTUzwrzIndf6ojKC8m3r1s7uOIKsWAL35Y55qUlbm/lqqCJ4Dlk8
zFDPjrBReASzH6kSoD882Wl1P0EIUNoKUfgyG005xkfAskJ4WEqg0vu6qbHS2ZgZ
sO2wR26fG3rMP6fpavznzISAH6Qj2BbId/fC7raux72A1ReGsTfXRgolkNAE83x+
f1q2J0nFcCS+RGC8GEpF9nHKqK9vHEWCzr9zureShfIsdG/1wOXuuNX14JP/06oH
tb2zvDCNi85PxGa11TITyAhmWNu1ve0CZ7OAnXMvmQt/J5Wof1e3s4NL96uoQRc4
OlXJbA8kIYPkRVwXog+IGyqPzf3OO7oaJ7Kq6k3LZG9WSHLGMCnX42HNnqogpF6s
uSpVCyXcuonrqPMjlmILqDwlyT4tSyP6EkDCbKsWUQz+P1tX9uyCQOy1gNWcf/aj
yplbuLmm4Jy8rD6VnglqMJztn2vN6I9U++k6N21qS1qKsRT238BhXOzFAKAi4y5R
AGvsqZOOOBTpYZ6yPJG04w3Ysf9v+8Ua+A9zujV15h4TquMUnIV6CdewQsSjPR1v
RL/uP0uBKAwZq0IOuGCeZ/TMWko8UfHHjHtrGl5xOMaVwKqrkhsthNM5OrRKlZcX
wa5xUo945mkdDbwyaTCwYJrB9/YjgI1qv43K9YKrsKZEX13LKuzw3EBEU9P1bn2w
03wICGVar8ZS9Kb9lJexKg3aZ5GTdisGjY8nXoe3RKFSHea5y9AXn4nj5nbz1UF8
HU0hh87ovf4fVIybYADX6u9UqdhAfANCV+cwOjKlxKxWZv1KeTkf12Fx7WBl8PQ+
/PKarFWxiTpO+3fdWPAvKm7KAnQZ00zqS6alD88yglWlJiZ/Vgdh7ONXmMZk4zjz
kFWgKvAZDdpekTV3G8d5Uh8F7eCKObi1TS89UY8q8gPLhAzMAMOspmkNE6UCtm0M
RasMjZF+q/ebfVeaD41ZS6UVxQt1mWIqkUOP8VlbEs9RNEwyVh55KwhKd4vqYN+n
qLFPkrf+uNY5tfyZi1gCpkB70rJZhfdLsvdKIqF+NNqqy8RP0siuyK/qBTm/Qvmk
zUHhPFQXPRi/m4u7qauWNRj3W/ClfDUFyMcMxjWX0aIeI2ya7CuiG2TpkxEb1hLu
xIrYmvKr+TLbDZKt4g9tnQ+Sh12OY82FqSZHifoECK+8XS9/x0s7peF3zrhc6mYK
4mAKCOFwdrZVqg/EG6v7a+vmO+4kNeSrBhv5PansZo6jx+pnmOJBmtFzplRINK0J
9ITuNv6Gruu8cInghvF3G9c5mRBL2QMf75qRnn7GUKBxTFvSLIdhy8jQE3wtA6JJ
plZQTy+GyPwNlhd0Tcp381Qaq2sXsI2NwPFTWddASnuwRJc0BgtNh0slrGPguQlB
NWK+S92lKoE8dLFvAioRTgUaRj02nlq3GFIVCha6Tje+LoM1XRCiwGQ4OOgWJEv7
18oXYn0Kq41BUX0Gx48UTGwdDNmmCG5yafWNk07kJ9OumEAG3RSa7Ft//2Ar+F0I
3465uvlKpwMNkuISk0NICYWM0IQqpY3rRYgZJ5CmALw1eo7QFEgUpU1li9WFsN0h
XJJvY0DzR0Z4uQ11onyJsLhMUKIdmA11XA1/mPpUy5QN26m6IpG9cKe+88pFMzXG
dcZSusBbXsuhUBDURV7qcnSBp7zhsKVTsSKSD7dIyxe2BMyWFmAcBwi0Mdsa8oKc
4rn3sdooym5eR697gIPynqwcP52rSfbmGqFfkjpgKKsYhp20iBaSwaON6/bsLXKu
scqG260zPVinYhlXCt/pDvXxepwT/E3u0Y9RJ7MF6Zb+cMMhSdq4jzVHSXNqf3rM
OVbrifUN7C53ypcl4QXfMeNoTnSnnHoQF4GzxsSz8KGKRhX7apHOI1xUoyouDcM6
B1aoShDrn+aQTKFLVhGRV+7W8+JNqqSEo031t2WWpXurWfDRW23fb1WlcsVs5wYo
vZJ4nYO3vCf000S2b1p1tcZiL/3oOHlf3qIUxOQZzX8QgCp4XHi62B9iIGAx5shP
tlIZ3hY8Mw3Ihca5dPNsT3OWuPoC5OcX+4vQgWtEv3cKQGUbkyYbP7LF4DckDOvy
QMy616DpUv+xrPa1WFFfUdJZS8YU+BviQ/L6aX6nChMk0pQtJ9RbVCQ2G0KQiQ+2
sgfYfWK6nRCZnLActjV68vBgGhm2zBLD4q50RBPBNdorLLHbZ/GvX4y/MKKklsti
gM4eAEZCkQcUug7TDoH3OdmYNtBblBOtjdVD9fkCR+q3fAeHo4aztHEOYt3dvaJw
00XPraycVdNVddp4KI3JIHfiooABjDu+KxFzQGTs0+9niLCeUj4IZiPl3B4vhCd0
JEsPUmUCKDNRagGwivG+tOn5PKMqysfXD3qS/BP/5RilXCAhyQgwAEsngfySPJ7h
VHWfoD8YYMPW/mKMAI6vVDtyqgvWinHEiixO/y3YRjd1BSKgg0rCbRemc/gTbiDl
9BPrQ/Qe3+kKmChFm4GleRxC66GvGkCh8jpYjXh7vq5vbut9lQdsajnNL7HAOw0+
xmpx5UKmdKsLuKTtJVeDEdGb8IVE4dkS5UntFW7WGh8kPx/gM/w23yL/ODOu0jCB
M6VLb6xvIlOiijDXDBY7mU6SQygjjxEYRrPE0RjB3u79lKwUdgbJ2BR/xKtBYDSJ
WZ0tJQqjOmHbq9S911O0SRTOPWyCcTbLrQuCaqXXwgMNZKyWJM9H51m1/xUeLoQW
F0XQMjhXHPXwmVrc3ZixnSnTLdra7XN4XCipjPAeJXesPVcpTAYvDK/XICAvktpf
HkXK++tYLyPTwr062y+40MikC6K036pJpxTvC9OoAQbNEeuS7ePgg541BT0KF3t2
XQIFWe/F+MtmaodiAX2DckEh9AhO/5RnOSDqHhQHQq34FHFGDeYRK7Mv4Ev7Pmr0
ekCUl72a8qqPk4h/fTkmtiiy6Cn5X3xXnBDV+nHZO3h4XZ1pySqfDy/NjLINL4b9
ZKHw151JqMTxwW2F2CoPwwxujm5JZvXy4UwdP0yJGym20i7XdGXMlG+79qalMtHp
vg7dRNOCNiIrhn55f7RH4l36wGKVwJqDksF05ZpcbUn742+DVd2N1PiaTK4GIdtE
uDS/CZ1XWFiSViJsnlIy9maQmKNeQQUL4wPzkOqhosPW+xX+qc6ZFp0d4WfjKMMw
A6fNSGMymjimzkoMIuqgo5HUOs+QaLbDKh3s/NRmoDoANHtuhaWrgoRn1lL/qeuo
9vnulM4qVP+ZHL5fNIVK4y5GLmSBpzWiB5DgBjTggzdUbh6mIYLrnEKh2+OYsdos
+mhO3F+ejrmp20ExkyEMiDGbJjlDy5XBi+mHdCC6fl9XinxGwCovzhpmi4ZPOtFm
rEd5JKCx6qn7/IcFhLvdrn9czS3TiKgclaUGCLwYaG9rHibIWRQY3Y2iKvgEzlHG
2NbN5H77Ahi93PDZh2ZovnW1jQ5Ez+4HevN2XkAgyLv4+ZfvtUqc6D+PC5BVXE58
FecBRw2OykW7/oWLzE+aV9BynY9LAzqktWK13DtcjP8szvhEnHMWRHe6/8AaUFHF
991DkKAKKr9idNa3nTbcPmnftNNFeL+ZlBhqRRNh0ax7ANwE2uqTnvGNyvKMJ4We
0O6nSkj8oHScrpDR77mtcKSZrgB1Wsw5uqxF/mUDBc4CjpUPBArnOH/id1UP5Nav
MgZYFwPW2Y5mXx1cSSmBMYct2yVQlEPb2iHYHU0+yS/ufXpttguEGpmyOTK349eL
evrF9t543TP/QDWD1GjHluNd8X1umKHqlFYASsRTunHNEZd8D6VcCF+kl9jZ7QNE
XF17JIzNu0UvXVVMELrmoMMEZK6wC6iMdOC0Vn2c7lSUWAF2S/ASoXyr7PS7/8gH
gUv1peOr+N1VvzMARUMXbzyPqrqzsW8PYpOVWIoamgebwWpZBhaka2C31sz/9O7h
rI/P/z/RQcfEhZu7YR/UPBKZdQTBOTWTJ7a2haz6es5ZRJO9WDROZ7U8qm6cgW6G
Ichf1V+XfKBHzflXd0C9Qd4/ruE88f7mgYfzkmTdgLbEPRbsQW9GzB3lyfaJHLAb
XX1zJNG/T6uTbFympg9pVv1D/xRX5z97UUvEf5xsThq4K5YSSpRTgMedpGKQEdAb
zo2tBZHtPaHSqwUk4dQbvjLb+8pTVRPsn55GO//G2i/cA98TQOgMWE7dJL7gRG7+
fCb7AvILMaIdWakDEM3F87XdOh9YS8yASZWSOqbmQgThSNakfztQZK2XlcV7z/wJ
cjaPyQxdOTfXLtrvE5/bujqAI5k7LtyWSlFz7q2sLFxEmjENIVXNzFekP3+ljn2p
X9NOFwOZa65UhMHUjgwNGEWb8c58Eaj3EbQNSgeW311aotJITkhx2jvwY3g/yjFg
zVJSYHhz4C0i+cz7VUdiXY2fZ5gpijhkAk16HifIpdFXCbVWrEtTTouuapIdGLHY
OVoPx0D7nzTlnrDtTiUIKVYxtg7eAjh+fNNMc0YJF8c3LR/MakFE5M4uKhqydepL
kQNvNiIeWwnsIJeESBJdo4cpnWtQg40m2GWmqmuIe/lugxLn+/uMcXLjYRvqva90
Zia79UIXRdtM17JPR6YbbZAnTAPnwUZZG33/2P4iNb3pLUlKC293zO5/x6UQJdKA
dPSENzIOS0JLncTWqOoL7Xd4fmapWoAf3Ri+RQXrWiVcCqgkeLic8TOKOldPMtpY
6bXffzcgbDk00rZYaWDAD8TPgdfIc/Z+NMszfq6tmjAFM5Ko4tUAE0TN/myeg+7D
LAvPKv1e9SzFqx87zLVrt09FlXVTcWPrM0PUfAOfn+Zo2Kh8+2R4pyYq1bOVOP6g
dxFPzNdSNLw5oPJ0RHRnm1AlhnLPzhJvPH1jeFVJZFYHJGlHLx3de9Mq1BWOJxQG
Qo+D26b+EjVm76UUAdGKth4lzuDMzxq7elinQw801BzDxHiYVGwlyupgpnBQ/RlS
qsHR/39eAImcEP/xkZqh4ZbzsYfRh0D7pTZIboKEWMkfbAvv6Zr4PzsXn5malV1E
GzfI+6pLDf9BAZRpPoy2CjzbN1QqFTUEIcWBSErjifItvDmD4gma8CG/8sNAKZes
jzb5h8gSpQ73yU5PLPoK7zBuPnxx12On07vfDOBP2OY/FNwFbHjcxJF/2xtec66X
ENqTZlQG5lbRGNJfKMaVpPdwfBSEgGrWYB9Vr4AUUtNHsSyjbYJzCDdqbHYTnm+x
NxH/f5CuIjQjsHaF8p0fhp8XSTR5+pegoFd1r4ff1gBqtAT20Js/meAnzjKGxwXM
a6cUqBlZJSGeYWmomDSA44N1So4wIIuyRavd1Xx+jaipPI0lskBWFoEAvW4lQ0dR
3Xd/bBgwsyR/WZ4iuEySsG2st8pj2pr2Cky65oBmAJf/+0bXKcmAJapDdFkytL4W
Q+TkEUyUlZTn/Pdw+W11VrYsT1e9nT291OnRpdl7qdibJKfC3oyXXc3nRXgLksLs
VKy4/OlUewGQvnrAnVfqt9bobMbzakjJVjU8hN4v+nZwSIWpWKeSG131te6xIo6c
GQRbeA2l1GU7U7bSmAqbo6/Qxcn6JScelIJwAgdo8HCDNm3K4Pri0BnhGb2HMQfn
x5EJoPSHIT1fFpwcgVObOm0lbdF0VtswZu3j52dlwiwVnkMNdpQgcfY3eT68QF8o
Gzw2NcJXv/+utN09zJ0c+VXd4lP8Oe80Asr84vkb4Ltj0V1zPkP2dxQgPPQxSR4R
WYXglk2HtwZT8ebN8TLRSZbxIVer4uChClNcjxTN6P+oi7h6GUJsAdOaBjK7Icux
29Gk76W6uyez2ZAAY+03darmbQkLuPqVGXvH681Ugq1ODsDI2z4B4nk6SIX4a7no
cUTktckgs/ZakjHBclT9eb57OZNDiZBYG+UbRdrv77may9mvKSRL8eYii2olW5id
PwPDObduEEwXFt2oFrRv2oV5Dy8y4UxKKO2fNTycSgzY4mGxnnJq02fh5b+Hd5TI
j70lmnDwWKcVlQ5f1hbfyH3806gEE14XTYCuYP2T0zMYtFCPMIE+OwlUw9hZfj97
vln8qKf6OsZzdlEHOJ+/fOLu6IT1HD6bUf1B2u+ZW+5ibd0Ifz25QkqoH/HKHU4V
QqJan6daggOiIcUQulnxiHZRK3nCbqtpWsJ2FpyE9Xez74vTejCYYZ52pOW5Q7s+
I5lEKo8Nd8Kjsgfa7hUY48p2Os9GJyXmBCKVRsxpUKSYJLYZf6oaFIE7TIUC6gco
JsEZXX880z7XSQgWvUm2u8uoFn9V+czrkMAxLmzQQ3QQ0roYHucXSE61tfUZWGTz
EMtL9CWCG0Dz8FFxaitVObqsdLD+alO6dZjKCzNEsklMNIEUSDNH1WvQaX4F82tX
umGMxJdU4k/TsJK/AG6T3bH1ccMqoZnXS/A6iYIv4UIxJ1JBpndICflmcz9+XRy8
6bnCWoYA4pr8LTakmhSfAv2W+5RWA3FL2KxEd/9licZjfdJ1TXiLWUxIpSyRYLTh
RIHCoLcfloDYUhjUgZFqH9r2xQAQ/gX5gIFici/aH002Rg5d+4m+Br5Fs6JQiWk/
KQphsspUen5Ar6jwT1pAruA8ITxr+x2ebeRLwksUjahR8VulzJfu39pNDo9MI6j9
6C6oudLf2xr0ab8Js5rTqg6tR7EwuOj/qfIS2d8Fa0Ih1rygGvgnpln9ZDHP+DXo
wsi1/uoEx6EcnwRjTBAJHzx7HkdHiLBCSVcMotm2QjBCxTs+ZU9Qr0Cb5v0fj7TL
FsN8J6gWkY7FmJe5jRxDdQ==
`protect END_PROTECTED
