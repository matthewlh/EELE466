----------------------------------------------------------------------------------
--
-- Author(s):        David Keltgen
-- 					 	Matthew Handley
--
-- File:					interate.vhd
--
-- Create Date:      03/16/2015
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity INTERATE is 
	port(
		CLK				: in 	STD_LOGIC;
		INPUT_Y0			: in  STD_LOGIC_VECTOR(31 downto 0);
		OUTPUT_Y			: out STD_LOGIC_VECTOR(31 downto 0)
	);
	  
end entity;

architecture INTERATE_arch of INTERATE is

	begin

	
end architecture;