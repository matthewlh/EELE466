`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
bgyq9gorR/0vFmXAf8XY9Wc4SFEFUmhQ0Ga1Fs+9Xf0Bl579HemIGrvhVj2WOTHK
oUODXEUj8IpFUyPyeLxuD2hTom2erEe+e+uOjCrjxin9MB56KsMViucGpg9Fvk30
fVaHNZcmU3H2+xrs6PDiKEMeIP//9I2DRnNHY7BPDbppEQQXR+7asPvK1L2B19nw
BMlUqveSTp1Fuqszegtsm3kh6l0AqM+vsWTlOJ3Gikejado3j2irnWuT05MkVOcw
sU+49GbH4wjnK1B/d44CTZunPUXcmPNahbl233y1tfNH0N9FxPvEzpE0XAiXFtZo
lmpINVT3cwGxVeWCjtln+wwe9xY2n7wCbhrsMiS18x2+MRLvnE504/ihfRMX98Z3
+211nNAhRZZ0ODQBiT3C+PZm16vToV1m9zmifh2fatlPt4eCSD+SEl4r5PqI8obH
hCx5uEZFpsUyjm1sEapeIYQUJVRulPXJMoTiEVrnYCkHkCfVJ8zl9dGUrPvbuWY5
CTi7gSgwAeVkJPCYp4LT+GqE95/DTdn+zEbzhN677cUwd2+ORqHqillMwWsge+g6
dDMa7iuR1TKpfK4AZmHS/fQ7ABF6HyqRM2vayrqEU01VWZqECSFQJABZMOgyjM9q
rWsQd9eMmx0NaJ+8cR2irXYRmtREznRk4hCwrszzXqcOGOkztG4xJLwfF3LhMpdy
34EuUobEtFxgRQV0j4HvKq8U8CjFVXAFud3wQW7UwGYy8/FWYHv1k1NYb9CnIgDQ
S9feTkS2T5VBsS8pOtKnjBGGF5Kqf0ybNDUzplxkmVkgmsweED4wisDpi3ZvTYF2
nnG2jtItVuBB1E8zHwsBizerobb9c0kigvpAUSZxcdbZd4kb/Ak20Gj521TsKcoq
k0QS3px+uirYN7L5FdMh2WIyIFnKTQ8zFKe3cdudH3j7R9gpXZ6GOwa7LKmWi129
uVzp7JWeUt3cwCss3i/C/FkJNUgSNfbs1lx+Ue5emjbqkiwK4rp6dLMrOTr6s4aa
MzoMobbCyQhItQWqOPLMQO4BSh9gEihCvsyiGcTV7jrpTOLOAJlI5J1/rkSci0L3
`protect END_PROTECTED
