`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
dvZuPvrZl/hII3gyHjq2OmXYhNsd5iOwL57HnDWbmPNLYwMx+TNqRD+KX2XmEWgo
TUlYD+nR6PFwLjsv7jr9j1NCDxMy7dwcalhoMuR7riI2G2XLWNoQHCZKEOCKniMD
NEouGBeiWPGb/tTVtTLbfWELyZqSUEvrQ1kx5k4tRIkxtraBShkc3YJ+0EeHe78X
zXlhdTI6uyL2VBmJEbeBBGh3Jyz/eVDCzGTefKUB1LIjGPzTYCyoY+EpLj0Y1ga1
SzOSaZe0vg0UtsCZa/H0ATU5TC16UKDQ+VMvIIHxntai9b/zATcZUBPNGuKox4an
S5hzpymU5snE0aIc6n21z9nadguztySR0sjFza7NGttx06KyjtnrL0ltWfadDtsv
B31x+neu/UEmk0n4OtmLX6r4VJzc0W4asW3WTTkXb3iJG6PU2M5rdNvDoPBiqvZK
PJVW1RLWRg2FX4pvhDaVbQ==
`protect END_PROTECTED
