`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g+q13J6lip+G6q7gU6ltHmbKn/LD/41JtKs0z+vxYHveg4p1GxgnL3NVdXb/6TBQ
f0+l02Tj0xarp6RZX9B7KEa+7hiaZcD5SAOvjnFg06wFJJ8IhUVYqavT/kilXWdd
v23LDUseH38Q7s/K+XUp5Vt0XJ9Bf9sb7p9sf7AvB57c6+M48risNAOgLJcAByev
QOQVtvuAAnHqvsOUhWVma03QF24lXjyGyGxB/N4+xUaY269oDINmbG2kTw7rvXm4
cefUf7YHvdQsznLQWGGlDvg2ojJSuXXW8qjHpEpUrdD5ZF0jWvOV+lLUEGLigddJ
yHFBADbl8fhwuSleWI/PqUAhpAj/Qz9FL7DHmWivTmorqFKjyjgaHO875pBsEl+e
GDOXiuHRg8eWGGP8cyZww4Y0Oe6sMEyVlj4cYlq5o9OXrWGrz6Rofo/AHkw8AV8h
my2NFiQIkjeGhcXTghmAIW0f5BwsXj7lXPlK9rowHLW/yfLkGM9rSYEY+BdASE1R
gpdB9hlFwELVvh/oQoVLTHr+7ChW7/K8wk5D2j85Dg2psQg94QznbGAvxH5/qRos
OBLYHrx+5AAHxZFfbCoTwTCfWQhf4x6USpBsl/d4bwJKYuvbFLC3FQ3AzhuF3dW/
RUnjSVLM4+dMIKkKOq2XjFhpyTkIIedmp9XoJP+GebwLhU6hmpgI2MgRFODobyS1
8mJO5AtW6p1ALTAC3zPMAxNkjqt0L/ZPI4G7m71Sp6XToz2GKJioqUPbb/p6doSi
FN+rM8k+Z0iPCHFMIcd7ZX7MAXfM/Y1dtUPqVWesQnuIYuqkMmJiO0QQJYAFjXiE
Yl2qFJE8D3F0JLVcN1OfHvoVR6P+w6Rpel/z3XtWPEcvZnDLRPYY0CLsAVNq0dkZ
/ddE7Xd/G8g0kB8I3TlCfWBZveB2RDvBN7FKf64nH3HlcbP3ww3eSIvhYqMQFiTy
RTdla3GeNqYRYgm+JZIYJDsPmxYltzOEZXnnBgY1pucdMN5I/7aBMJaSLBF6fowI
K683TDCwHvsuRDNc1B/g9QDOYFyyvn631iopwT6Q8BKn6dkSRdM6FATFxP+UT4eZ
3zEeP2HUcDYMB6AF3hJ6N6NdcIywStlZgDQkRFvVM/YvjhI+fPRXWaiSBmoUJdd8
vmwJ1NIyfcL6XBqfcG9GPuCsdaFFF6svCl7VKjE2OjKYWCTh2XvoaIISexJkdVLg
WYurkoZ/hqyBKL65PpGoLyVf6sse2/Y35XQtSdcInhW5e4afmKxBzjGP1NSsn7oL
YtW+sMNN/FbUgzUn5vgms5ubQY30fSTkIr9lihWOCbFgg1kmxADFoLgG6LYyuNgf
pp88qb4XefCTdsz6PzzJE5AKjWrdVySSYavbQ0UpEI/BaTMg33oSqEnK7yehcXC5
7UdxzHF0ya0zc4OvAl2NTQJUDVtmMuI/+NQt71IzoyCCg4Ox5Q5mDkaA9C+lle/g
6zLGEbr8Qys9FNIKXNR8cwz9l0Ch+FZtsWaNzfsUVA1QTDhAbouCR0GN0WLGdHEk
0VHhicIkulmLuWnD5dTceDdjdTbC/v/uBk4J0vW5D5U2GMTUteW0UW3jkc6qcGSK
wPG48qKQg8iBqP8nr6iWe9tMQg072CMyx5VvjrRf8BsxIEoHNUebw/84PfmarlGP
1mBYs9t95HOxRSFD00mhbu2c1SpYtNjESRE+dhtPn2TlRvhoPK8jvHX5OVKe93Hr
mUSha0npQ99bcpaQOta8xffoYf9IV7goQwGpxpSbqlABov7D4KzKNjDuEWwbrRFy
Io9aJN444M8TKxRw9CnCZytQzymBHjaaDjjAoummWcJ52zqsK525h7ZzAgUBzUw/
o0dWYJlvnW8HevSvzsAb4MLj+Hvpttsm1toaflSQkBFmGAI1hwJLDtB8DEV74eRM
u/MILrOOSxeWGRjAjjosVfx2TGksMdYXDJeexCfd783vCGGABXBiiNNd4psWFV5I
a1q6oGxjxUlYUD5ZohPyvtAruVtSMByOZqHwbz0MNguh2G8V3EdFc54NpvWmsgCa
22YKCNhRGqhxZaN7UtB85kayDPx2BRwQMuAs1MIAr4vZTvtMibKW/MTdkRd2P2/I
as6RbkuCqrtJzbZ7X6ieeVME62hldcZvnEkwkb4CLsDfzBFMm3NxQXj3bjJwdxkb
9pFzdoiaTlO6dhUtIjpIrKBwo6ckh2m5Jsnu28eE31Z3NAzEkey39BD/fDyzHKIu
VEVlUYtJeNy6aq4FtHxXegsXZwGsBr14o1bATror+3KmwndXxkqSUqaUuKH5rrhG
r76RjJTodcakA3kPrn7jyR6M65raIbKyQAEqf04HDJKScxRX4fcEu3WCsQH/3ETX
aUDhFM0O/d40fdHvx2plyELkyhcpUiW/4MzUzCeq8DFntQHlMO5O8dHb5/Zk7EoR
oE91G2YLXHBVTnJlcDv6Fp7nlE+ELmB+hFpWPboXH748JiIkFp8PWCEO4lNBX1VD
7rYMy+JjwiU6p6AJdq1LbJUBtKgVQgsNfG+zcmQ/cLvo3QpVisY1K30mopuCEX1V
BVS/vEzHZ5s7ccB4i/Bj0+uOvdLopDNWB7BzWNTTIYu8r6QHYK5WQUVIzUok5CcQ
tIWW3ihCpUqxCsMTtUbdUtmnHuQ3ZHWJgYHlgDte6ssbdHRhvUra1W3UFW/GoaU2
XbY7kBZCpH6M3izYUnjeMudW27kjLs/eI1oABjujJx74tbeeraZv5IRVQsi6wmCc
9ZylNBqGrvS5nZHpi30RZmxTDNNsWOunfXaXHu1Ng1RczLFkwHmuZBYwPcPIGGk9
fh7lGNNsv3hJKlMZg+Oqh/EXYgAZ979msN9OmYZhy556XmhzojHOi1vfzX72M4sr
x/SVyo4jDkcRruu7m1lEwB3W9eG6hqZInlL0zvAh6tt5AYkd+tXwWNyVfq5MTI5/
d5ihMukUsiAPHcgzBTFhIiyfEUclb0EMM9nJzsoYQBb1/oQcYGkAwqclskLcVdZg
ekyStZXWmSOmk+JfLjJ7Nlr/iU5lPzyr0BrzapJfs18m7+NjFaYsQ7nuxui8mhPE
1rVKmU/AQuuu/eOS5j8gjrcOhB4lCKjl1ChLV08VCs9V9vllYPOtAnl47AmUBk65
N8gT0gS+I7/pM0TpEacI+NfRyFqogPR8s+XMfNd282wtc9SLomW5dzAmfXuyBC1R
AoNsjv1jKjUf4nWEiZLNd6OvYJlA4b/vgL6iVVSu24dESP+OEGWdPkxxhKOFOQYE
5kns4JQr6bPwzQ4HTErBrDeeqVQnZn2bBlRG2YaeNkG9X0X77GCMmgKH6J8/VwDz
ldw/3xbSplsvUNrzGNSmuYhpL4J1ons0WyrCHtUtShYP687y9PMslcOMJXIRuJyo
7SKt9/b3h4gj4jERtMy16TBp9LEKqLBnpNGrVHy3LFDZbMA4vIiq+gmLs3ZxgoZx
/Q1+yrxnEhY1qqpwCoI5cg89zEO6VdigxeVKdnDzt/JahnI0koe1iAjRQ1Zz5zcr
wBnMhasRCF5FYKoIdkskMCE5uJPRc/T2+nXtZg3oPLbyH8IUY/weRbcn1oaQ0gKv
8s8mf7GV9IriLz7ieqICtJArDDQ1EEEM7v6v/+gS1XQ5ogzXRPBV6HDUr81rV1Uz
ST+HFm8gS3ZNxTPVjC03xEbwOnD1JcmRPDPnqC6rnA9vaTOj6X8+3uJr2qnX7yFC
bzKfxsop45gFu8xpTC2pM1aDKij0dB4KUaJN/A+X2CxjQF1sqdE/d6ml0PtnPwNL
C6UHnVkfLAqLpo8ojRtK3c24f9S1vK0l4gN6X7dA2PUFLEfuSsa+E27lK/zKktrs
oEqm+3GyMFtlb+nVYDNt+uidGA9qjk8wTPb4fgvdShcnPOeOfiCSqy/ha7pnObfF
PqB1RchJk87/Wa0LkiqtxmBer54fe7mfiFbcAoI6/HguW//aIs7va7RBps3ypr6C
0W99YJHwRn1mcJfA3Uz5Z99vOTSkFDeNIjCqnsQHqvkmZoS/5nhkfPUKggFxhuu4
ITN/qFy0+kx1NavcTI0cm8xF7TlVA2YZvPmyu+Z8t8Fke/miQoI9xvd3XqTeAMhT
S3a5tbsWUv4uI4QzRVkg6HwpWgG4+ToFlJ6vPWP+kp6dt8zs98xWd0gEiyhS6teb
i+VbN5XXbIaF1fAnmd/IbxxaC6Luvw8wLlKniQqvgEYg/kAa8LA8zUW1mRzZ/YjV
UXu1MtExvqV9ZN81FpgLYhX5ziLxzLV59h2zpr1wnm6SbogfMKSkCM6JgVBlceOV
+YRavCyOzjHqbI40uiZ9X2oZJGZmZ+zSoqqeq/cO6dC1tWIbSp8D3PWR2ugnzWUt
FOJYumnUsNUHqRFSm7zvzgqm6iRVPupsaSJMGoRAA2aNp3i/8wMRZLlCcYZN0cM/
0MXELtKrtfc4LB35kblUOdqpKEILOHH2iW7PAw6hXOLw5YelMsFNPWSTFdYoCVmu
WJw710h1dvItmze5/1/6I2PpATQyvztfwwVQyc4jpDVlOHxK9T7OB2K0y4DpEuFm
9nyOa4WTsntsWCMpprgAKRWp8H0rc2ZiF0UOO1kTA9i/rNwbxxZ9QcT0waHLiq7K
YC/0KAd9xPzp4zDdBBRU5Ytm5j8CPZMJfYr2LX0ZoYuqv2657EROAxZB6u7bIToq
Hd0E6hS+5/f2qTJuInBVXEaXqvZEmbN/BU4oFTfdbkdhWKovL+1NJfyq8LOWMX6d
fjODw+b1Cdi/Fnp5+ouRFEsFvNnFwrTa00XUy4qq+Yf1XWRG5PaB0wppgvqX7Ags
kHdMtsDxfiE6pyZITYq3qTrGL/PEslMVSDylYljcij3SbGQvMhbeunzbOhLAu/A9
B4b6a2N6XWEMuC2QIaU79zHQHf+z2N3f9rDWQGj9YwagD3ZALJyKG8zbZybjmBs0
X5J3YJSL5nUqK4vV5PqXNfmofYPeQBboLLIb70Mt2IY0ObQpf0XYDslqz0bcUHWk
ogaXo2b8/U5GilNutKzqRg2LBnycJ33X2BXqZdEaHUIL9tWFrPEJwpM4ekmNWQ3q
CtI2/qxgcXWggQ5HaZ1xiA2becc6RkRcQCMQZB/+cBu7YWURbVdWb0lxdLGGYhyk
ScYhbRJviqlQhS9ckIanwzomZFQ3OhcYsDghGxdhqlk1MO5Ipl3Mwesx0gCQwEh8
xzPMJYKSz//bfk0MK3Avx8eJceK/Iayth0zJxSNUJ13LSm0seELznOQGDg4EVRx7
JD2AEaLSgJRi1M87PDYKCtMn0kFwrMmhpp/0BF46mGO8xPF8R7V+l5lxDzLXoIpO
kaBXJZalDV1TDMXPeTyxdJnbwejVekctZHLfSpjzu5p5RypFYCkLS61WgY1p4a1f
ITxZSFWYhBWYDxEiUybOEBRenenJVdfwIYaemBzT7OCPnPljIaG24P45/5l7db4q
8GPG42KpbXlRHzhoCkrXrwDlzupG6flkheLw+1Ey7j9j7NcbSz2ODE4IKaYnm6ft
kN2zZWn1Inzb92iTq/2hjJxbHlewjuTTLFUncxBRTT7QwXueRBCiQl3bTqKzjgq9
yk7bW8cAA4dn6M8q8h1e9sLEKLW3i77SFOaYRmiobcn+daAqR/FNRuz5ZujX+RIp
o1THn+QLBRczK3usVc/af0JgsDHUtWe2IZq0RFrdtszlkUFS7428WRWeEZBm22GF
byTdpMB0NQkV/U5t99SE3Y+IPq5YNRP5OhxXevpRWOiJcKotKSnJvYx95BM4SQKO
XJKLcS+uNbMav12uYafLkpva+3BSDJEvjDjU92sGG+1nC/rybr0i51z/dlJs1DEf
2DGKBjbd6g+s5gagaXnyGyAt/2DfKa5//2DMJDIDP9qre6sZKb6dx7gK0Q3efVsS
sOYz95xXixkWD8OdHP7RCz4jvBr58MLgkmnmhRm23M506h73zG1TzVyEbFRSrVbA
QtiIUNS82BU6CtaHSVu7Xylw4vzfUOMbHLudC4bEbZ6VQPV1EEG8r338MXKDSnpS
OOCF9fQQFnFr+as43KZdx9PS+SMDlcOh7F4/LQyiXvLSXJLHnb4Us+zxIJvgaJ3G
2ZjP5SYKfprO3jwY5vxB44AvXFnaOJ8TEvdEQAZmbWc+JUwr1RALAHWaL9rz7Ibe
d6djkJNpaIzbj5tcoqvZ1NO9RFxH/YU3yat9p3PEAXvRKOPbQtWhTFGVIq2+DEQD
qoof3rqgoXf97pl9d9H4FUzWDZbwXHBB+6bHkSw9DlkOpXw/WIGUTD8aBGcASVNZ
cmjXK6SP69ZL5qRj9NzD1yxBfgpmZ2lMJh3Dds5/rlhl70S28L5eowQpnFKHI2n8
gXTHHEWT/YylpX35KZrDm0LF9MAQyaw1MFPLwOvj5/FpK0q9JXa45nwBXVQ4oKpf
fJUXp3ijSES9GnwabfgvWftaaRx2eBl4YkNiTi6iyo215hjtjctaLIBDIP0Fi6vh
1y6TD/jPdLDj9fxbFrqiCNsWN74tM8BnhUysl4UB2+Vn9BKxSKUn+KOkXPMmf09J
Ogmxj8r7rMqgUKkf4+0OY/aqDjl6W6afcwRMt6lRzM7mjPV22YVSEiqA7H4jLl0S
WfRgs1HKte7+ElYIqOApbvgmAH3zTrtEYx/g1t8Qwxc4jziz4fv6IhmVwhhqRLGG
plpujfOlVBhyaRZOmReIjs0pCDoZ0LN4+BtIffWZyVSZ4HH/OlUM67QIhO1lqJ6e
frqyC5z81LyJzyKbQqS2AA1/k2095Zrf6WAzhuBvQPhGJz7Jqi16CxF1S6wR5aY+
c/4ULbv6Pq/UE5eZ0CuzdKYw0GZh/xETWGP9hi34VXEkBS8274dsQmptBqrYii2v
0jMVwHkok+cd4JBIebv9bqGCIZZGE0XNffmGgrrDc8ZlVTZqhGGUxKMCD9XDMF4X
iXKaXHsJord9TrQZOBGeSrrTI5Tt1zmsxXVjSv3TfDiPF2p+EcM0OnE5DibxWEV8
+IeytAutlOVij4wF+IdvpLd/JhBFTXnt/I1im60X+enQZHt6mrOZ1qbnJhGtLg0v
C/PR7FB5l1Y4UVT0JXkbhIPmwyw6KcLU0CB8JaAZY6nrp5mCgwLHVslf7t2vm5Ry
uyhCgUDn/LPiFXRVViN3ShfayT8fvSqWdqiYOmoFXu4ZS9NM3lmvFqSRQ9ZHXZhl
CSYcwZL8aJPTSMoxteWbUM3bIiybsaHsKTM2CARwmhrvSlsP/ll3V+oZgBJR0lSX
9MNcp0k5/0o5lEK36+WAewzRlrGrhnQEuZsjHtJdJCs4ZUA1DmtvsbC+ImelFb17
116MtQlszD5cQ9Nd0/7pCH6iaWir8JIb0pegYttmWN4kiNJ7e2WJtyClfC6nUJHj
CvxyBMYy/CjNosWjP7pEa0gV/jqAJJyWKtb2kSmVnLa09nypVQvrPY0u6jxjtdn8
9zMJlU8HPxtNmltZJCfwwz41ZOCAd6Wpbf/5g68WQOiqf9I+iH425ux6NvfUKYoz
a24LX+VA7+uWlICYsOS/DTlHIGG1qENeU5BVtRxWCeaatQsCMuxfrMUChnobK1YC
HlEyoXEqurRsWVLWE2nMGcyh4KwtIMenOjTriWBuWP12aTZ6yl+uPwyg9y/Z+WN8
qlp6JhKcBOuqnxbWwvf1Rj5bAKYJf0tK5u529wQrO3heAHx4fWck8mzEOXH6q06P
/vH0ZRhBRJ7BmJRmquk7+SL0Zmma/MT3j/9jAPeo9JGdFhTs5+HJfhKuSHSYjd9/
dzDK+lPWjzz9tKslilWfnGEbXnuSIilJdLinzhebRoYpoYRMjHPIoByH4bQ7A4E9
Spaha9PwOs1acMHOyuj1MiW92HDXywR6Q3c2KuYFYQPIKIpBDvbXo/fs4kk1TtKh
KmONiASAB3rPLOhfFTb43CuBV4IYaLiBh4jdY4GtJbD/eD4Qmgk/A8nJ0uLezs6c
cuANpAjhQ8syGP9HkGdo+ZtWXtiomLa9ePUFOebRGAQJtAAl4/xaN3YDXxvdI8af
kB3KpnauCbYpT7Wx0KERtgWyUs7pm7d2E2zb6BAQgb8/moOt4Y9IIwqVA1zIZlez
Lx8df8oIbOhd0mMZGRV22xLXqmDZwGV6DO8cbpldxvHRasREaDLSJx59TN7gjA32
DQuv7xDtttRItvroQnb5UgIu251rBvU23TLldT+/clWa9q60bM23s6IjVL8lZFKT
W9+q5K1pPaY8JRhTreZ4wRZRTSt8GJyLokLY8lq3Gzpo0NxVWOeS7nx1UQGezjSQ
2I0vQTystpI/Ib5m4dRJxe9Np7siFU0CQPIX95coCEAm06XWEeEcrLI0EQsOicWc
wWfJoWD/5TOlsVk9vNJmCWVp/QK7fkzNQvdzAjsx2IkoRKG3yEG9aUYcdul6bxja
1tdpgUpTX5Oxh8gY5chUSbBIIQwS2J+vVZpNhtLjNJrxglQ31r/cDgVIrDjsN2Oh
MgWcITwh6611rVN6HWRg15OjWvPtwZaKIlLUovWdt248qdmd8QpVgcJ2+zZlKlIb
yK5m7eqoCHIY9d9r7uQsvKWP/TQDhGRt4LKYmn/D4zpterljbVmTrvU2DAs3JW/D
C2BBgEcMcrwvjTE81qJCaK3zayeQIkh4VmjdwEKWufyGWnfnLmgKu51cZnlNVEku
UNwi725nAeNfC/1hDzQ7roFr6cCHjfOsLKb2WAVM3zHF7BnYKMfKp9TxfYCXtHFo
/Z8pNb6ooMQRZkYAiPrN5XTAEAqfK6ImVOIGwYp+7o4++8LBqv8bkFux2grPDsTA
CfTee3/q3h/kOcTPrc6la+6H58pnhjxGo1WdBrWI2HnvfgNdhZM6Av7Ao+gh1LNb
nbal+x/Q1WiPK9ouLO2os0yFRJfLRcT7fwriaoW8sQJlYDiz49MdUGtADwZEMy7Z
GZiXcvTawnblgXrCbVkCbXz5zRNjLKV3XdgQ4a7dUH6sLKctDJ4xiCEGxQftM95K
aWXuiOR/a942O6fKXKPY2nPvdMEkqzyzQJKdtOenwKAo3zp2mdpxtrLJCfNzUPAf
F9GCcK+pVa3W/TgSuuypVO56MDeyW/MKz5k+y8YGana8fGqfQUU1Qa6j1heN+znK
d3XVsijQhfzj2jm41f8M44sC6ft5wqTo/s8FR1dT4CdT5/UI3HqstDvdasoAc4be
sa8duHrWJA37CPNK6XF+Ua82+rDWo4iRRX2AZ5dNd2qox3P3ftDWqJd31ubGRz4T
0lyaHCNiLf4nLRmKaktu+pA9YfG7Wf32XIx1WJyFcQMIAVS1yZ+QTm4DsS1FNddu
/OvEGsWuLw1GfNGXbzMvfVLSjqMnATtDGCC99T9dK3AgXakyu6q0mHey3qw4PYhr
fwHuz2A2SxMB7gIrxIcOd4XQ8bGcZK+63aWWP0wlnNXy+WOAXmfmy605Oyi/XFu1
G6VqIDcieSazo9OhKQAUnKW42EoTy7DDq7jBZinWZdR/sgSTYASiiKpq2+xToukA
NGjCa+L/EB6spbSZNJDiBUOJ0jeEcCKAscEIh5DlC2CkR5hfOf9t8gu3EqwEKKig
Uho1fNY9Y2dAXZFlMvMG8zEZDtsShlNnC5hdWUeZ8wl6W+kwme00YRb4PtOKXzr7
10XpN+3gLAxl3G8Y8tMStN8UpgilmGmrp8majkgZqaY6CCs5cfc4FxU4daS2g3MS
rCdlZ/BgHaZ2e+o0tKerpPZNv6q7uCM81vtJzVXk83rLwWJlEdAwdugAYtMMzEZa
hQ6C3IY+X8uBaE9DbVQHvkrdFIDFkjgPimrxhrkjk3dczdkt0lZy0nnKtON2gfNc
g5znKHq0ADTcq95b16C6dOf1cc5+sL7cINkx5VaJfygBkoM2PoKEKI/TVQYv7tog
+miw4+8Xr4KF7l3+NhCOtjhi0+XG5aKgNkl8TsEOFDECoV+btdYyVr9NB3bAXqpj
G4IMrvqsd2t+rB1pzO6awhcUEhNxbl578P4ucrWM8dt4QorD3K4kdHbMs/AEn6/N
mQnKasb1v+jWjO+f0oLPsvseB7jBBgDiHLrVz8nmEoHvdQcleLafTR3y2vUITIi4
dNNrQ4CY33axcESRyn/59fOkUn5Yd9YrCJs4aa7Bmad1Kl6nVS2/0E+0D5YPx9ys
0WIv4K05q6aRPFluPDTso2/4dQ4tD9I1vYtaNue61UPQd2O5M30Vx2ckDnvIdnbE
1LuXLvG7E9OfOxJsTuMVs2gq00mM98RUowzYFd9x038GDY5vW/W7ooKl7bKn/XEH
uIKp4l1i69D6zA2NPHKitMqI5NoUt6ogdSSYGhg6BX5AK7JwdtLQVnE5Y+t8Yxhx
RN5Gr6s73VbkmDttqDvKuQW9wxxWSaPyVYHjey8kUW0Hv1O1wAQ+cKP1Jc1cSpO6
xYQyQtIVbCLqMJV5LkJB63DE56lsX7VpBfXFHLD1QWXs4b7XTn6qKUvostqmj0eR
qWrmtykoXPLzqUte6MpMbmYTse8agjHKChIUUfZq5UZUc71MPDJCMwCRwbGRFlex
yeEQTFZh4L5lXLkDWGIP+3+4haweIr+R+6AULasSWSC5eJ7pD7CEs4mMHTt84JpH
XR79Rl7BRi8lCHbtxhBdAq1hW+lB97NcmQicHXw4w+SSP7wCn6nG0906ZX/5ak44
VLoQpJn9gdtl2hkR/1sNyWrjv7kHKnEr4K/ay0+iwGBeApAKSQ6WPjpx6YCqwUAs
9paF32MKI225qj07IGV0DiOtH2DFR0/Ok1DummLloKVQEM5aVH7zXJjOVqCMKeRI
XUUPEh4fbE7wKK1Pxme3URrEWEt9c0HvBK0Yrtvc5KMgxkfg52WpVz9Xr2Ukvf5W
IzJRkhWzxtYjLNIMon8YlFRE9GErTw+InAWIElUyoHE5aYDOyfArreE8XCg85Fwj
xSSJPt37AGzXOomGxYG83tW+vxOJThkHxQN9PskHzr+DTSv/RM+8hI1agrwD4xWx
vTPUTOJEyw31Nm/f4jH/SKcKLKVJAWIYCt3s00U+4r9B8Tu4sXqoa9krrK5Pe8cJ
OP3O8Sx5SOkFumyG1+o5GWlyIRrOhzeTpYK/XjQFN33WnTOv8m/T5nAsvVj7ff8+
jVaUjcW+gKmC7wOditUranqONkaFeyBLOl1BMiL7niPOsoh2K5/8SVXe6Loxz/Ag
GQThb4eUKFUGOBqA48hphcQBO7ka/1ZxnusFMsOXwZ3R6wm/vLmnsVbIMgndYFku
EgA4fLNnBmhkilbBaJPuGDkyShI/wsVhfk7C73y4Xp/529zldkF5xnxozuE3Lo5R
E/GObgkMncoGiMekbISLELuqCRg6b5So4jL4WVIPMlY/lbjsRkxrTBxMwAtCqICx
RZntVvteA3YxylCtPCNC402e2t2kYU4yqqAc7EjmLarYCeA5pb6zO929qHM2lGoX
8FizxH0+n+0u+vZ52yWH14pdgSZag5YT0bgcfs730Rm+Tq8nYi2cDTczGTbqpfbp
jFC3hA7cCiSTtM7D9Ci3KAj8dknciYWT/N/SZODIt2OglaVPKuuR2BvvYpe2AEaw
0B2ZGYHXW+FBdk6pQl+8qrSK8n8xk6qFLebj22LR/ploXXnc53nsMKNJQPfxkrz+
Don14WH05RDc4ZR3dEPeuXf/93mP46dJ4l17/eRVW1rNggVk5pOb4Eqvu5AI8iRR
RWsX6k5yLhUPBzlyVaSkVjhpp8ZAyfWeT6KTWyoUkU/piJKsUjgpaLUXgeR/AX5x
4SreW9nEQwOG4LTSvDDabr+m0+cY+CGsrD10mkkpig0gSY8JYCTQ4g8cWDvHdWWk
lr2zQi14uiJ71E4bo4p9N4pTuc9aYchsoGcdtYhocTRDFFt4vTyT6J1WWDOIr4CO
+4BMty66oiln30ZGfkKhXtqEeYtqC6gqhURCszRgf17S51GJVdAM6nhzlaOMI+yy
NWDcoIqi3qIQ0/NkJRWe+ofmE3MIlEMCOMgm6LePkx1RqS4pV5zE9M+kTjpBF+4o
9IL2D16sZ2e79O0ET+ZzoS8zs91RLpx9Qov2zj6q1JnR7TzlITRdGrZPy8uKWKf4
xiN2ryYFzZMbQAn2Z/cGL1cypmTb+0smI8bG1wwZNq3ezF+CnnWcqw6+2dhp1MG5
rYvvbiCiwFYticqL7iCS5XRWoy1tgiBklI+kUyHZqzrH7HyedGMO0AVekFzR5bgO
NcpniDZcnPS7PmPCgiJKyuuo25zbiznxUNrJgK/nGsj1jchSfJ3wIEk8rM+WiChr
UG7mlJcQ7ouhpv5eA9aZy/cj8YugrJi2fblhxYDD9kQYosZbcpO2/4HE67574B19
fYHw9zx5guCrE1BFRPYo7vMlnK5CtPGIsqKQiX2TIGrhkZmqFrZJRGzcierOTdak
cNekJozbnbheD7C8NSqihobldyMv8m/OTJY/aEd1puqcgaoGbd2m6tig5/Fa1i1Q
J5iA5tDLJzv99dtmx/P8YLluV6yIqlGp6fWPbV2OhD0meFtM09L8AQpJILAF5h6X
v3zBqW7sYy2/HB5KCmZoMJEwFs5vKn8QNSKdwvqlkzslzlKrEj7jxAPBFEavVr64
ObaD0OoJiCdwOnLI2vxnC1g9VwqHUJGnkp4U5AIG3zO29oAuFHw8Dt0U6FADXuFc
RYRI5jyX8FbC/ru9Xt+HJOzmazHyZY+gMDxMe3Tc00PjK25xV+AZALQJ4Jtc0Xlp
/8XZaZbeWwwYU5YpdqmBJy7PtLXhNaP2VHCHERKU+c6rlmACJPA1UzPvLgMgjvYX
/QTc7r/WhzhmLgkGDmmjZ5Vp2HlJae1EfTL/pi/a5M4m2EYRITa6uG38+8+pOrn9
Okb50HuLlJ9ofAInuk4hS2Rct0tZxHNZyjv/j2NGhmONVNZMO/RBYujTd3m8HeOG
BTeaI1BMcfq1bG6HDVZHl9lyBYxwh9Y5iIZp/FORVK2llJgBXuj2Wo1HLkGYTqLJ
qNqFoETKpbt3jV9XZ8hP4Q5roDcHLn+7pElRdLa9Us1IxP2QvGNE6apNeltmIP/a
re9M4WPJVmpX58trbbcs2WE7oLn7+o9xTCXliPzRZ3cxYvO80ZNfq1MVm3pBz5OE
O1tQHJHhXBhrEet7SYMGPk20fbMPM3vuyIMy2OKvKzzbOObSVB2SsEh0oHE+BlAM
N8DUtgXtMGFbxb9TCL4/ryQdmc9rdbof1OHUKylwWwjSLXQw9MrM0oF4JS/jjzIZ
5aUdpZJYXiVGo+5kpsJlvzlLFljdrwoIHWXDFyqVPE/So4YGNOGl+HpqgApaxXBA
CrahNquPadR80qS58KZNgKfzFNUWjtYsRh9hRoJbUZsGNrCwkpKamS4wJ3FuY7Ej
ejVTtrybeBp5VZ2jAcPeCuZ/GDH/FSGccbQwDoQaZSEVh/sC4r6gekoMmtLHam30
Pyxv6L+gf+H+HiEoMe4ILsuHgLVreZziTPDQk4ci1jlbQ97SK/YRFkk0j076gEy2
fhGLyTpxwvRHKqRtbiL0DcTHN7VyW3qPD8NsbhhUsk4PXQ+GblTQLzwG6iuWjqJF
Tf0jDufDK0LGBwuxI3pP86RHumoXrbM4oY9ov1Gpn+kDansDBJZ6CO+Fn7hbVM00
VwrKL7lhw/3rXHOr7PUAZysfP+GCQZev8Tr96G62JZ2rR8Ae19fRBpDq+93GppaR
Irlxk1YQ3AbIgT3NyJ2jATqEN64njUKMwOuoYOsd4Ec3hl6TR5ZVAjMMhPL8oe3j
DRGOGcICnhjXLswJ8HEcysu07mDNS8nRMzNxGgdDLwNu7n2swRVcCGIeNP9U0SQF
fhTlKqqdNjMM1zRi262yZkpDDOkXatTLwaRwm86P3goCAGyb5sOCl5N//F42/1CB
ixcOQ24tZTgYidTD9W48V/t9LL7YxvkgFtHern7PfEA+8uvu0d9dB1oFJjp+v9cK
XTxN039mFVL6On3U6Hx9QewE79p1nHLj8eapncAaTZFwggjQZYoMO9VTgcmY4mb/
Qkf+45vTuMVny/W3u487FvGGYfFuerT+hlxWiY/sTkbfTD5Zw/u783yHSqkuHVJI
T9D2x7U98vEVJhTGaEV+p9PRnAiUOoDKQDeVdoKckcSAS1yNDuloFaCaKW4JjXUd
M9+TRajkgk3tENegl8XYs43/uQ+P3X7w7jO3F0Cystm7xFryMeD+LhMqTxS9wR+V
lEdP9L5rC8gecPksRQ71+S17tJxUMGdbetjyeb8pmP80DhAL3el+pxgtJfk8JP4K
7vu0WwPVvXRBOf4nLVdigxwDHloWX80kHFw1qWRTU/IxAtNnxgCethy42wDGNiM9
vYqMOQrJU8vbiiZ42uTQKc4KuFwEl0/EN/pL+LNiOu8nt5kFX6YV5E79RiohTw07
zmISEUFTReL2EjwXA3DQIyLFj8g+JBorRd3P1FFB4q82iGuXGRyD5Tj1x923L/X6
mdfPwyM+D4xWILX92oxvmT6E7JNtIV8rafR2B+hHZG1uc2xn5BmdnIPrzWBmGl8H
e3Dd1SkTuRP6XMibJg4slBn+CA1ufXr1JBQSojDLk59wJyjzWiFmtK5A3/OE60Jd
bWlxVaWNrGigYm3kb66birhX+yvOiL/nb2tzjvsIR7dUl7qGb6HrDs9kner7DGvw
gW09z0ZzUPfhp70jdJHAezCVyiXQI8/nXlFVxO1IahgheFH6TvPoDbeLG9TwIviq
1Ur7u6me/AkM8R+7TAJVs30aGUiNxYq2Won0C8ti1zLMLqH5L0n35zl7bj/AQMoF
V7cjsBbMzypUfXzhwQo912JSk0J+8jX8dV/+2lwAioXmQ9cVGcD9MuA36mR+81Pf
zs52A4aZAxxaiu8MPqt+oGZZvwz4YysLQh4iG0/VtgUJhUssTSvr6IbBNiF9o75X
LsDRx+ywy26KwzvpaVSVdFu5TLqdxJ0xufAK3cXePQ8ew1zDLdaKMCIkz4FSwtna
eyc/u8/S7ipQdM4g7vxKpL7NEGsM2h5Dl5RPoxZ6zvt3P87g9rm0wehV3vi1OKB6
eWrfaaVR0oNgjjMOOgXzNVeOHyjKCh2cQgCvnGPeNA4n98Jwt/jiGvH2O7mkuHd+
YBi1bP38lBaRDhrfReg7ED25djrGTGBq7EsJ6dHuu1SX2shsATdltAVJHveqVzIu
IWipWsuqNLSee1V481glwNnmqLPalpKnGlpbIBH9pTEIzVHKHv8yBeQrYQ4VqqD5
GsXRVm5As6FvVOkfYo4N0/IU6bwIAsrBU8l9+PZWBg+KgRO0n1QbFllOCapKq5Dx
YDXdchUM2MvlDnhQIHh/vAM+cyuTSwyN0jR3p60mcL+Q+TNmisPZXhQMEjeaN1XK
Buh2TYjEdDn+GqYAtlt6juWgRjdlAcHzWBMH1dmhfx/FPAGvZJa+c9Gjm+Fhw9vI
hrQl+rNnMWTPiNr+06wH4L22cU6huriRKD+S2HMCqi5GXvuDtiEHaDiV+1X96Cyz
61LGuYMj4XkGSl0+f/l+1WBSKqcbS3RD9TCDWFVhA7yGXBt1ZmMGkvpxYH6MJ3vT
UPkCSl9V9B4nKK3hmIKv7auvQTrRl0aMlKO7AM+IRs71+zAK/sbuVT56BAi+YDVw
2j+tjm9WfVHOIg9Yr8fmS/yQwY4Ch+Q4zeMpYdGf1yRfM6aMvyA94yAcrKj8aolv
ewJBk5uQxe+Sj1NHNOmFvq7cImiL7uS3rCVDKW5U/apUotvAOChhMLWo6qmRcmt2
faBCvUhhVfK+CtrO86y6aE6vNV/9q/vpYrCyyT35ik36QWZlP5rPDiKxbose3CYh
6DJrbYKUjinMZjBkpahP84ypJE9AkuYsOZySTcC7gajrshGtFL3Tsr8tk+n8OjfG
mQMm6vIW+WPkCA8EYU25NgB2Fqn8rsFXc+YFBr3bgG6FfXnNUH7GKt7eKdad1uoj
wY+BrnrQUaoLC32/sRrhcZGlXzhufu6yErTvGo8t2YBXJtCTtUxzxNzTiqvCvR+G
hCE2ZkmMFif5AUS6yqVIha+VlG6886XiIOvMFjFEy8jKDGUy529/oP1Qocv4pMVF
RM6kclX3/7lf13Zg4v4dNuCDH+i3qZ7uHYSDyFVKkt9BJbTDtI403edE94wVph6D
cnDqliUzfBd5bifFPaD0yTxVEUgPQI6Z6rgEwJMiSN4o3LvetA/l6dULcbyw29DT
edv/tCIzJfZvgK0w7n22T2ILb2hFiuZH+3SZu+O47W8Fvik4d1SGgM8KHZwWYQgL
aZTphyDBqmJKl0kONF8Vg0eNWCQRy9UXviSNxXIPyOREDDBI9lmbDIGR3H1isqgH
APXqA/aUVjBN/ORPnwf3dsevAEU47zKEGS6L9L3GpuBRClj+PzRPFn33KMfRl2L2
q12Lxic3Xb/msZb4Os8utnmgA65c3FWgePM1AmiDLte7CLI0lU9UsjkHDdhHsxH8
/uHYAPB1Zv7QdDQd8Lf9amHbRaE0f6zj84xMoDJglm6Xs+9Y66mgUW8cVGanoEr5
S0IK5ggJzwVtybmqUOn3SHDpMAqV/Z3b8DRizSjBPGbBqe5DH7NOXg5/nEWnEsPY
4pjAt8HeHXdU+pmiN/4kGgBR+c1+12+xfXq4FcvNaArvrUIegWUlFo1b0n2PLIEb
fIoJ2B/594LpFTUMDmCIyWGPbFTJPKLSkamwh+VmfmRSMTMLwhPyL6n/gL6RCn/9
vZ4SL4hDyJI6sy83p7lvbcE5YGBS7MOq4mfhmnzKEcNFX+nzThepcUq4sNUzN0zN
Ztn6uvjtHeGzwst0yVwCa7ZUBf++zJA99r8E92GmNzD6r+drUX7XIzP3Gf0ka0ld
sb3/xjSprmlIN5N3ycqn+LfA6ezfvTnjfLB7qdwNR/xFLbmkr5Mo+iJimta8hZ0S
ukyhCcmgc1paQK0fgFsff+RlNfUJRtnzn3uET/GE4ULduh9PqQzw9g1rB/qx5+gs
eEw33SbhQcUe7/LUQ+xCKgXRuqGQFWagN1rw38KGDEyvH+Rvo+XxCgsTe31MnqLZ
GNtt2pmIZFWcEShNfU2XTUW7e5HQooo+F9v/kizTi+DCwKC1I5bn9uFYSLujPdtS
nxMcAa1VcBjYTJziCGGf3cMOhOfgWRvRjY26kig5/5tizZAz/Y8A56jIOC8aqvzD
OLbUnH6UozlC1LGxJRScI29y+YquPPKQQVtBFKAxNleXoxVopy8ES11cUlM3GuEo
340VjPskmw0G6eNIPXtUcSaaZiBS93hj5saGH9gD4oIAwmToyp/SDX9HKZgzliLT
+Kg+J25qBR9MGqyFN5/NYQxjRZSqNhc4Q27tEceAOdVoxGZcA8e0h4vQrET4FY4i
HefLGB78VxPlDGhuenTcKmT6QEXv/cAKq2qETiAZadwXN4wiCZMjcfoZhkZBHnjM
gs9kIbWnq1oHUn10pzjxjBjcG8VyCF72T9QUtP5oJeY6i5O5+rV6UL8SUrRSjjmg
XEOSJvdQHhEFgKFYqCVjEfEcvLDDJt0Tdd/WU0nI+tSh09qTINeHjEONtkelMdaq
1aKxEX+fNso+HQBPfNln55yBb3ylagvvpoiOe1SRkwG7zlyWs/FwZGxLqAfba8gs
Gj++AspbjBMLdjUTrTkGyNs1ExOSSrb1NFZNWlP7SoDUhXsiq75VPvMK38FD/CAq
/0NpsEQuspOaQ0tUtwRz4HprP9VugWZnY5T58d1y4HN1ytLXPgFk9ZYeAceC43ao
x9TuQ11xwMb787g3m4WV5FIECyOLA2a3+loRu+PHE2iXHSqYDsJwbAWGW+luJrbK
+KmkltWKBv5r+mX/RZYwNpfasaeLkNjYELZSESE6r1A80nL/QXAMka0GY15AtoXT
yu/WerAa9JbDG8L3xxVyNVLcsog1ZZCNXyjARi6d70pKLOost677NkKSinPccq4/
HTGwPYRr2WlBKjemR9ofg9rmsQKaerHxuK/b7WzdSsC0UUNK+CGXbF+7azmFFhLr
F2ZXod0A2uxRckE+6FXiXmGoWgjJ0evUrx0zxGRh6heHZoWbeQU+0BBGyQ9Fl0w9
8nybp/Fao0scVao5cilD0qIT7BxLvvXUsjOqDEEkOe+l94SaB1DANqRtnRD2JpyD
Ab3hAwnUIjeB6wwp0dGlxHn9iHHiCwJ5vwaXI3nkqC2FXWCciSH5hUMwM6FB+mbL
FB9h5vlHbiMVYQmtVnEEDFzomTDjQkClPaZoA1ueL1pxF6Al4oEosxEvnCj6ftFp
qfntyIavLbmQP3cPZT/1xLwB1gbXge1J2DmsHR/nfECJ2v6H7lqOjoyTBrIXpRSl
1shqSXiPm/pfmUVs28QBqr4dWGR2U2baeq5NeBcQYi2E4fDX8gvwXE6qtU6M4bM1
eWdrSmu774rBhvYkXR1gTLdd13KkEka5HdrNO39fMa6SqocdwA/qb7gy07CfHkzm
zbhyjUT9Wan4sAmWwijikv5sM1xoH9TA+8INuyyzHyEKyUPDgNKLZ7j6zXliuaC3
uSIQBkot3kiV4MdAD8kpWWjGzpQmzo0yfyyUlwfQ7Azpkt5tdmMloo0vmJ3Y8J3T
Ubo1IxcbaTgrNgmD3AdR2yVapoSGe4YuJ2MEpewuyFTnwOJBab1JHMufXYfpr/ah
9zpiBQqfQAwuJ+bMFSg/s6/HGiOiWV1pBn0242kEkzfxl5tuTMS3cNgZCJm5RPF1
C3zKt2rudsyHb97f8tXA2HcSCVj1Vx/qAKzCf97akwnpeoSkdZl5/xs+wCjwAhx+
ToqQREadNgSPp7+jyJlZGnI9LQEDf2K8AJ/EQIRgrOUA9+gXttTPXmnYOGqAKyRM
BxM1JYRuUuD3uvlhjwBr3MMP5TLAAWK/0TZsnoTJx9vHRF/Bio62GSptwI8unHpW
0jqvbzfsoZohPxUlTUw5pTkE2+GxeCR1Fy3y26qwr9e0lj/2kxntAK1GWI37Bh1O
zFhNKLFhPADz0Hq9IVj0atKBooPlG/WumG2MYjXyDlJGvvbVtTijS3agsCVMdfuu
oJ/DxBYu2UPh6izywgG1yvaxwuFM/52W2CVpVNnypQleHGxbCemzQtdXDhrH/Lsl
fIPYQGB/Pe/duHvVXNMzpWMBz4XnbzI0UP451HnjCnnlaIqU/9mSNtK2qfi6x0bG
lLefQeSo2t5y7PqnDlhU1XocumxkFoao2D7Vy1w8SHbcqXWk6glPkF9sWXsiC5cJ
SlBVH3XvBuleDkWHW0BXZZQBjQfq+4gAaYygJTzziwuvKix1HGtMwQ+EQuY1bZdc
nX9W+jhk0DffTExIRZn7Rqf3N+G4SRmR3nuigYo1OjyRvRURR+u/oR6bTgatgIX1
R4/ZwNtr5BsvtuRLUeujyikvLSwhVGxYUrDL0GhEwvK2soZNRBwqTWs4BshAqqhg
sV5OkbjMw7htqX5a91Dgms+7wb0G0XKprfJRZBMugo1FYwVZbv02laksJZq/qIq9
92Wo6W1Xe+1U1oruAvs6NtQB0X5hIc0gtJ2z/l2A8j7YJzH0JkTSa52t8v9Zw2fG
3wK4eh1CSyMWI73uO7X091K1r9yL4UHxNnTGInTt3GpHDtCExHC++yyn+/utRp1b
y853Lh+jGlpzfQtRFWsdo8OqqJY63UgXgJ+nuoULl0kJDJSmo97l1fQrLBu+8ohU
hLRZ52/uj7mLy/nP+Gn1Tk9hNwKiSfiHNjTkDQyHPrYiwSAUjoYpK3GOVwXb5euJ
chE/A9J+W3d6ScTlW4GdfQoAgq96azeC2bNtm1Zl5yFbzrg0TpamancdBFD4jHqN
GRMbj58cwE85hZgE8L77xMC7HTcAjx1+1O2DMXN7XvBT9TcHf2GVxiVIkB5FR6w+
ck0GWZNo+LG2jA2YctNHvbiwHZDNfCKSiTnHjbnKCntIGxFR5EN3Oi0KWCWlv5+r
yvkKO1B9Ci+6YxV0wFAyjELkWX5a+TuLTL9NP9VWQu2LRWSCmYX3a5Y1rwKOAq0l
YsL/0yKJwc2Yjmn9cqq/foLc5TXvLNhzWnFJ7qokWTewEDJOStPVoJBj/n7DJUw1
sPUWAqztK1FX9n6+sLE3+ezSCOZV1j3orcMZ0Wz7enO0lyckG/yHKNLj6J8dyxvS
qRuGWHdzyVYc6cj91JcUDI/mTsgk+hmfmHrzrMzq4dg+DQqxZM+znhIjIr8pjkS5
/3FNqmaPPXOyNzWS30OMmnxf3BRvBozdFPdgNuYni+uCqqBbdejuu7aDEWg25Ega
Ofq3B7e2Q39VE1CCtaHd9J8M9cDJikT6kNBboSTd9+gdQl2lDcNRWhTrNf+WHl24
gN3RMLgZK8UKWADCtJrFdAwWmcRXvfi22hSlBpsmFAziU99RnpWP+NzzV4u5Fzp9
GCvNGZ3psqzN1lgfscHgDBr/fekPsWGrTyyzeGYQTXxa+Zlxt9mx0Z5jFtG0Zo4K
6ZWoo8HZ4ckAbp+R32JJqn7MKAtiQd07UyChNP3P4BgNgSia+SdG4JFOJcHmjBIC
yZbLYwyV3VoY0WE3mqBPAfP47QpGrykf68IJRFfof0ORBtavPo6K/UyJE0fPT+hD
7gZbsli4iTRrX4dQWgDqSmxlV0ff3S/LinPXY3cOoaoELzHDamGCEaE6tmVtmISm
M9YZTNzwf6XhEBx5UTN1YILmx642iT/0d1cE+oboyeye+8HapkyIxrnmNPWei9X9
aaTMljvtdzsea1ZMgLArFk8O6mHFW/+66c7nsCDut/gvfHabrNkMwupM37b7Xi+K
u2OYvexQx6CIHWbA5vZbrUYGem0jXd2SCWQvZQjLi7723kS2OtH1QF2MsQI117EU
E+TTDpFtkLA4k6IUZqNYQHdjR7r0snmDomZoa+FUcpfopQmPdM/tJAEPxm/W9KN7
YggVTOnykHb3/qzpIqY+47USbJfP0OCADg1z/tg0xIgk8lsZH89daruktlr+upT7
fcKzMtkdq34xBv/yA/cCjSjkYu5k6MhcyP6XvhPAP9q9jz0J8+x774/rPHixheSa
10LEBh+3Wldkb2WJhHGVc5SoZoiBowdoCNc8hP5bdfhrOZ8SZmfhZ8ffaSUkj3eG
prJZ4pj1bWv5BrxAxKnUewiIQLQDLGQ1nSFbzzu0JTwak3pPQYUeJDE06gbmB4KO
dD6hZmg4KLK2CcoOVhVLIQJKQNE+9P/xcK9GtVVDSWugFfErEcVAOD5kxfaDcQZc
38F98alpFCU3LV2P25rC8Jt8wJabhg5tEMfLXTUfBF26tHNllTmTgIWIKZwY0ImC
Yf6MMZwK8Yn/nxIoFCWzE/g+MFvj9vTY4wVLD2Amx6XF957Y1uJb2ng7OUawcRRM
B1dWPSl2eEHAsy4/0+z5toYI4gL0DrG6UOjbfCQIh2lv6ZH+Qf7t9lnrNdJPAbXz
hvnZhWgNN9HXojNzDgRkwrmR3Hoj+tPghqwH/w2/kdoV/DyABaTUB4JOCNQaZq8M
1SZrC0NsckF83KUMzaAmZsa9Wahqun8+sP/Lhay2L/+qwzVhMMijf3F+FT8Q6e2b
Vj0q1ZeWPep1ZKxO5ko8Sv3EIArsiphW+5r4rNlDaoVLu6q3eTviglgJRRcGGr8q
E3v37qevdJrDGl840u6aRwtLpP4YBp43wkhBdPa0l70Byx4O+t2QlpNtk37O3xJR
JMZVAPfJD4OSNzAhcxJNbitq+NUT3zJmXNjM9IkYV9fPramz+3e1EHX2x39hJa3n
t+OlAJ75XoiqWiNwzHAVsf0fTpyDkyQ4PZAXctYecbM84HW+rpzbZfYF5KoNj7HF
ppDZhxUx6u+2adwZZqBOPtD94MJz95DbnCA1L8CkjDSFyIEXEv7VmiUy7ejtjdmS
fnlAh80hBZ8aS7evQuGmkYme+tFlEUbAApVydBP2u+EpSUiOKb+I8wmG5tyMZkIl
zGNm2bSId4TONt26V9Qb6g8gelogjZR/DBheFijqI7XgEzmv91j84eI9ZG2ORPtD
LxLa6YuXd/ekBpJvaZxtJhY7e5CE5lsU89OG9xHxStVMRa1/HE1wuN3WXqCCCqYM
n6y+u3xGe6yHq2gsg+Mc7q3u/gbP2PYFKR5vvb7z61Q6aq3D4mEU+m1w8tEpoYDw
ETExJVbLqfieDdWGwqW+8l0eFOUQvDx0Wt31c0xS20qhTWCp8KUW8jPYE3O25ZdY
AAvPyDWinH4KYKZiq+H328HZ7i9VTRL0TZVxZ12tuuOTmvldoVqrULl7TcjH7chU
VbyGT9KjK61JQzuPBR8/04Zqd60EY1KG8ySM9Lmz+BG4ZxW+kn1f8rw0KTJaXeEj
1+YZvQivgW1Er55ZoW23YRZGdb7aBC6W/mqFkan3F/JaBvsUXlNJbMkcGDlZMDUY
I/9K72ToBociCnuzje0pgSqGSaJTXsW4cSwOvURDi+0c8NQsjpFsis95K7ahLNW+
YsADsBDT4jNgUqPMRsIgTX2DiKbzfFpH6dykj0wvYRCyptDnRoa6ldjRFAh1s+lQ
PulbU4324o3vEsd99A6SRuKQBWCTAS6L//DV6waggZEKDPGHOqNw9MhdQzuX7qqY
1LjVOa5m3cbiymxDmwkcO9nwBdQIwrghpgFFCT09nI5exMAhbDptPeHIN5VP4Pno
/seIu3AxdTvk2cVt9rDvRR58d4lrotSCXfP7AZ0tXHJesFaT4k3UnE3DayUzewSG
DE2ONmr0kQ4kHZ6HhUds39VbJ97EURGwJuNnZLHkaSrCM8znWp5KsBulLwFGJD/J
yXcvWy2lw8GMjKgWH8LlCYZHxcnkb378JVzBG3j3Ket3Yi7recp8YMqiWO0yTsg3
aWLxP40ADmAyy5161ZVyMQ/CVgysvv8U75wydlgEXbP5UsfzOeRWCL2f2dFKlYCv
uRuTQysoIH+qMQpMIOJlFZpmDGZhUpzyjuEfstREbdadnO5KwmF9MXjZsMgW9zaE
UP4GYmYZ+Sr4zXFZTPrn91yFjx+wGIMvZVxP9dkQBpAcVBXCM3IctiYCNFXnQ5qG
Mcx4qMZr5oHrmcSJ5Vrh9jqK0Kw9Ieada5ILoXUB38S/QIed3Y8a/usj5Ub0P2mn
p1n5acUXVenMB/riqzv+BzAwo2NcfGIxphr4C5ODOrzsMmW0557MkBF8yM4+eTQk
tGVTJRnLG5FHfTcuC9PBt+XJm9JscVUO4CRcoy1WIE10i+YkcWT1rXnM4vdoNdSi
O0yV6iL4DdK8au/476pcdJkLX9n5tBbn1+7BBRwmAbYNj0H1VoRqjfB7DU9jqPSm
x2EIrsTi7wcSS3VUIr1aIHjSM03nKL1koEJKrvDjMQhrh/8feIfBMhpHDa8VOBHy
LCZ0Cg8IXS+/XreSfJJwLWMRPtS1gIzHlxTUU4B4OhedBsfjjoXPvStgqpwFd5++
y3yeegGOdYCTeQJblptGozvu3TAcv5jBkJeWL/38FGC3yPttI8d0wMR9MNTxQ6rX
KxITzZGFmY8rWtRtGpwMKU7zqg7Ps4wVRhbfq5m5/kKt3jByx41tLcgNqhRFIaOD
SKHcFii9QTQP3mTS87GrFzbXvm9ERmot44jgzoSWSzr2IAO/onCn53hOEHykARTa
bghe78EFRR7GkUclv4QWyi3Q6DxDkbxH3F1NhonBHZ7Wy58EkrTuD597Z2qcYhVh
Jlt4daKBsdxNtD0aY4XJ3BrrG99g3FBdwUoF1vDbicxScednDdP6/R85KqS6+Z5B
UmlQBIr9zDJsJVUTuQM5pAS+jdaIkAuItInWacbEtrulJ8UW33xmhPepqB/Wlidz
r2JfZ7mGwASN27uu37+OTaDi9jpTfAKTmtAANG7UN6VGpSOw1m2R1PAlVsalEE/U
4mqJkW+s6O2Rnl2BOt565wWmkmVi/VQTD3DKPgstxNQNd+SfKR3qM77qiqez9Imi
zSFKN+hIGm7IwIQytFc1hQHTQt/MZGHdjwW/fxwMkVVFyC4hMgjw5TPNaXpBY3NN
BcnI9HzIyPoZ4XrHTXXGpTvbhwLYwUWch4uw+Qz/sI4PvrqYjJKaBjPMfNDIc/6U
WOXvH1jPoBLmJ9i3VuE0eSR/21hFWMbmgg44XP7Bn6P438C1NGi6f9rUaLspv2CY
vsDoBhZDKEEDzy58eXC9cGaLyHS7s73qks109lICMlJ9WzXyXs40hjS61q2kPW/t
czNcpLcowcMeY1TPZDfxcrMB8CVwgPCmOM8/gorcaw2OzUnsLaJPdJ1A6JProY7d
Gi8NOVtJcIcTtUfJdQYj5c790sHoCwYXxMtge37Hwv75zgUgXi3go5SmbOzU64Zs
Zu678S5KeWSKK/WF7NccNIW29F6xTREK5YfHKuCq0PqjhRoPeMdRP3xtGhg0brvx
0tndpKJZFp7+ORi+V8pI48sGlXa5wF2rPDPWWN17hvspIDqiCwhpqgKM6gaizAnM
suneTwpHKB61QCH8JGbi0GF+APNm0nJ3+71MvfDPa+6WBL7rG0LUjEXWHNhx6Q3m
NjYTwst8zpzbN8YMARRUWmLJWiXOcCo+16Lk3GqP8Psl/2DmTw30YwMGzoGcyl3K
Do5Vxz8fLa+ndbacG3zFWBppWIKcuHQGfaYB4zHPn9ovZ4KN2r7NupXZk7GFYg5Q
a1xHGNglhCZ7yEq5CnSv02/CQo+y3yNNuwnQe0SeNf4HQ7/azzmUrewyQASN8xtZ
lk4najXL5wUTjKBq/TKs0XRJpIySM+8H3Q9yum+gXDR2WlWEuM9rQgOjWdYMjHf5
iimggN6CO6mdjd2oQwdjsJYxwgXk9jUxzqFZHXMgncGNJm8lH7TCT3DCwOCSGSio
XrnOS92RDXKxbYg4fsuGyP5IzX7UN0qXn24RwoSoYbKKsz4lh3hE14l4V+KS8Cip
4bp4+Cox4TQZSsSuQ0PMfxIOhdPS3ye2Zt3l2bZ4kfssS6pqgtSpXNadaQfRpWmx
Xwf4v6+w9iHTYYrV7r4hLBkvcYCHHPKQq4fc67Tz/WFxy2NDqsNX26ZucKbAz1Qg
qiKnVrBelSCQt3iaBadG/NgpIHssgQPXUCOYOBT23f1//sYOqAOOIv5K6siRyykV
ZmM0CRWg0Gr9fBqsDRmaGDvTFMpkJ52sQ/oHw37OGcHr08tZi1c7bM1IEoZoPwRf
l00VHfXPjCgl4kD3k1qyookLJ/wVry1hQCIAGsnNSRFfU5Oqyx5Sacc+JU7fY9TK
Q0I00171Mcf0Oiv8OdIkUIk8gxYmmfWUfjyRH2bSRdUITXfvnfWMnCT3hTBwTJFg
QhYd6u5fAnYAhlvFE2GqngwJhUEYnqpZn2WRW8VLy/NrkJg1FByeHXAfgUuHzPKG
4PNc+BmxT2iyw58kYq/NOAvuFM4tVe25kebS4wNDGmnB8eY2cnAfBoQTRMQG+ezy
SkOUjc2n9TYaxtIMoQU1TsXC3ZJpIZO5a96LozOcUodVZmwKwsvCZzIcgIofGZKu
VWPq3Q3CoMS0mqEoRqDLesKgsUk2Z0l8CAlTbFTM6ZAKBFpeYnwtpYne/f9D65uy
BJ10z9iVllUiSXjpWK9kpoABkfmT3GMCNVSw8wlKg8OaoMxEUxHyDXGL/fM5wjMO
g2+90q1pQkE9nima3m8H2rpuhFbVZHI55TNrpwFKAYqrKW1GMXD/+aG8lVCGWvWP
lsbAE/sKLSqGlif70TOyGhIrvO2cUZUTjPDn8j/TjNLl0VHbjrN1osDnlcTpmQJ4
BaSAnT9nl2WKjxwZzGGTVBaLR4kz/VJUda/3i+c9qCLHp3S4O/Swk/Ye3YAX/r37
D6DM1c6bUd/nIAjEu6FaS3llSo85PPXOQHQDeaoQpBMARUKg5VsLCsz4Q2sPjAwB
hnZ1Ze7UvMQouDSbDGqRJ8VD9aVVgDJgxhlTlXVpcGOr5UKLrWa0v/Vn/BNA0tQO
0M+UjbjX33St2sFUc0FbeRvg7plFobNVk7yiAchUhLreL9za0/UBMjBE1rMDxsNS
vH/UYlVziLiIQDMtouChL8JXLBN7OxSOPkr0cqHCLZG0n2iYsW/SLqOZiCgND6fc
0ooKmc8LmK5j+S1FTJFUFBlFM6evH8OrDJEAsB2srKzYYnBOTVbAnUSUCg4+Fgpn
nZOg/tFjl44n11T8HYdy/1WpuejMWjupnqxhrbCaYdJlYBQPvbQruS8Z1tDkClwW
ls4hCl1G2On7Dj5KS9M7DebNLyn7n6LU/sPca3atd1abxT7hJuhBTD+vfuQN+UKJ
EMrXG9NXZP3TSbrM1dZB4xtOVttk9K85/EKN4GwCcX02vddOFIEbmJGj51YM51r5
HA2Xp3pSn/0SBkPe+izMdzvKEgD+vS4RU9nW5u6WLNa1ySj6gd7AnPWy6yt3HFGF
FxyP3y7CVAm9eCWgC5Q8/gGqpaUU4F0IOB7yJl8oLgjIj/z0kgpE/CMx0cwQNoDJ
1pxmJwHPrcTitV4sjQrB3xlxP0FPjZD48lC9hE149bnqT2ibZv1py4rr92rWdOBZ
q07SyFIs1fYNLywXPLFMuD62HRYyj8gP3fF1PFaacUjuMDodPxuasSTeqA4z9RsY
Cg5coZewzBq64Mwk8kMbVC+yd7CrpPS2PHiuB2WPE5W1OGpS9HPPL6kXdBy5kFCy
2vOk3rpEqiW5KijckvXDhnK2VekSAQelVBrMRCxUec5YvyAQ/kGv7Fu/XcWUojT0
yIoRbyRtr58cQs36bxY7AJFUrRpxztUfW/U6fzrHaEJArTndCabOrrEfIo4BAOKj
9zBfqj81ZRy9chS7L73wcSs3jroPo3nQwRPOj0zMqiQzcW5WRkTnRzMQZquKVQNM
8AaanvPOZ3Moo8IXkru0JIN1KIXvBkxP/VjYArZJ0F2O/Iiv/RQUWlA4wsA3rJBJ
lj4tpokEkyXpWWOfAHtDq+P2SDYxsnKfVeUR6uPknVduXek+naeYiZEvavpY9He5
N7P6kJwblfr3nSGdMyt8PEKVOWd8RD+7nbjeN6KFeqWdO9ETZ+6eYJvA8yActo9C
YSNZNyKUIF6GexDJ+2rkwJYfZo3PkdZkmW9O0ouw7FxDyDHRlB5E0sFo9Um5rCSP
5q7xzyu4m4HGXNgl9rRXk0gqpRAHWW+9lrtlGScDR4rMsFcjiSlL4v6+LaMDCV/x
YIqHTx7KVgQNml23aUGoUZUbfd1UGAjvWXEkKuZGBcol5FaciMwq/GwpqSP7iywl
wWWS8CBVWRXzNPqo722/MIES0ZZQ2UZjfzoUH1tBXOvBU2NvvEHx8PPOHNu/9QL6
kgf8QXI4e/WIXxLBE78N4vrw+Y1aoHx0O+GHLsgEyu2KHxojLXgzov6Fwilg5MbG
We1gC/RTZ6SBxOSBndHK5LfaUMwbQebNT+TfyXisJRGrovNDWyp2Uv/TCkfnDfA5
p+T+Z9IWO3GfpiM2d/UlC7d35UWIpKYPVCgWcwA2qa662G9UXOo+KyCd1FU8Yq6l
+2oxWdrzyjwdbWLFid3Jh96FqkSDw7GyofoehgL9vAtI6Md90Qkpgt8VtLObbN5H
NKqrnVgxIMLzoG8UzyWA3aqQDqPZZJRe+KV4Ibq2+LCNN0Qlo+T+LgA3XzFb5nSw
9GGzjraRUycPgeEWaxdHDyWjtFGFwQ5a9c/ZwkqEdQuHW/+W2UvlTeD4fWnS3z4U
nBdyU9G313oMqaSpIvBNCStiI5R48DhKL3rA7jtB5ls44OifwadaSXOhr26gHQlz
mQeXQ829wa8UjpMhPt6nBSwxCqRFQuUBcfa3iDPh+gStAHryemigc581B+mdDBmc
8MQnaUOMUY5HO0qtxaezPZ7z014ZTt7NwdWVV8uMtc8gHsfWyiT2Zo2Byzbhc++R
0IxQDQ6ab87FG384AyZ2vAeq1hLTxHN/r+kQjahUK+hgwg4+GSlSs0eai+joovUV
TZloEaB6MlOoXiuXW4pm5RGGb1r0GEN8DgDDERBIY/E2P7/nwqW37vHbAG/GJi/C
OO6dXFwfVNpgMordWKHccUkFVk6QoFQjaKkmgX9PLmOEHoFUzf6/yjrBnzHy8vnd
wXUvLLJCA23YnelMHBLV/J4VsIU+1O3LDVMfeGh5uhM/qqIWBjEkZ+S0azMwuzHt
TbrxULRFdXFNEZnWoKCO++M7TSIznf2MZ7F2UQagfM3RXk6FKmD7n78UZwlEF1VN
HkRA52RwZgYehrejLx+nya0rkKJS3GmNucRN8siKOjPMGjbzsi2AvLHfU8K7SieL
u4hNS55PB5WEMpHJH824w5Ev7r3zOrgrddi5hIE6r09yHHgOumrnEVPO31/XV49r
XPX6Jj0m5uKyZSiGYRku2qijvLkCs7RDo6ykgjnrr/xLmol6WH1rtv6o67svYAyw
CaWq5TyvGqwyuUfQEE6+gYs3k9iC4Gkup1FKxJWblXuMaaYGfOhw+02T+noTuyUb
sQ9AF4M1I47HKSWD5TEn2YvEMGar3jpi4rCkP6qdfdMi6/nHDPj8uePVTpkL8xvk
YzmJkgTwsmkNuX6AUo87X8fYN5/emd5cohLkwXI3Ep/gfHcfvJnJ2kWR8G3F3fs+
rDfGoC7Fo57IoOgDmC4DOc2FxjWuqCDb2CEbQt6hgWLAWYrftRuFPyImDhagInWQ
iMy8rMER5xl0ueq8s0UsE1Pi/LS0BFQdD3mEBiY8XmLA3WTtdFXZWudmMfvZ/kw7
oitpc7j9ql3c8+Ue+Bd5M+mHL6rD0Jut9RMsf5Lj0/kjRJVJ7nfRPxom/0h++xlu
D7k05DCo//ftDCs2l7JOgvFXpUF+b6ypaIusofGnNVrkRv1t7OBT4/erQO3rqudN
u/OaaRQ4+jnIKr5BLCVmTEGXu/NmgWHKi5+pd/Z5RE61h0q3fI/9gmCgrOc2Cmaq
pGCARZygsn6nih/Q0ULWHuqgcvQ70oy7D2ePHSjIbLyrwRmaqc1452W4M+t7gkKH
kS9p6efzt9Zztqyngb/th0XfHWXP9SjfNoLp6x2PWbHUuDfuOIPOYzL3RIBhj+kb
/lnyp7sYapwOk7przFmQhmGgZ8AMLZfaHiIEJw6HNFVykXNtiNiggb9n4YZrMJ8T
F7pdbnxYq0tN09QsWOZSKgeyOFk67enjr+fc2pyhfwuHD9Hk6xGGMlychUg0iiEv
l3SP7HVjH7xMHBteGjABIY5cEF+vUa6+eORKpyoVXLbFmaxts0x46swjgHUiV/zb
XX4PiQ/mFp2RYqNOz68oQZthUhJbg/q74gOLsuhSIN+HuJkF5Wj5IOxn6zjnTeR2
aw27pgT3lhiwgwPnIat/tQneWRthN9fRSzq8G/aMwx05Dv/v7cgKc2Rh3k6lPO/+
klE2hk10ARCmhISKcQ0f/6NECL2OOedyk1sXYd+nGDUMpT6pN8ZL7LfQiaZI5Y3D
6c+sFnlaSuyj2Vkspm0u7mNtRuZhzAFhxRb2tomZLwbf4kYSqg09V0viT22og0gV
SAR/qvrwZrqRY3MI0+SMl4NesjZEfuAF5G+isV47yDvKSfFsKyvoWHwHhh3SN5fN
l7AuYFFtDDPHfUJpo5Kk6O7cQYHC1bVLzUb1ZpI74bad4Gykz5hD39ZuEeWzczt5
NP2TytXErl5RQZ/0/t98BaN+lK9G+ybjbOBH1njekXMZHLSngsiIaqwC7SmOmons
0i8q5EfLXI2z3e70s7HdSkyqVu4KiN5orPhOOm7I+jQYx4ENHejeF1O/jNHD1+C2
aGF2oLwsV1vJzauI5CL8DYo74+E3vNb47L+EJFZEDR6ubE2tXTWtrmHDLWbpe4DX
H5geU3jcmj6tybTqIkMAKXM/SiiEKN9fL1l4jS3wTFo0K0vP67urTcg87FYY+rK+
fXMjJKcf/B7EooPyRLG6sKpLkwKNrrgwAhbmDZIeNB7vdkfdQtjGEpgWDXEjl6jR
QplFXRVOGUWz/SN16ihayDk2W10zP2vRD4QJuJDIsyg/3rSysAqoNiMREarYy2Vx
Js3Jwu/YyB+2K4l6KDeGD3qn/sGqGiMjr5OaH4ujAJyQOXARfn1lnWaIszmEvatR
x1A457AbXR7xpIiD71NwGmg/OXa1SQp3Eecr+HB78URgZrsEQ42nDSbKle/I1b06
c5KxFmcGqcdbusMokGpj4XWTyX5uo5DilTt6FmHKe9XwriWpNYSW3ikUxqI+waDk
EN1d21vy27QKTCJcWLvvLTnHJWNrLtduwClqtQaogza6VeB9pPeecUcZs+32STvy
dR/v6mhqjUDhvZJlk970+7IoK8Wa1ZM9Kuu07BSLyk/6ZXtUuZs2FtCeKMSMz6Wk
BhoUSHSUycj7nn6/xy/9zr+M1OFaHS5Sm0F7IKFDvoMPky961QydVdON+gPkx7Wo
Intg3jCkw55+dSHm3tVS8SYnUqC2aUM2unD9J+YUzKv5z1W08wLMm3GqxJUjNvq/
Rvg2E4GXroM74hXaNnEQT5DS8YAUbLXytGkAu26nsk+k5xGnw3bHTgAMTahGt5RU
rWBFLp+SPnrO1y2bXvcjvutJQ6rM6FPcZC8BP7SeHcxyaZ68sdPZaXK/xgdOp0nG
O32dBqtURVW5ZzMDA7GEx4CDbsbgeFx3NgwNd3QPoeX4BracI3bGAUtCcRPSvCD7
z1cWR3Nk/rL2BcN26dG9JrtDJWIrcjOobG3kafFV9mVYS/kPpv5MJxoY2mLhw+eQ
tNYQti5fF1FKEecsvPyj3lXLLejXMht/7sFEfGOjnrdvOI6rUjQm++0YAyEQYoh/
gPjDoQOtmFCHNnkcP4vuCoJM63F+kc3z9eUN5z6PQnHrkzR2hLPpUK+/hTnwAdJV
YxEhIfC9K88CTeg0cX3hIKBfNp3PJ6Pj2WqN+P+pDAF/neWQuJZCex3KSwlmweKL
vplAInjSVwyaWWrmXTodYgZKjIDMH+FkOurTf1U91gKx3o7yWvzGdlANPGclQLsg
ppDScAwLPDS/cwJnFsRcA5ELGVEyRyq1sZIP7UOm6cf9ozcgM/lJHx29slxbphat
JSB9TviJk/UBu7JoTFEupvdTR/tmFZPrp4FMlsP9xRMV1cFUU4NLE7s6WyTgPH1U
6xyK2fRuMycf6laYK5Ena2JNZjAmHwT/+hG7M7UO4ci7LIlqNx4zF8zeu0pjJkb8
hVJZnTUfuSLKRkAL0lFiDLt0EsMExSYhUHa1m5bxuxCw0MrmqxYG4vgqS97Z2Ngj
ozcgfg2It7pcDxgDRSSa2k3YN1Z7BFOL4gmxflHsAc8qYxlu2I3GT6jrj6xdWv9F
50YUVXqS+cj55JLN8wbfdujdeOGwYgUO7VI8gU/cXUdM9pibkNvr99I6+Mm8JlCY
UcajvdHaTjTsXIMTIBKyfr+3X13kHEzLPBlWl8AZ2DB+7i/1wRYmgKicIUjWklMh
rrNGuSbJ5G8u9OGAdBItj34v7YIy+vHbImSfOCoxXudiAoko8YnF78QLaRWR4y+j
kivrXP8SL9Fw/mrvuIPcfekCYT6ZoX937o8mqd0EUAMzUbD1CRZCk2FbnUfHZAP8
OSWt89Lw9HHv8pBH/iDY6AQPz1ZAbG9X5Omgl0/U1cfdXMmMdMzNDzB64Ho2zmER
eDwkjOGwf4xm2h0v3gGycq3YNrbrb/fg/iRZTy3hOYF5zzk7jcN0chtnsM6W8WMJ
dDDVcQTTRk07ANgeF7zHlgbz1dPpRXmKJA9oHOgZzbT2ITjS31fQMcXEEgspoKmQ
I96wrEBvSQLRpWeaZKbL/GEmxu4NlB1i446tdc8fNbMzRxw9mx6wWUx7VTcHOtoB
CkymG1ZqXzxYRU6iln0FxwRZ+eGKjOYbfiXNYzuBEdywpip6tNlakjHPvexXxnnw
+CTWHi4SB/RF5Kiqym/WjvdJFcDvpngeEMWL9ucXX408XPug6mbaGLc2x0M26bwT
JOMx7iim6veDD5cz/kPRzIleNUFyplMAitY9XWEFC2d7Yb0SBQUH43M7axgnoptd
DITQQCCOYg4GtH6RUmohFQwSBvWu5CtH93gNdL1MDbfDdZ9+Uwju2CiD9oliR6iB
4QdkvIOQtlJM+Tn7Ov6ytKRHm/YhmQe9ndVE9paJF18tUtqpQtbSrY9YxVuN8HfT
bBnskesgO04z6P7k047bAGnGfv+6mNtINDmaKON/d9VQC/Kcn9E1MOtUy5VBy054
VDwGIKiiaKiWuR3tABJ4H9L97vylrtjBP5NnI/nybl0tT8D8NAecCKWx92aCvzzo
kX+EJb/Y3bAH22qFSFNLUOu2JNDJIm+kf/X+qIp65OkwsUiihoeP669d7zL6Gf8p
M8+I64ew2bKLOqkcgdoJlZejI7prRZVhu7/Xe8+zy7IRp4MHhq4EjpewuAnn3a30
VcYOxHse+PrhviJTVwOTByYJyfJXlwEjgpwXWIjr//JqjmQkDPOmtGZsGasxGHl5
MjB+PrgzT/huxfFVGa95VbWa8spTWQVcxf9CR2gwQUZalXuiPEO8AuBpINT0lIZD
zp11nAPRChP1goXbAis4vHcaETn9DWs14CL+zb3/Wrw1TrLqABfTFPuZdplpGdkf
g23fUl4rHOFCTY51GISnVQEubIEJ4SCR8aR5StR1OlPmrh281bmtZwW81WkUg9uL
ONXkfsnqEpBMYiqxzqLFhXFMKnXwmLB10CvPTULYt0gVosvGOzW46uFAwSrSM/Hh
Yo6B3qs/Q0LAbCyh3XFpE7xaKA9JbYZ8EYBkwiuKzLA/aCxSB37MvBLvUub6UK8Z
m1hoZjpWZYYxJGzBi8s2iAiiFBUpkZdYWJ5cFqi8gbaYuyvAoQFJBJp6ztYm24zW
K3L9lbC5mStT2mzqQf7lheFvUaPeYTR+Q3mrBjB7dhRpoohE7nOj9+4yP7dgqHt2
UT2TSGe2WX/NVUNB6y3pWDrf5z8CfSY7Cy55EJENTcY2xNw75TXm62oorATgmsuG
V835eo6NRWbR6QNV3TK+0472bAkAOtMQUWMACKU0rPh9c4YCGqkyZhwbvange4lj
68kYEOrn9e5aWo4uNB32BoNBmzfZQmakZd9jD46vO0n49dy+mnIv5oeamQ8CyO4G
ZXumcVIse6bWgY0dQ2Va5qdhA2MxX7cdCsyGax7YJQUfXS8goHT4gB7qPLwM37Kb
QS9pTM5VC/JpY9ulwFHQMbidjtl0em0mBVIvs5cmU5q7RHsw2SFuxAIRc/55Xy1N
8k++kSISVsF/ZbNQJ0ociiQuRRB8HFbTiELuWI/F/gfeagp1aiL20kOaP4/HTxCQ
qar0LuSLtyXXgCBBN8lgCS5FjwNFokgAIBvRa7xxGww3BlmUGfg8uCFXc/Gdra2o
ZWmzgiBMF+hT5E6ijzodziYl1IBHaWMclTemnsH7T/JkcOvjtwIPHr7ObG+WleMc
qZYZoL1kFFpq3nXHioQEdm6yWSEXdZqZjlUUIGBAq5Gl2vawPSwaZNIuxbph23tF
R6gT+qPEB2qYaADR44awuJA1vdKagJYOl4lASBM0EcLm1e608xyFwAXaxFiplSpA
qA//sVTfQb0KK3izrzC1imZY6Mj+7PufyhTdYe2LseCJ5nm1AgxUYStkoX13PXbU
YqqMjueEz53vM8wLK/+bk3ZgMEZVr7gdcojfPYDZUIvd7SdJIj/6ZCbxmBxyearV
/+vidl2Ex7WoQdHlzZxzHyNJ8GHez3aYRSitbJBEsNrk0we77ghO7/gguL7otKTn
kj24aM1xpG444XfjsEoiFa490p87yyKHoU7yrlPxNqxWbs6SQbILQ/D0DvM3UEww
onsnNmlGeQjLeJrZwXL8wy6/o1BJAx+5DcKPYSheGmh0gxfSz0Noj3KuTkUDqkyK
/7JDfnOctaPFc1hYnRgdmea58tWjISaPDQvTApLlT4wRaBS/DZn3SLMpNSbxFMdy
5dYmvVedFyi3ZxXyxe+3k0GfRl23PGDJJdha+Uqqj3jtFxmSP51awPNumyo5iBei
+R+0XuyyDqzeATx/pR3AgEwX1bJn6TbcPi1N/DXPA1AJV6Ow0oe4NdOPS6NxpFm6
A9Fd31t27qgJ+HMuYF43Gdoh4MRWLsNJS1L6t7MdrOd3ISSZ+qp+4xr1h4Nk03Ht
9MAltI0xQdiHygRQOFxwb6csK7e6FZ2ZHkaplF/tWACgq+60hbzKfaM8/6LqYzoa
x5vubKRCNhduhnV6QDtmCbKdGzJGXzYSBv4FQCILf1/qBDNrMv/QMqhE+YO5f/Hv
c58qnWgbrJyTC26v1p5LWNjxepYXexRA1IICbQceEjqjh1sJTxqTDX1XenbRb+r8
wK7AW19olSbkNNDJJIANLVdMHWlKpxpuITMLoa8LJX7XtnZ3bLJb5qbPwgujwkLk
tmzMaM8H+rnmRfZMAobp+iBhui1YtJhQvLuPCsawphFCsxQXPgJhyF/q7R6mBmWd
h1oJiVeCNW0yX2vhnQ5YKiXe+ALHjWaLxhwA2RGFhRAHkk2I+g/ixENNj3fTrEMh
Jp48eWxo6E6utqZKVuConrkJCYQNromG/jsUww4ew6vrBbe4C6/vgVmTtXFeyUxS
y6Ii8W0lHrZWjEYGU1GIGXqoZqBZ4/WKMQLRRBuJznSOEUra/3QkzYlOL/GUeZme
/dfDEpVcs1HGsrvJgekRIhQDPX638xwVSLtrmh63UR10sbkhyqy+FOIVfh3lm9D4
jB2hLyGwV1mbpmAzeKw8sLhJSunnGbWUTSlQjV02fg3AhQ7yTFFijEJ6BukxzVqa
AzKCHzrpzV4bi/VRJB2JdKTus1z0nSg08w66Dd4Y88Cg6/m3RyTo3zJ+7qOddsnJ
uOqIry5JLzMJxeHH5Tmuvuu8QfmObcfIG3l40YQWlMcmlV96Ptf9odf/Kg49RRfg
7kreNZ7JEy9lH98KA1OTT7SVfiDN58TClc+ebG2eVAN1GrdhEhk40TAauYMx4Rp5
g7qonJekIJeivI5i4TGK/A0/jA6s0d6FAfsOByhzn+QV/XQPePIP2mts+JHLz89Q
2Oj9YZsR0QLCVRyvw9yvXWf0PaWQ+pC9uTko8inFzRwqoROw5zgsXfqKdp7OQ6rQ
Chb76h656gYOZZgxK56eXtQtsTkLhVuW3W+6ULAzcDqfHIi37avEN/VDPmPbIS4k
/benmi2F6ajBogc7D1cyo27JV38NEtyjdEpGTCL3R+QdLmHC/AApvfVmGUyO3s0T
8cAVukkvIIoHv+Nqboo/thLw/YftpLh+8qB5psHcxZWdvMt03apCtz47n7Z6dalE
AEvgWZmsQ5SJaVa7K3y2DZfwn+7Iuxf42fJOYPYpb3S1je4PRryq/cJuO4Zkhlf6
Cd5Viobxg00VuA3LoWrnzoWc2wHoqc2+Ir0d1HViGw/2rr4K2AfMMpx7KjozKkV8
Qk/T6vw2405w/PvZi2Kv3ae6iJ2BJMGb6orLXx6z3Sel63BGsfhEwPl7l5/DOUvq
ko/78UJzgg3fm5lYga/0imoTxXFoZqxXxd9lowTU1UalaXZhUoJtx0rh1IPfCekV
98hTCTLTMA/495bINbHtE/OP8KSMqfft2hs9FD5TgZVKpAxtQoDFptntEglfp6ke
NVPNBuuYmEHeRL9Vmn4AlId4mwbjcISLz0DBK0rVFyaKU1PP0V6yD2zMzfnynszx
587Pte3yS0sdhUtnnzaAmRvTmxJTP4Dj7Fgwbf1AbisnHR9EcDu44COVaLHNrKko
88NvX3v7OqhYO+rcIc61mKc3tvAQ8rzRIb7OPrXNhyehRD5tWZr/Tus3NF4vj5Aw
48UJuiczD3SM7ZptMSGayKzbMascAmlFvTioSUs2i6gVYM/PyfIhgqo86OET63KS
XPAzLT0KXadGatunPb03uan8dXDRrPfKZdHuJPrs+/7laXQkTwBJTwzhMWuwuh+j
bEnvPwLoxMgemPOI5MUuw2GX0BMdZZggh9k3SaLofIDsyOeWbk7+ZF9vHkXA1mQK
PkH5U1wcTJcvWw2JZ8by9HdPklYIu+jEV4l74zNnKuNzdY+Yj3TjkY9iT1ON6N1q
/E94nwLc3MiO5GUPoWkcuGkmOn1e5HV2tTwedsT3ezlYVW37FzRlrxql1+aoUxqS
g93OtLUvoZt0DCEapFalXM6st7ACeJ0/VSkCDpM3m/GvGBjcIMP+UbVE2sSzmzqU
txtKfA9Fuz7o9rTv1/NAMBVmrQFL2Q1Bf49Fzg8vN5hXvtaJa6n+4U75G+63mmTx
eTFKY+GbiIoL3iO4N1O3h9PQC8hnHs2dmH4+gB0Z9qiVI2CZeHAl+/2cC36sAX5u
ma1uDUQYQ5mZ7mEnOQHsRa91WLHfFzVP9O8LGOuVeay3Doa/YbgrqtehN+WUMAs+
ouVe27h1PjLq5WZkhw9THQje66L3SZOL81CaB9ukp33bx8OoCpfTEjBrhpSrOPcB
AbAikjzXuZnVDVRMRahS0iWBRmis/MvVikrELi/PI7bx7/GA/4hQjIaqZ2HEij4c
FMUgRPpzAImbkVVf+8sOdmFbt/KuW9n+M3Z0Rv/FRK1yLo3/ulmv69owzIVgx7+2
lrS0ILxnETm6tt1s0ikm7wq4TsxyBI59ztn8JP2bcr+IPu+4blPgAD9FqZDhYx1a
KkEsZNAoeAQ5vxyV9gw7bNbqIzVkDF0ENudx2jaxKro9TTseNuVs86lKGCd3JpXC
gm2fGrxn3thlrcouWh1jJB0yqU+2zDFfZbbnMKuQF/cbK7Z0MbupBfsth+uPhUHF
EZ+DCHIkD2zd/KkY6fwiLiI3gH7zn9OiiL1MJza5+QK3BVSzhIKoS5jIFKwgyeCR
X5qgUF+o7OhnKpXQHK6HStB9WB3Hkn22odjStFdaf5qnbsz33eJ/mdN4lVicdwwE
sqLBErGbcVWEAR6ufCfFJV+JWJlaaS6uUf6m/04dBzt8BZrNy4H7tXJNAhZVdroR
d5MWO7+e7rFo5Go6+YpCbqFOXDUyYlP8HyjgJIuI1IABMkgOfDSBg9gaw7hI6dpT
per9ry3fbnNt6xtbGNBefFlhdSzziReGNBy5JcH4OuWbHY9jWE52rckl7kg39QGh
9DBDy1UGkFYOsFHTDC3Cchh4TjzLI03ynnhaDuA8Mrt2Awq+xtNq/DR7NLUuQhfD
7OwGkYZ2bx21YFGRJeFJ6Mt5A8BkKJXTQQ1h5JgAqewq4/rf/VMDaSR7zkg9N3UH
XdKcqnqUQhy8W5S3+biH0gm0t33ipn2y/hY3Oi7xOHtR8GUKUNA0oghUkR1Gw78v
O65vkIzuKPEuCO3wgDzlS7ynEk1dArTA8PgnbninRrSLrzPVNHOfLfOVqV8NiTuL
LV5sknoz2MSiJ/Jxm+mAczMU/n42+RdX9lVn45i5VkgHvMpc/FX4UhkrMr3rEMEW
Fe4bwfcjsDfrcs6y45YFpi3YC1mWuu9Uo6A51AH4sIl3wBkAsGyr4bO9WjMWLBuq
DULIbaKmTnNAJX/OBPx/7OEKHAvT4FuZrq9xofLELd6IUKVaTXfwwUHZ5Hd62JYp
kDxJJ4PwLZLkDWTDTdrHWrzdMG5nBA4AO8OMFynpLqaf5bx3gVYba1AHnss/WdOu
QCNXyuVsL2tANCALsnov8NHieAuJ0CyvC2gtcHLJ2cEKwN151WeVjhvuUNJEiu1d
GXaCz2U/FKo+Oqe7EealdgyBXuwBjlYd5SB87//jy1xXjqhL8B+Bpx97c4qnHHC2
80Pj3XnLZjdwFZT9UQNhedmHHLNii2IHarkf/RnkwFgrxAhOJ5fNLAb9+cESBoCa
4W5GJ9ZYw9YOhbyegIWjxpsBNM3FsxnOK6qCxllj0wQA9/AA1pBNu7b6g6OOwdql
Mdy1Byqf0erYw9czfQu/jPwAoOmhCbUV+nk3sdE0LRg+eFbLp/JwTQIAmSbRhsg1
VwCoV1vfabBFMHpbcGRXFdLsLoj3nM+Dn0TOhqMCQ7A0P+hhKwtmXWzA01+0+acI
XWiKq0b4hStub/2aujdOs72+8KBpLCMC/VeZzu1k2nL6+6hvn1QOO1KnaFf/CvzG
oYrimX1NgiOijnsng73RYzED6N3kvEMCiHXS40ugYMPGaXF2OWIO0TdVjpceNxcz
GJJXSjEAvHMPDzO8TeC4lAE47mRAT3tmdydkZP5YpVELpX5SWI2CFvSgMOnhBwKJ
Hhynk/hHdt7yq77eEbcxwlSudKqfZZ1S7ddBLvTl7LT/wODqjwqTbSKwPX0NyWCs
XgiGl2RNkMtnw96eg2HkZXG7jj2XUYMvSW4K3wJbF23fFH7QBKWdmy1HCdM4MZRm
BJqdynHgrx9AlsdVecVUeDrLwZvFMxCuJq23lo0WJftQzUumYnpGr46j0ntyZH5H
sNWWyh3s9SDHfx7Ng1LoaQQ8Xv55/w2sdVYZ7Hko7jEdYHuiHOmrIIKhhCOYqFqU
EwqV+uxBTizqCfO5QQbd1REdhUqLFx8ahWytsbEs7Aa5ugDLJC+Ba4dmnlJfjlIb
yE6b6j2nYrZS75hz+sLCrN0eBniOX2ot+YMbeQC9Uhlo6nTERx+s43I54/pZXF2h
MNRtvEbIHP+/iWWWPvXqy1+SiUmt0gxEgGtoeGUSSmNgdl26gk0c7BkBrEJK36kt
2rXghmM/iqV5i7UGt1vrQkJAu587b1Chia+MWasP79ktu1+VIPGItXlwOSah1N+4
j1v6THyj+IqlPi4g76GnADQnKu+lSN48zqDqgXVJI7mPtVY+Xx2uvufVOh+aUPoi
btddYvDrSOsbud7B881yCLmhNyLtk9PHnJiOi+nvA5L4oSerK4kFzvJ+C1Q1RPuh
C1qNZt9t2aErdDz6xl5SJM70KC/a/KhsNJN+y/Nwi0egjrBlHe2Z77wi2AzkSIjb
rwEbvOcComUonXQq9i/kdncDTcVXK3eVqeP2lpi+ECbYs8ObLZRMlxlSZW+YKhpq
erVOdjTAwrg0eFvItYIXME+G04/3Uae3EaTZhS+fnNtO2FRlHY+97bXJq5F2WQyl
NWai6OwNmVc2n5at0+gsnnmmecP4DENcMvelouhxa05WvkaS6T4xKQrnD9ztiq5b
jZtzLkU51RpRYFQiKq5+Fgt4+Tw/WUnenv/aQ3PXIiDC3uL49Nor7OOquElW4nO1
rcOtX+wtPUrgPGa+l24890+LTo2cGicYOa6GkyGIO6Xr53DeW2OoGRkASqn+UO+o
7GLlOztBp4DezPpG5rg4DiqMnKvknlhoIuN5B1AmGJBP+QY6soJ5HYig+Ccpx4qu
KOnjS7o4bRxWb7CdPGtAtvJnobAizIjSUQdXMFyCx0VWqnsJF4WBzK+AXdY3OBcw
jGUenQpb2LpJDDOGwDOju1D3/ugMo/5l7HwO2BqgskGGzPPiQ2Z2PmrCbYvGSW+Y
66BuQc+vJc0j4P7f++gaGwGxzwD4ZXRwTcwY3H+068/C4cg44w47EVO5p7rgK062
JYd6mCSVt9/QV4M7dBu6t3sxSFMe6vC+WwDNfddqCCMJ+nvyDCae2UYKiqrV/Gol
SkNckSbFuO0p9i7MtfqH7vTYebrCiJJc10ydVI1/LFUrmXAyNF8t2JRfD9JpF8GW
HhQvhy0PMD41FIBb1oE6NIIdYmNFt4/kGOSMfCAcWvHBZrYJRN16tTdCT/XnBf9G
Tir47mCFHr7LihYhtmI5c9DEikAHiUZVcPwDoNt/sfR9inRam/GRDlIUqKwqMuIr
YeVmKuF1yHf2VZTvYfNzETNdXho0DGzckNb8xPBx28uSc1At1unud6BsOBPPEl9j
69yHHH3uqmfHwPLYFqkMZHzmV/V7XT6l3Jn9pvJp1RNuh/UCPL+hmzLt2WJRosag
jZGZKvLPr8jMFUe8hGVHzTui5bX4MlFzZ0Zb+tvJWL+1vgJXNoIYY+dTbnNvynQP
v/ZhK7xcGvUoFrykIHwHUswtw0ZAZV++PoVIFc1jwcBKhnuPhOcR6k2fzi7nZD9e
Ozc1DUOW7I10+zogPmVla95lh20qcc8gEJ3qUs8LKlJNPvMni4OU3TL3wDhg3+Va
v/CTRMV7xKauuVbrVMmzGiuXZ7RE3WWJtoJsYFQY/JVmk3Bjt8keq25gB71NEheH
WU40X4U9BYcXrsZAYf/8414wAyWbauawOBNO2JshD1cGsI2gGROxMXW9d/FDYCiN
c9CfaDeyPYf+jLovYT4tKH1/+rv45LgU2Sb3vKdhFJMwuv0UC+WX81IoNlGIKF8s
Ie/XlyPK3DRce4b8zYACfpGmVrPe09nZNAulti4dny67IMWrMC0AGBaiLlPWI6lY
a/3EhLuIiFlQ61/ukhNye8oDvBPMnauBsmJkX1JtTYRMzkJeS/UsU8M/OezahQkj
/w6MTE/qfbBNnI2ddw5CqWJJZhGHK/PaczfeyrmlK7t5HpCJGXTj1+PjE++h8fLX
l4YQuUCcxilahCN8QSdtIRVd0OV21Em/vzh5Nxb2VRZVu7xukno7WHcU2qTq+GPf
FhOfRBuL4CcQiA2B6T5rD4OzprV4kkMNwT0M1BfETHRXucu5OLK4vhS2WGeemTaS
oRPREu1lQUXtYwp8US2PQu5fhSq1pZFvTtT/z1c3At60oTLa/vE2/ZB9VEbr0RFQ
69wKGChjCO2tiAKDI1HaUSgk8uARwRFA4EnKeNLIQPUmPQMYVjQTP4JWhNRAqYQS
hazY//5Rcmu5+f/VB6xOVxaDwWfBHU9sUtmR4zlOMwvvKaiZYL+jXWmILRzr1O6x
0Ve3uZ6vxL8fMAv4VTiyy+HNfWY1JbX0n07XfAdDzg2j+wx4cbAEaD+2f5LgECA9
PyS5GB0jcgAdMBV8KEW8NbMPJxkg91+j354kQmtfC3h1Db1+9TsukKCtgWL0qJFv
OFe3cWYpwcvVkLLyB6JLDEWZMK0yyK+p/Vujrh6UHXtmDw3beEkaYjGXKcTHioVC
wskwTRCS8mX6+rMT5Y3S70MoWlMQ2WgkRqqex8tTJWz+a+YWANXQ+56c4j2NtpWc
DHKTzkSvEcnMfiMIP6xHpQlBRD98sUaSF7Z8kpc+QEAPmyGseTv1wLl4ENjnzRCU
LuBEItDoh0bjDZKncrBhGEJT0EkzmIhZZ5vL6XsrlFFxXriScxedVfzzRHyhNAX+
55yqX2yDVuKakns7ODtF/Hd48pA8R6YD3yvjBtuHEZNhvvng2O+Zmti8Fy/rwH9K
qRwwvogg6trnTTo75m29sRBdGxL13SpIjvolRy+2CmEOTD54xVTi0InTmY1z6INp
7+LAu+xyBBrKNZkIPcBd+m3FiONwv7Dmhtgqrhojq/Batp3AQTzegYhdx52krDCn
vZ7KrjyWqVZ8U0yvzi7FodKjdC2g9R7f/a0XuB4ejiZuL2F13ogjaLA8guU0KJUt
OwvWyM/4d5vu9nIMa4HImdrYgOfBxHViaV2FuZfzpKLsfsQgVCRbQO4GMKLMCnUA
xIziYm1s76Z7vHE5miRG13oJFwiD7REVBlTDX9/Zy4D41Y4XVRtHIIM5P2jp9DJ5
tUwTCvb7x5hXK8vY62RGIxhoW/X7ELHlH9lGrULWeJxYw6PqLMpzbhs8lowAq/Xj
fHxZRMebb3ckIwtenJQW1Ro3HnBNH9y0hZ93mOb0WApAchJKzNX4WReIQCAHAz5f
1QfSp1+ClNzaS2X86SsGw2VJyzcGQS13P25ku2S2muzfFChtntR2ykHzqKgo25ZY
Ue2PLlpLO2RZyGnEip9uBAiywgv276HOmoRGqIgo6HKIC9qr3+lnUxfctcOrOI5Q
QNxYiezXGRxbc0ZuOD0ZwSBvFkbSsNNWMHbYZzYjRpycbkCmvtiBrCwOmIPjcC8W
Ts4BahSQz+7VKg3qwGAy5x8eGGfd4an87foTu4/jDamDbUmnIJzQXg9D3/xZVOP7
7gYJbUOhCcm21vI5C8tpPq2MgQFtI+eKk54tbfR13D7J30i6/KcwfIFr36shm686
BMEe6KXf9MyEs02vfBHh3AbUQRYyv7fwpA0bIBvxYKN0vMIZmip7H4QsqEWC5EA2
ATYJLOiq+hzcRyncLoVYErrxhI/Sigl3eTRf1xvepTxSdZnVmWglfNzFBl6FXPJd
rX6RvC6VKZlxQN/2le86aT2r4tncIujYi+fwxelbzCf8JwEP/EbOTta5Q4rQhDEh
itedA1EHRJiQTBlE+v8RzOKwOmIvmQAT/kj9sCUhxZT1ZG2geew89q7cafLYgHo5
wyvmVEx09GI8flZi1gALxFwxmrEU1YaTracd6eR7MBHeO2CiNJDStdaPLTj0emRW
Ad/tQjpv7blAOlyxRdAK18lf2gL+CuNuE6bgi49wjLjLTCv6bYkbKRlCijbjOOom
GYmDVBNNWKtEPl1fRGl432Ng+Tw2P5/HYqQV8vjhG/ULg3ttidr5p7dQEuAzhV8D
7o8IFZXvxQLaP2K3TTTbiXYJT+2BhIEnvUhqw8kKBtLieYBB2PdOjnauQItCVAbJ
m6YzyjhlEGY4yfflZ42nF2Ip+s6049Lgjhil1HddzgxEDSM38SCiM1cuhn29OvyT
ElbbL2LnqryN4uhTXd74+dxzKJl3H/fuXd3ZVJ6EUTUg/ZmycKtNMVrep7BuGkGs
9ifHms2eGeZl1IGsfJOIdOrx0sHI2A2zJRAVlRdZ4WUEExkiTRQ7LTd4QvzA2EBU
opqmI2IrRt48O9mVHM6XUtFUAMbL0usZVtJ3uLFBq9B048UIqxBry/+HXxeoSm/n
Me6XoJ1gSI6SbCh8fTvt4dDh43CZeYNo5mEPuC2gjufdj2USpuUhMG0G3Rx1nPNb
BnHNf2yA4w5W8wqOYDPbLIb63imd7sHGDrUXnhbeYFoiqQoqCvdA0ftEuHoiYrO5
1d5LTzWRWuSjmKutfnEAbpY3Tp74oL2X/QT3KI0ahqSQmCRhoQwdP6bypJuLtvRW
HOtX7H9kwjwzfhjKLChWYVTVi1qIKCKkbq24E/eHNVOIjviGNanLJbtKv35A8kgW
CoY2BYUmBmGjw/IJuUI8TFrHYoaUF79Gydfajx8t8tOWUuu+wVt4YuvRTuZdGLF4
vtFbBmNckzziJX/k5AoquV/njlj1+WRzlhXC2mt3VWdA/fgkBRXPOw2eqq8Zk86I
eymvSdtQJgPA3Z8HP+TXdVqXfzEvM+1whgbvn3RJfDe3Vzsr52Pg33dgIMXdysWL
CcGrGiYne/qNj5WGXcZ9p7GHziE6GtmNoQvkWA3nDQyNUMWgCSvpiE3qnPv/dGH6
vQd+lfyCrzlFV969ZJHhrHqn9WkaqUZfLYNIrS3rtPGFUUySXhGyT7ALFK78cFDH
n1eNPJQDLbrvJ3CR6E7MK5ufs2OEyO3s2JwKE6E5plFPcv1W2RQgvvUyzTfjUZ5l
egVxya8YXhthk3LkjOROJ/V3QxZqUW/ShOfdd56LqpmDLCkcYNzmBkfAkdRKUVny
jJGXQwBqoiHKeakMPpaCGGQCmKzTFKfMhu3+rzH3tvCDFpmo89tO12hkvSpNbtxr
yva/jwpQTjh0z/lRMpLXA1l330JDS6oT8p+EmiFwVeDX4HfQesfZsPaFNGIDaqqt
vtLoWrLNHyp2MymdgfHeSuqAL7qh7l5hV2j5Fl4xDlpT8J443hc33VZaw/6nZXu7
aHY+bEtYNJ0jKtzj8YbG7HRhcd05ewLQ1LkMAQZEVdKwMjADvjzMBOBl3O4q5CSt
wF1hvABWnf27anwKa6NKxg2pE4bdulxEF8bZ/fu2tgtg/YF4V1jNp6i8LXyxf6Gj
Grjx8VZERA5Dd+vF27Ri/dabkiY/b4ZXktRp3r1FF4Ezt6l+O5Yq4uTx8dwMwGUK
vfcgawIRXH3qGd/ZiK+Ru1VJlgdMEPo/G5daoRId3w2JZX++9Ede78jjVeSxdppt
y/X+ZoUZ/po3gVZXLFY2ZWFZs2WY86ATloc5lMreakvp4qYY1iWtJKTpj2QMjrZi
Wx+7A+QUo8NNYDoupjCnmdQJ40oKCXAhCR9/WLAIw7xkqLyyeonkhhuEiKuGShww
4kuqPXV+ACrUC2U7I+pyBiylYpy6MpzRf+XN4TlaTFB2gfj1atQPQghylPfztGhW
B2hAndQ7M+X1zCMxsdw77MwRCI9uognQGJNCnQkER+3kI9oCMLAexPzQn1bys3iS
jwy5iZkSjwFyi9CEbQ3sCtp4xucUeQy+sepByoHPbH5mMUuM2qThhoVNvGL3Grkp
bFRVYnsm37RMBNkmQptJVktT5ev2Jav8Gy7LQmQ5IGpjupZQB8pnatfgoSh9n3cq
+LdRguI4lanwlktJBgUnz7vsfSNEbD8XSXkqqf4/8jUFU5F0C6SdK+PT7GOSCtgr
blEKGdItC4UZjz+Lv8dWl6RDynHNknsdQM5HOsSrFe/EA1QUspfGsPVw3Lp3U1JU
xWLU5b11xn2HyX6qz2PtM5Dvh+yUTS2kYwqAqF/ySkA142cKghp2cK1UNWi+w58h
hl0Xt2m2rajKaXCyVhUBWdcveR9s3VpCa2fi6AXpdkky84VQ9Re2L7c5iYM+KtiZ
U8A1gdlbSt8ng0DGdKrW/zRkXXgsMYl+XPZGTyGAg/8GuLUbsdlVCJy6XioQyoNw
gjbuIRouPDfldQU8w1KYq8TaDP3euaCt5X6PE0qlzLkRYpOnj4cYtiKEjardye71
Jg3D+gKP1ytqMjYr+6jkdFnYiei8h5d9Pgob1yrC15InHMsWCYxnZcqq11AMb0mV
xEJqSHlGAJf7dEo43GTfdz8KsNP94br1vz213s7gIj+RyX/klilebOsrIW+JuYTS
+nEbR5BuU0oLkEur1BZPG73HNc618iUTu2CuZr3gEGiww7y2evQG+GeZeYFqdzDn
gF8ihrl7QbnwOIV/2uDorW9lO/28H8eOaQ1U8uXjSqP9kxOhg6E+STa66Wi/mYDy
khMwkmFIzzFNHvT+QYcPyFU94vuo6JOIJfMFbWMcz1w8RTpU26CGqu5y9NrKnAwt
anbuvuJatbhXSLCpVKsiiz6BddVHUFLihF2ktgqA5aehpqemLoaxFvQPDDGLj7Lv
pzU6KPyTRLR+Km6bcapcWST819l4emghfKD8Smb/2fxArB2N1w0PDixB3cfpFbqe
6TO4CSZihFV/HUXuxA1sjAnMJLKF08rZnTFtzrn4GS+pLLH1CA0TUFJl4QarvujT
PZVVaHbtw1V9Ywfoo4mViU9+BeV2maTsfWYvTRmKYJrG/X7jsHzP98w9FpjuaHiu
NHMy5hrh3/TBIvDRmpnOb1cWpP1eAC2AZwjQjSDqktHCCaPug39gJzIdGMNnlDpi
2UEae9lWOCpccNF4vhU8mcp5ZNh626ufOVucrwoDrgqSEJvaLdtWdOC8PjTFB0ro
We/ivllHcz9++9qpoBKLxOoVq7XDl3O+cHG5XrRyJwhbXu+C45ZIItk8dAAX2vyA
jXze1ToG+W4yA3fmtCaVhQ0ZPev2GsCQRDqS/ladqmHG2mg2/WFmsQnkPivTA7jU
C+kxyDm2gkTX+ACHIra8XHodIyIBUE7+A6fxRUos1EQxPv5qNwOVH/qFS98ojfRH
oyM/Ae3SyzVCQIBWNWksPX6MHvRHyXRunrE3mJxvd9n9Qy5CFrrPyJzp9eFkrN9o
sOUVHc9uY6CL1sp96Gtjk180kDw2cXSJ+lOhWy5h0ow6B700KO5EjBFsaecXlegv
wvIJZsEgs4rytdismig5Q6713NczkNxxOByyVMg5WuTry8zMSS35Odf8vU410rDA
JMoekHomSWV+w1bgOxsHpEfRPp1tTRCcoG+PhFR6udA377N/a7nKuMJqzId8xpuZ
7ynt2wjI9UEG69Vk1tYj5tAqk987XVuf3uJXnkUPZiQv7EyUw8gGrlMcgzyLKE6B
L9PWeRhLSbvBR+hi5Q3Q+k8QIxp2gmvLJJvLOY2h8l2WSchv45Au13mHEtcw3Xps
TYAH5BCXKvIHXQNG3qwOB/X+YiDSmbYTSJdKlnQLO94Kg4JDonM7lutdsCwYlt8N
VbHAZNgoy6D3NXeKx1dThvAuU74h3zHH6odq1LJQhp1BEOhyIekbiEGhmouWf0s5
TDVIjoUtMw/N+K8tz7s7w+aNr86LNqy0pdjPK6fPm0o87dtgr05z+ezlDU1KLgIF
mcElkwZzY7OS+QZ0IsLrAjYoHdjixU+mEFUUNJ9jSAVYd+mgPNFsnJhUR2cz/W6b
aE+c//YaI1x23FpQVMi+S6m1ezDPJDccXJIcvhtD61JDVkflwB35INwPIeUN3He2
fIkJ8+sLDer1MSfC4QS+FGPyeTNU6I6oLmNutVk5gACbP2FpVyM7HQiz/u5HudvL
SJBqWLKNTCEMR/G+MRGSzz+4KVEyOxG7NHCwM6FPjzZ6/qRcobJKDdqES9gHKNOq
vo3lmBdXS/OetD0ZZLj4l5k2ljckvqMdWVWeIAnEPjaz5jx2ym1Oh/obpLirVjEG
VnwwWQtFFldZo6Wph4BrhWz88SRpZ7v6C36ZKJS6l7FZ3NA4v1pvQlfI/5raBTPG
SyuzPZIwMKnTF7ZoFBwD0lqVGf5V9cDRnU4NzZplkF5fCuGAmIubl5htsrxplWR2
TZq1rRXppUYe2jPiFHqsD62wW0mwEBnQzwLGoBqorL8yKdEe221S4jWlWETJT5Pl
kFRhrwB86mQvR09Y/XhC1wHe+3Bs6l64TSLhWdyvHgqAyolFdHLke3QWKw3xcSsB
p5b0UmrGv7vzTKCLIuH+o4hugfJaTZbhRZxod8dhvrBct47B4s/wYB9KiYtz8N/6
C26r+1+z5hK3LbQa8U0CM2tPnBnNgedNhz9f2UsfXe1X5W5j6VO01Es3qG7frbO4
VEfBUJ4S0B+T+i3QfwC2LlK4LkIIMy3l+mUjj5ovPZx0fObNgFJ7Ngl5/jZuDsKZ
TXT68Iq5s+tlpClnijbRVT+ggy93W4HWQoXjp75Ene78XC4jwFFODIG1XzpOxsiY
Z0nroWPgXJGPJQEIyt8yBGnImjLON06P8tfS83hSq3MrhfMegEH2c2HCJ0BAci/s
EmK+Vgw25BgKlVPth/AlC6J+ejMWBehr3/6CFU1QL+xf9YFngat/+3fPLXlzfCLT
Zco1h5nJWP1PbIcB+CWqddFXpKLBe/XVFTrJoIGYcK5EY7iZDww57voxDL9m4IfF
dxrNIqRSjPhlTylXbkMGSmec00UQbtqEPkl3mBwQKFO3KCmjX0wVZrhNQLY98Z+a
hphQwjHH4+Zab8GJLhu0bfgn/8CNttqCLWxk9vJlYN6nP8L6GxHaJQ53G6fhoeys
/4MsE2TOujFGC22zL8yfw7VnFqWKzwTai0jU1qz8beQsN4rA8opyyLGUyqAugA4A
DwuoeZdyD1hDgnFfdbnKR2jiHNRBxIEW+i3bJWqY06fyrNKjnS3h9qwPF9UIjv18
3QMGApoFsRTV0ej1oBJAB0vyrC3BZBsNicAxb97ZLWX5qfEec0/lHybcVvgO5h5T
0rFVnmIavkedKbX0FgqSgl5TJx61rQ+JENZ0GJanGmBOi3pOeLRazxBkbQPIs98b
R6DtbcbXQ74rc8XObacyENXFurY94rLIzl36BGoXpLoKImVUlvDi945vIHql4nMC
J0G7UmlUhw8t2YCthKhCoulmhovwSrOOCxlPgKTgzNGmGqBFGaQJCDyY7HDevfD/
SCZgohQIKhLxuvLrMS2uY1kle5kSqLYhPrcT6Z/7aJzDMjb7WGp7gz5wiWraZfle
yZyQvTm5IjtHdBt9YvfGWMewUbEBSOI1Q/7nR6kviotTJ+DxXJ3+hS3yz9ClHpZA
I5LRCTG6bBA7g9uiX4WnK7eOeBIkCIENtY4y/yOgRdr/e70Lifbb4IZPWPxlk0Gj
GZ3kquzBBnVsC8Dkb44Mi6+xVM1WbZEiCXdobV4LN6MK4UvFwnlq2+20Eb/0HvKz
EFXB3AAhITz0zb7Ogpfp2n+uCxjoRo8fsRqTKrikHcKzw9vm6avYIaz5zHEH40xw
p7YURoSLgBwaLI9JRai0W09JyZUWtGqZ908+I2o398MU99r+SGgLF8a9vSLRM+MD
XJ9O6D6NaYJDtwFbTdUnRqJoqe9SbvaKeZIT+2JrPcO7vNig3wiWL1Y95M1pyPRY
tWHkCF9wVwBE3+Bt8KS36h96pP3gjd9eW5MnfZl4rVA7wWlATFMEfP7lLtDlAiO1
D8EjIVRtBhcrlkCxCDrXlQ/l4JIi104kCryvGO+ZVg7wV/UMTaCSls8Gfg8//hUh
3M8BOxnq9H8WmdGZI7yoxRJQhi4VV+sGIMzM0YKjidnTYezcBROJu0yfSsXXDLr3
wEXjHA4867i+EANM73VBai6wBytzMd8O/9K4jBpG/ZMZkpDwUK8jS227ACxxH6ZX
JMrU4Wbp02M15oGJi5ahDU3pjRrrJG0N4X1TPzvaASh+wW7aybDpNpasIBbo8onv
4XAeSQ5kv6LgOOGYp3EobKIcUErDZBK4iBctwk069BdWhTy7KihsvJ22FRBri2Pm
w/4n7UjTUURuT9ZFMFDc6UaEHOfKmcGvP91WSItsumFhZMeQMwP4ZsoNg2exEHRr
TprPb2MgC1PkM4aWWYQ4//VZEGpU3q/pIxMLLD/YyNRePMQg7gpMCDKaOufHheWa
ixRI0FgbJEg8DcrbBZUvc9+UWEeZS9eoOitIpxqllBGvZTNBMHjmzPf9lxc5wyfV
3Xia52xaw60PnD/Hvo1An/9luXOtDvB+hDRlo+uNH6cI3VO4Mz2fTWRX7ZQV38Eg
vgL4IS/k/Tho26Ej1QNiWvghz8SccTiGpYaqUcZ6DORO3VGsdvBcsUnX/lUMtRBq
L8eVdZLtIcNehrlEoOJjPuw6UcRVygsH8sJicPD4Fgwfw/vwM0CMUYyu2nxU3Sug
0BlvbPrz0WafPGhZwOFvQSvI3on2lc0yj8dQnU0x9Wl2mK8nfTN/6sD1kBw5f4Tp
duri3uV0kBDR+GtjIA7U59Z2ue4WMKxdBQng5e42Q4e57xcXYV+7drLLvk8Dqtt6
ApC+FB3k+ONG4G48LAJFCJsqMn7T8hTrxdr35bdlVfatjt8ICGk9p5lyOt6FhMR9
lEWPRUJZ//WHyJqk58DRwaLtMobDkSTxESgiIKEgqsJsxCD2OrlM92nCKWnZbJbD
uVsJtRPvVNZLIyF87E/Y/Bk7TB1s7ocADEywaCcihMPs0Xp4yc90nHohPxCd02S3
MPweFrB9I5xQtO54GfAb1mDzvZAh5y1kWNqB6IaLREvOKQaJz53/7DorVcsAlViH
LpCD5pHRFCHnrWz0ieZ+/O5dcV4wgZjK/Sttw1/pYB7Qv9ROGmgkwx90FEUZUoWU
t0wpGBqyFTBjp0fDNf2JXHMufYD/kVOlYxt1Rvw1vf3/B219rD9QbI5/Tc5O3H46
NuILCI0miTwCHOG8rrpEK/Rb5KmMwftDZlqvaL/A9iKS9pX2RGpkLW3g4T3xD5Kc
Sk8YsdMxU0eImsKcLd4ubazxrQ50tZsDZ0zxYIwp1H6cMA3YEH6l6ouEFvQP4wMm
fgnehqsfuihkmKjYYY1Abd+eOVo5d2YnZdmrRBsAJUFOUxmHkCRRUh//rbhPZPcF
Doe28KZcePg+Q67cWz4KeXRrMEsqYbtfF6usZQcd4UBDcf/8skV7hgVztnXVFG5n
/vWR4/qdo5Y27dMKHsKSCdB+14cIL5BUrvdfFftjOap/HcnCzmGy/Z2Tma50RN+I
jX+H8LfyjwgHlIQGSGxdd0cd+7eZ3DntzkutbFnCPWuIbfeMV+FXJdQgtSvXlgqY
h9XLvx6pNSJk/Bs9MdMt1Gh7U5HwLM7kJkFtw8CCal7H11q39FReX5VwF39MkbTl
Dg2z0smcUzpXr6hXZXXd2eh+QuuacZ3kGR6pn2fczX5kGh39OY6r7PLmUY6P+BMu
noeHTXuqWFtaQ1kpHbGpervCCOSi60P8i2Nv0nQSFT02BGtaDsFpTSzamoCPuYuw
ftiWX2LZRsFuvEVJu204McOXO6gNZ1wiHhb4mwhehJAmjTC94s3tBuRu2NwN2ut/
SFJZUbW+iyexjHDpMmaNsLe8fzb98QbKy75t3Y9t+pAFdM547T/dMjd94nRF0qb1
fv+L46wr0UV3ZFtVn3BLuFiN1yw2Qfjgi3qzwVQxmQCE7f4iqNhD7+tJWhAfBEhM
IgEHb3Jdr6LbkEejFkKPFHCLbFzRVF24j1FEzK2edTZuGQWB34VIYIrzkVLrbB1u
SVOD1XmuJznkN8GBlTuvJrg9e+f3ihBFDjdN2a6RMvmm8XAnYWVf0P0PueNymvv3
4PAEXCFiCmfL0pnNszX9sqK9JmpBrKd+/5PttP6OFey7TxYJDqTmkppNTMdbFEqA
8tRCmdtRczrRbd+iB4Q7HPUj9/aRiat8yIxxsOX/saQL6rGA5vJ+Pu0NlMZvfAyv
qox4kooQUytHoh8kydJKfoXgMYeOUgD4tmckHjoKR0k5M4xaN7tUCw3vbh90UtUQ
JUixHs1jucyUvKl4npGVKLYbyR6gNBqHtpO0psGXnr0unRviHUGZqkmha198IDzE
`protect END_PROTECTED
