`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Ov1Q+nwIk7qNpFH/oRX9x8zb6jNNwA6rYuq+QBf/E6n66jH3Shyp655j8ILYNhwD
MjY54yfj7jQrI52CglMR6OFqgvzTAbSuEuBqV5LeLYUc2sL6PWgD3QpKXi/B5rby
rGtaRfrDxQQFBPu8QCsqM681zGA8f9//RpIgdonkyYiqvZgEFDyp2+feNfxRCeur
un4qpev9vl6CI1e2YWslj8nyCkQZkPOwYMgMP8L12pRTcQRwAZEHfdwzHZVMeO2s
erbX/qZgkdtYJ5iHCYXn6rzXz4Yd3VjaZpkuRRA23J75dkwkYLOkPS6gjyN743Dm
H5awJVIBBOVo20c5Jkvw6d/7cGf8LYce6dNsX3I3l8sVqljpWNe543espIKjjqjt
/PTurFoC3EK1/ujnW0uEUhp+on5dZ4w2K87aXYE+b3Wi+8bYWucE8X+KcFbiRiMZ
uSItzE/xvZy7F2EELXvVszPfEukRiFMmcrWLan3ZHlrdSYkgBqAbPF3UkVKK00mh
x1+vVZx/AB66+1fE6EpwDvh4Fv6cAmMHd7MpWnlqCiPTqH8hYCSifKS+kmk6efuY
7+YZQTkeazfIsUmuOdPvqbrUTzrkMOJFJd/m/9JCsPbIbb+W7qEBWLejBJdc+ztf
tkeVYf0L0zM6xgj6cuXX7JU2yFJL0d7h11YAQ+AhbT4RqQrRmDD5HxliKhQxiwWL
ZXA1YW+VJlFChk3v/gwvLGoTXnclwLh8TXQ47vrEt3XkDhkjG1XRDuXE4YoeDISA
g3VTngsekLhFbwYsStgSG8DIvWRVXWz9ctrMBc8ex/ABIcp4zxrg/1GQiTjbF88/
3KA7m4pyWjl9kdrOVYEesGy9f3/760SrzKGX1+uIbhswlQRb9W/yPMYUW/bi12Bd
yLNlDkr3bbhdqR1lqiq+EJqhGT7WtZkXDTAShk+W/F1D2z+Tnbm98rR4h/VutvgN
+5WtzVVEWrcQ4Lt8rU98Sg7uhmiym3OCE9Tvzth2L/nG7yovhp+jV7to5ehBZd3a
YvGltXLos7FaX0nfL2hOGBO8KOwogwi6tZOq6LoCzWYZ6Lru7ZRjNV4HeAZPd9hF
wGiJgSsgsOL+5RYI9TGDCoAaZSizb8jEUKIr8wqAAfDsdpTMSdv3rut6a6N4kQOK
fRory8+pwopHfOIOWDxdd6s7cibBBZZzc+zLOvggBtQ9mLyVrOVxvx1qSByHhyLL
NOMUUdGoc/O5GEPpOhm23ZRwhafaJsFrexrKTi0TFRH8/e0GjJf5sLhIVbGbd2kS
8tEnQasVEKIgFc3wn4CaFh709FU2vD5ONojcp/oMemLKmWF3NXYIB3kxncrbz12F
VdcC51l5n0ooQbEKg8V70k80TSWENS0Uostxh53JJ+1z+WdYEKxB0zlnBOgF6s9B
ZoPjXh3hMUUuWRII6Cx6Vfe4v3m105F4WHmk5G8Ky1caHMi22HG1wdJMyMFy+Cs0
3MiGipKpN4Buakx5UhbNpPUMWa/Q2kUxec8vPlAA3qmepg6ZPZYpm+ERxJVuPt0m
o5Rmg+xILOQMj62lpzaK4jziTkYQE6H7AKBua+/qfjk/0RNyLjB4dGmiWPoZPJfJ
OSpntMcu3V2LaEYP8R9kNCvE+AK/J2Ivj2OmRyt6cMHJRE0TtUZ4kScUvroiTgfZ
P4T/EmmSvOAXteBydzqyfLDimCPL/1oJNjSTk2ynum3Pf4VEqZGg6f0nAfnbdlgh
oBJ/4zcMnGwwLwSsyfeXULRi4fTGu6A+DtWkDcaCfA3fneQHfOyaBnDgdcd0/irP
O/kYaDwkogC6pcsccdw3Z4Z9u4OrMhg++6DA+s4fRnWk2LO18woM5hktCXmodOxO
XOItErQ3LTabKho4LiOyUZy3DMBMCBhUl9A5zFosxv9dW+l+P19rlI572slDnIPs
41ELJj4/TDuarNgu2tSwQv0KHC+CCgr+BI9B2KhDmD55TAP8mxuBqs2RUTtqIfRf
T9UvpDF+MDmSaaTE50wx28s3l+a+73oPJe58oQ25N9Qx2Mjr4ilKxZ3vw2isfyl8
Z5MOdvtwCbXJyO4QGvCnzBJuqsylh2vV1XdxZk5adpgyg/8w3MPUNHXSZrs2vs26
5gWNaqI49j8AyBJz9+LzvRlh93yKdUYu/ky/58PT3L04p/HPXbfeSYV/1wZg8KeK
TuXpEWjYBmjIm2/3Qd8SNzumxFCXP1KUbrk1fCCRA/bHPpH7cv/LqobVPyHzyQMa
qIPHCbeDBZXSNiPPc/Ywuw/eXnpkGDb1hvUmmeot2TnzD6i8Cxc96/xljkNkOLHv
14HS5bZD9mm6Iw6eyeAYoGlLZHtmmrWwzFSP5lmdouHwh3WlCtnv8Ar60SFB9XdU
vaJWR8wBfyfl+++UC/Q6o72t+mwE7TV5tVsGhTQCWXyMJYH90RKOYq7ffpvFPK67
vL+MdhfWL4gukeWB55iTFxe3LhQF5UPVni8a4Khmjbcek8tMOrc75qZcFftR+6Fj
mw8taPIgpCOBI9DJ9bgRabFTbeHZxkzZ+HxxHJId/mUzApUIyFpdtl69JLo9jzK+
OIMmkD9MvECl9QnTknsOCEjOckN+zSjqIMGPN608Gv9/gohkunm8t7buKQ9Hbga4
+UuC5NBpXmlRFOiqstB8XnMn5MlUwaHikmzgO/VD/JivDEiAa4X/cMbxZqmiB/yu
81WbVaikgvqQpp4qsHJWzYE8l3MU7nxh9/puv1ZNP/FhZqZR1ucMEpxUxfARVT67
YbUB/pzK2J5WgpIQMFZM+5/F8oeYrsJBu5YnU/a+Zu5AAD+dKxy4y+JYYViDn1Rw
21GNmF1Bdt0XOnipcilCMc/CZfWO7aiy4PXv361q4CK6gVR8AVMp7qVlg5uKlQan
G7JyhUgJTZIZLWQqWuSPgYBGiF29N2lWoSIEeCr2FlnVKUlr02Q9g2okwVmbt9O3
8fMprjBoTP51QsZnA9SVvSVC8nY1MQ7XXuafVIKpHXGmwcJGNs9SuYlK4pW60pcY
OZT5n3wTl9NdHKpScFMMFdvXwU1iRCtzBRV4cuy/uEscVBCAAykob9nRR4enuAAG
rf7vB2NakZEvF+TgYmFKToTvP0xpX6c7n9fsvZkB8VtD52xqePtDHLc19Ciwl/et
uzRV5wTCY7Yw/enNNAKlnvFzmmJqVIY2rFH11dQUqL2mbdRocJCAU5O1cHo4jswV
EJdEs57wVNWdEUdOFlE3jf14KDEqCvoTPI2Vcsfp5D8RygRX6Uq9SBmMw3g7VGbJ
4L587enfAJTh1ge5r5qmpoWCsjLEYQkZAth1yLKJ76z3SRe4+kJmTnl1Tr0tC5MO
qgwquUf4pQkH9UGf7bLPc4vfXB+2MKoD+bnYC2i5S49/6osmKnTEBspsvAdK+/cX
Jq+HBSiPaScbZoNI5zjmn5ifQIFu2gYRin8/GaX0IqqMx7KctXHMspWm0czrWkaE
0+MYKeE3KMO+cllFAkZowh6mbG5wMubO3+zlgumaSy75LHoeOb1S9ADUthqujDG6
71/b0Q3bQjF9s+GZrMU/l5XibBha/B4c/6mLEcXIUUmSwakvx8C4yn6g37JdM4EL
QiZdEAzCgPB+kWxdCZiWWI8V4w8/7AEZLzygdhkmbcZO9wMg3j7owF3F73moi77W
Mr/p63Vw4KdxeyTWBNMxcN3IsF5wdwSpts3M3AbX5fOqFGAWHvH7SKQVyYdvprdY
0kNpK/7U4oiDROE0QQpWnA==
`protect END_PROTECTED
