`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
L4JHedbfqGie+O27fP4AVt4EIPihSExc5zbyoeJ+NIObpfheek+zLTm1KMyH2asw
Ku/u9A14xClqVfw+AzA7uCpbts/VjYeCaAKDfYVwJg2EhYxxVTc2p5ggUw9ZPDKa
f5/C3/P6YuTyyaBLlK3JpaOqjzP8hD5OUNdePQ9ClLodLgbba1QSKI1EJFcS3hSO
DJkwFUHX21mEYJDplAOq+o5zDlBWKDidkj+sHkXmOO5XEdd+Bu35veP55O2Mze+I
Hv8gMEbuWKpLQlbJ5qhV8cwnsAJt5eTCTVsCS1/+MeJbKPQMCtIMOTFZwS3W8fZC
O2/Uuov08xG/V3q8r7Rya/Lp+159vsqoAoSny4ONqfX/tBSz1CMLckFG39rlcsAQ
vEsikwoFvgy/0HBwOC2ManjGQxTSBWAgSn/I5JwXIza0A4dzvTKdfHWoT83Qcl+g
MhyRpw4QNBz0om1QHkNBQ3we+8PFIafajCT84gERO0C3IdmV0uPhS0LfDsXeTe6M
ZZDtptX/t+ollNM69Mvnq7rqWjrhytLfczmvARJE6QTCNBxYbK9IJqSlcn4hmceQ
8QVI+vTPy/FgcJX9zyN+zjqmxRSmUmd2zvtTY3XuIPpBepjkPc4ZGwpGxC4ML3ah
xj/h5xBnwlvB4+zNF6sou5ci6bSndsWD4WMHRtYLKJVyg+WF1jTFTW18yRXbTwaa
I4QJzQw0YEjLChCSJ/HU0NcqfyYde9hdYdmJoZRF7IQkLiOvYU0rNagaTxxteotJ
dUXxJm6btJ7Q6mYnSGvk0BgiTmpatg3O0VCZtRocl8BP60iSz5LDS/ttINi486U1
pE7InbeK2qgTWO4etx5Pds44IyPNWRufDGL0yHXvs5D2UPvhRYSnOA4NNq1w6u2+
a7fhAixm9u95kJ5JQUd5XZodfJD+HllqW0jYJn0sw1ISrbB7Cj1t6/gs+LZhZtJV
RdeGwRqn1ueh6LqpDfDtNkW0mqitkFuCvuDnmMsu8z9/EdNUsnT24Z4rCXSHpr/l
mpr0vINy2QPdAjy3WOjFoCwKxNxKFXDMNvswk/nnulACrg7rKJYkOMsQW4ituJ7g
qzMlt7pQpcKhvzFiKp7NKNNhQb8Mqyt2zNp7sIufMA4rGuyHuMCU4DpRr8PoIdY4
cGROl9OnmQDA/Ubkj6RG6ins49rZS/zIvZ7vH+gD55kh6km0++797dna+pGeDh+G
hXPd5FT+gfUDPeQVMVr7CNit/HwBjuY/mg2F5IN45x/f0jC3JRvWkX5GNw48pWM0
ZjC2HWno0FJT9Dv3UUQ2v6MeVfUY09sbCuyv2j1OTRVLVWUoSnciHPc7AwZV4Zmg
5ABGKtaDGo1ZjFnQIh2bfIBKyb+lbs4mMXvb3Xn8Sf2XtO5P2I08k3dg4sTmc5Ia
LkqQdZ0Wc1/OAUcMKFQZFgDst48hkggnjJUsKngA/nsH8mnmNtyBECx13XInI8tw
qM5GmHGYRW8VRp29h0WygBRJtIqQlAVzm7KNo+opFp3H7stjIQ70xh/onqbRdvRm
c0rIbOA8MJCzSkjLYMnaKf3AXiNnPkhA4c+MCdOAwBpPCk4qaI+TIdfRwzvhlp6w
mBV/RphhlX6FkvUS7Clvn/yqXWpCz/ZE5o8y/P5KeaYvWroF3yPKZsG+x62WiigF
jDvF0b4SDnAeonl6a1fGprqFqUx/LMe8JoZBh4aZzmwrwiW5rLjLsPgKYS5MIIV6
VVhUjeggt+DRNuw4uEz33kcBku451vad7y8sLUvH0SdDLpE/xyEafGGKbCzD36VB
eNqhzfXG/lMQ/sJr/AkKJLDJeKvez+mcCYbluSU7OqdbZOlI0J0cKcv3w5iY2mxl
lAlPYN2p2xJHq/65xkPw//Q8STCn809/2uJRlhWX98nosg1dvlv07293SvAuZHyo
GGZ3+NUnb3eaymWqeP3KxZlXebuMVeubFdp8m0cgLwvQ7kVSYnAtOEjb6K3XL/jO
W6EBsXWGiToPVFNrk9EoRtrrGQOm0ER5xBUgZ9auJa652KvD2x2Rm0OXHiExizyK
/OqtIlC6wtSD90v0a298aHMGGYMj88AAhK5IhYVivgqIGh+1ihs0ambHKvnoMVtn
5OGyXyDGfnC4jhqbV91vLrbstJBKKD1dDAQMCNBlAe1sqAYDajUiDWnmRO0hBQLc
3E7CRdBYoQbO2MKKcfqXHZMKoTvunxwpaO3AuIq/sQjsYNvivDkPlvY44ABhY1e7
g+I++B+h41Ii6AhneOG8UFD3eRzg2EPYN8qH+cAz0oxrQmpvi7qUtnQz3tb9McE8
nGuG3NjPiuAdxvVKkJ+spuu+1apkOBL346AYoFCM82KLqD3IiIlS/tw/dhBI9NFp
tvFQly5Zv6Dog41gWjq6izs7HiR4qBHxjplk95fBpPwVvU1rMCfJimDUfznGXjkm
zDHsddfaY/9uY1lsbAAMqZPymXXIb8SkvcD//LyqNQa6zK4x3TZcXWr7aL+koDmT
RlkfWWh7gpnbMPxQUPWM8AsjZuqUnq+84CZ9i6vzRphdmpUu9v5uRra6KEOnGbEP
w0JQrq2kTOpaydq8PyQs+sWYB8oZ2AiUALjqDXGcGpzTIlhZiy7adKH9eFjN2a/i
wKyM69zSmY8slaXp1wX4QBOJ2HtkcjIER/ieFqoIksckh4cuG1QpErHXmopqs9MD
kLnjbt71eNFgg3B0Sv6fxI8hzPz4iIrGa2CVzB/4/bu8/6di2jsvi/kdDOTY8iYY
vR8RjOEsxYUa17prRqVsr94bGk7qJkZudvKXg8VnQ01sTjATYcyJc7PYuCSlmE6l
9km3IsekfX7/Rg0QRDU4WbgaD/POW0PE1BERda/+I7t80oe9CxguPQhqyENDln2P
H+YY+UjMxn9OBHmgVH0cngVXoQIjkGtaRTmrp+iFx01RwFtkgcSwqf5xtryOoIFm
ZzFL8feYzONsPRMqzG/4CvQ9YY1JzWtFuFKIo2vVyyDW5ItF55GyxgthfnurYvwE
V4H1ygBomkva0PQkelgjGsdoHC4Ympcz+laK1cloXlgG/g7D8C079By5IkyVC++U
RGog1L723qZ8zLOPhhJhQd+goN5X8gKI36b/gLbLzcx6Vo11IalktkUTWIfXS6dO
rjXBaq9VmVxfSU6UXBH947i7JIz96kqsWl70YJ53nOX8282IxAlfqs9lNOInhndb
T9kdA16N0eKAAdb+m/SVEaocdeYJSIlhJ1wtEi2wiWiDxF3S8pyXNJJFWpFqwgEw
jl4YSWkMqp2dL18pFXVbvjiLIDuWtsHjLMuw/LpfBVfYeMUX7jjYCjFy/9pq0wa+
S1ggQF5xJMKOezAkUUPrAqHbeZ++TCNaXPoXKLiJqsND8zXuGx9rMmH91X8YQPW1
sZgIiloOZ8R7wOgsqINE0r8dVcADreIbYCjR6mdMaBae/alJMDQVJ55gZ7obIsWk
+hjGnniLcgJFpgIiEYBjvMirJM+EC1U4dHmQFUNoE2dRmBt/5APN5dMejqQ2dN4m
rbsDYP7pvwCOfJiQ8WsrDwKTVevh7avrf2OLG0L1lCBLxZE4VJyRiy5JeoON0tAL
F7oxD5VNQOYY+2Iv+CmQlN05WkzY+1AwcBHNaxYLB5J9XV4D2/THi3+SvGX+/hE6
Wo/3bHcHWFN7U37UtZ56qA/hbfLSjHpPnPXvIZ78Z/qjNs/U6U2UDpy8c5dMiEbf
XXziZSoDNHILKswry6u9skqGzNxl/Egy43yFxBo7wernXJmhbovWbpFZcnMPljCt
7pKWCZcq9M8q86r9b2OfLUEcSrNF2Hnd/ygZMdVY/EwoN8xzI9kc+4lclLf3QOlZ
yYvD+uIPxwHZUCceiygoGi78AJTG5/dOGP9+AyNIDAQ9qE2S+Hlkb7keGOch9KFX
0gXkWNrcQA0PRdsxcFvL9BKQLMPifhIfs+49wrEkMzGg32/D6fnuDhh/ocdpX219
Jbxfb4fqK0uGvMZK0DUZKpr9gHM4Fiq+6c2XWJKeoUZrg/zAteBUr9VbYWEm+PCu
y9sb52lPVfVIYLnOYfbmeCz9gXiFay5j09IiIfqcKDToPMeBNNwSZDOMq/q64ZY2
HEj+bj2g8V9AIwDDTVboFNiRGLYteWSn2VnkobPxCkNQ3zED1KTkd5q8YtlyN8/T
1RLWxJ6BB0oFuCUWpd2xNJvmg5LWFbMAbQLmMR9vq6MUmRJYexwilJrHb+RPiwN6
hymRp8IMXvQhja0fZLRPUCsKRzkXp4eygzfjvbn3H4kIfoU+strbAOJGXmbBwc9v
j6WX0jWn846rrRiclGhd9AvzAU9F1GOv9RbWm92bR0JL5Fm/yJb+i4k2poLmzZ85
Kz2nOLl/2hDF5CPj2BiTofqaxbx4ulZx/uITnM7WuOR6r7UjgOd62RRpSf9lglVj
6URF3nAqBcCkk1SFWEZXFjHzfyPrwN4sqdh77z18e7zQBEdK39nCR3P0VwOhRvBl
wc246gUroBvLhaLrqx0tgVNCFq7etQCry37kIVDOOd2vNe1c1QZKvxVdEOuCxOau
pKO/wHvWYcvmi1S8Qrxs7dhP17nmZ0JvIjy6xVGE7HPlnt7sCbPkAb/3Ci52ABDn
GHrrYy6uFJhsEekWjDkbgAWRj/w9OixYU5APZtmbubxZQBk8iuHGQLWcjq7kcd3k
XZlOqApYZu4iDIdzDHHfCQ3Nhtq/m1JuuF5y2SolBfxOwkAiuDXpYnr1+qcE9Nlt
FISc0TovzS5ZawVTpEykHME2vsCmv4elta2xM5fgA3U44jOmHRFH49/XycJWd0kl
UgK6Vyz8aKUx3/E9DMuMBnYgMgzZL06JL+/oDMKo2yPV9xKUzGNr583BbQFo+FEJ
iLAFT8/kMTQIpgWYySFwzqxl8+4xdKZ2Hh58Ooew6jMAqzg7ZgutsFhQyTMyi/O3
jFg4KT7wlAbGYcw56pEwWMGU8Hdg3vqXo5p6LEBK8fPZtf4FjRxwJ3/u/gBmXRzD
wPsg7GeNg5C/pbKvj2yJNB8iE6M6iGxykuImqShpS3TxT18g5puesZb+udGkk9Jf
KBq+Ojz9eobsXm/1UoRjNLAwBiiTn/QhobR6Mjt6JUGAYlaPtk3UscxrZjA3vskk
aqr/zUIk0ghHz99mXtypTl0VglHoomp0ZQHM4bawaX3fC+W+vuMv/L9JtzkPx9v6
BDn0JSYynEcnDuaU62iobORuiXvh0a96Mg8NErsIZ7FhvBtjHl9QeySpYV+Cqrja
oF16BltbtEWE6hY7QyKCc2YFdgKuLuppEaJjnVS7Qoiy9o1QQztVT4OEUJ+O5pWL
SPLlqz8UkPgev0/W3VRWgGbHR9HsPdguOP5G2qTGlwIsDOn5ZRONju6LgAEAS7ET
BYe8wJSbn1h1vVYprvCWLEs9xYgssVB8BODrBkMbT50WvAukfrcK1YX4ECfkone7
NqYi4hoVskNsvM9K6IP9H7NQxmm/FO8LM1q4aUszvMpryDlELQ+K0Cd08CAz/7LO
2mUWaO07O1A8llhFNYIdiAwPeQqnYp7+x5b0ev9ZDOxQCfcL1fdUD9Q00tH5KqAj
ybgW2PrDpdJEoWEvNExpPEDL4Va5QGsobFZr+fuwDcZsw4Ch8LHnIGBjBtf+HsCD
XCC0LuRrMCLPlFM9ie394O4goswJqeOXLI6XH8EhFuTJVJNVHwhK51eFv/ySz8+Z
0I2UWxcs0a1A/AiT79HH3URiywLZqU77ATRd+vASVMMcH/No2WNUJ0SCDHih7Yuf
UArMUOO9+FBe/fihUykHkIf6RS7SYX0XBJR8ZxrGwUk6Z9JqsInlExXK4ZroLgtA
xnz5Zy02AKmxBGY7XkJ40wt0zo0lI7zjIY5WT6pNAaV1lbr4TpRcYvHpX56cwSTu
+GYHDpdSxg8vOWye0LhFMJ5Zt5huGwTGMIML6Y+WxBFfgzQz/IGlPfYRpVQBMOVu
rS1tJS+I8wSU3pqU00YJiRu/crNb5DNmzjVH0BXjfqLy++CAHkvz/SbODn2ksbvt
0+kbdnIySRl8Q87MgLUbpOwWOqIq4IL4SMZi4ERhaUSUhusd06vYousFeRvxjhl8
3vPN3g+P+wFOp7E9QbDAn+YLCiqJeTmFIg8Mq5xPB1lHVLbTdPFwbfwuDgBWZAuR
Ybovfc0lMF+4zLvgvMq88+Ii8l34cmp+0Gq7ZzDxQQQp7l9+qGQyf7OrlSN/EntG
sbk1dl2fXWX/0NmnPKoKdwhupHJxkRuBTORfOYUmaxSXAf8mY4HPwYNKs5r3Gnxj
98Xoc/0684TyYpPTRISJGsD2CGRGwE7r7N2r19nLSjTLP8vxbUo2VmlrHt3RaVM4
9OYQveKQcVGInHTgjaCqB4Gd85E+p0hjvwK+J9FRsG+ep5T9f7brUpfnvSCFykeY
IfuWEeUj4ZUaeuWw0NkI6dDbfmPWDUzRCfRiE/wJjAXOj99BquV8XHwvWoPWi7jQ
thTWTowJ10JdaxlhIub+TVyOlc8mQJ371LyVsY4dmr/7iDlkwuJ0mnnRc2rxxKL5
IDWipCv/zxenRV672oCZ/HByeQ0rnlmcTKGz3ea/7KKdmpFGtfz5JOOipe2ND+pW
y5ZjC6J/8W0qh9JRh5cIHstGkK3YHI+84YbHyxI8EQ0FB7t312397GAAScoYhq/M
mLsLwvh5k/lPunFBxOVo04o8PtsI1m/au4XRSuCf7YYOjE2K2Yf9kSvUjHpdsTwS
HQdDmOgzlyOAo9FdyDds2ipqFL8j0EMSOFGx3DA1bVPDKjPK+mGgh6JxWlrLSXt7
7XqzQrVv47mbz3+Xi1cMvyElWTuCX4WFsdT5oOlid4l+I1GXTDMTWk7+gF4kZbuU
S3qZpfW6o7txm2HRafXboS5cfh6WKeUvy8vqaVBQ38c/4E5H3sPZ0O+wZqoA/+zV
CQkcsmbKagVLMB8bXVWvJNZ1O7arZUUibaPVylqFbtgb4lP+DSBHX2s0d5fNDNlf
uxwnzlaO4h8XEZlpTq/J9qJBt8Vz1/+3342CbGSRdlBvQNLltbRv767xorpbxZZ1
8fHcGBH5fnHbKDoB6U1tpUdhESwa3OF4wwx5nzTqIL+vqlvlX0tJ+oc3+rIytEVe
XlXePTzTrBd1hQhNtmR6TatMySK+hrQ9NN5qcy6EWQ/qBYrzuHPc0gYYXKPBLOQ9
ScSSSHoNe5M9yG0VEW4gAuwLUailXC5P/o47T0TxxxyxXtBSWNAUZeqaxHR3kn0G
b9QQFVB/fKXUGEv3ian8GtkfbUfEjXDe2YRPFVu2cVH28aA46z3QDSLWY0RI4NxN
otkzRJPFpzCBCY5QWSEURCVTvLorqzrcpahxITmVGIaYYl9rxq1MZRdRIpZTMJxe
Gx7Kpmh3jbolhORyarjnbHm+mfgg1Kow2A5L02m958xhEe0ZPr94M/mbXfPQNbRp
2hjQSJDPcRk0J3Xfpm5WR010qJwIlhxrgB6tpwijnKvuTVH0zWsiGW7WhOJyGGdV
lZd6jSrpgYLQeYGXcfRvvdQbLArKOGg+q/gHASs5+nl3v8djbMEnL+hpUGiG/cLr
vP41ceUFty752LWtNZKpa2jY1+N+Y1NilEVz0EIWiC2neYo4pjjv+uDwuTspmcRX
zIBauzqQXTxEMbbAoP0kpBg1vvE6+8RFXeoOEEQM7uZmIg8fXnWahiCr6Ej+dv3h
WDblyMleEOcokmtPsyMsOCv/mas0+T8OS99cItej57PvNBaqcFKM3NsWWARLpMwz
S/BoFxl3U/kBd6J7zL32LPNCFQ/BTAXkNjYyuu4Bx8b+wLOJ4k+19lIHIis5q0Aa
N8FTTbzC9jebOVNmpXa1OuIywk7gXjYDvpJG4z11IIL0RjY+Iai2uH6pqICvLGwT
8sHvS0lBtwNXYaytgU8N46XCsSTYQIe6paAGYDX3LE0uiIY3Ezs+NUICLm4xgqli
BgJN5Dz5iTDsOHluBQGQaaCexfeNS4G8EhOacCld9pe0WxdgwEY5LGrKctNaHEC8
aYqFC5VikaMb1YAdxWlpFlCKi5iuO+0vbsXVQ3ZztzxOtXTNmx1n+6Snpr4Q5ccw
ahX2WcExmA9Dfm0gSKn8g11BDeTewnsnwpswObOm9ZdsA3Is7U89kqQV1YsYj+9p
fDnhlLXvU0ywqVl7mZQWngr/U7d8OS741i4TtlQhb7eWuE3I8Xu0ythcq36WEHnZ
WYmRCCyBBecC63d8UWtnbxVF3a+OqVGCeUpVt00+HfO6QVZNdlFRz82sYjoD6LmU
FmxVbToNWMC+1AhhgieDl0xLnP/uh7QMSYTQkrcD11hN/K0D1jg61dq4hiFIqyz/
6E6RDDh5n0izHbbdHqf+jR0L++s43jfHh4Cx+UAj4wN2cNE9/e/1MvEpoJA2iA2T
lXSKj3LKcsEkI4wG3fB8GK61GDBeohzen03dsaPdwSPJBRZ6qVo1JI6mTviYDa8d
kvFk107lMf5a1DAvfrwZWNPwnAjQssQD/dVMrLeJh94v37VikCik6SaHgLnNLRoL
C7Vqt8QavuRpKvwnDX09r/37DBo9ilH9NNcPOQjY8HHoh4IEkkoUGOXHL9BlYmZ5
T67smn2zizteS/ctk5V4dO5sURTo7bFZPn2Jp8f3YtEKhaqtjoM2AK3V1Sa4r2sU
QcPf0o2uPnZ2H0nHRD1qt2myU9FyVlMfQPzZWMttLPXGi4xCj9bkWkUUHK1zMJio
Ogp9agqFAXkhdYwtlBZs9n/ozDOBWN7H2jn8RNBRruwEi6TXeyfz8GUA7edigQyS
LXtQ9WZjpfdc0bGRyO1KCJ/Uyd/muqosV9sFfpthuQXeO+JNNfxeWF/YjMUB/9wt
TdUXcGKDhkfc4p+EtBpUcRtQ+UfzCV6mds3Gh1SWUg4+UCMuDpe0JXOiHtZv4ghg
kW0QnQXRBje1YNOx1p5h9dlKvI788AYsQ82VjsTQ8Qo8n4w8wCdjbwZXAuRrcmmK
6n36JLpWfpTwdEJu+UvO3DsLf3i01bHedggFGbA6mcPuNDA2Q0X4oyizF/dSEIaX
7tFDVgatbAy08jwv53lwkJfVosTNDWtYxJfAw69hEGQGtxlpti/Gbtw3Tw03QSIw
ElLCGRg7X2lGJuPcn6Hwh9uMYGq5TLpoUjlrfFk3PZRytZi7NTsMzEiuEVZX5T+/
/jW/8E5X/Ll4zmEoC5OCSl1hnl/BSXWl3RZZEiDHCz18/G+92E0u7h0ev1ARngFN
04g9ztRgVQ+6qt5eYVjAHDEr4Spw5Yidq2dc4zPNRh2ccEljytufbzXstA2eqAi1
RQ7w8Ec8xImVfziH8CsJi3JPw+dcQFdcLOi+wvCyGdDLsMwdd9JMDRzML3rM6BDE
4xemkxFCpzBWz9E79vCvdUz06jbbYeNxoogWvuM1msWXBm30d+Oc30kL4KkGs6qr
e4uiwzb/sEelBCScPcIJ6cPlDsgiYilUjh9owroo6ugXqx/BhOXNAA2JibmJMLAv
fVtsCHY5Wn7ow/jNWnqSYJT6Q16yTEzsNqrwcUAChHxU/4b3uGFA8BLhEBX197/Y
+bTV7PyhepgnLy2FPlTtqD8NdlpIZor4FfBz5fSKVgNssGbO8QmvbUpvwAzYqgMi
/bZu3PJFkctzfr7KUgVw06GWCzn7ygL/rR71MVVAWbbljJhn5yCdBksh1OCVSNtk
j1Q31qCIDo9QGd/oxg4E04pDFvIUlUga9W18NxNM9O1NpuI2m+ZcFMj430J38x5e
K/4xyrs/vsreRn9wgbSnXX3KoIVFHW1As+vR/k7GRFEQJh/HS5yhyoHiZ+pYAGD7
fHlguL6vxoOh0sYnW9Jru+exhBlHMFjvabCnz5K8gv2sKy7TlkSqimWk5gWwu1GS
WrRZH3ldFCJ80FiCsnlji/MspgEfTEJB61dLCink5Kj0+m6QF6UC523xC9sikhtp
WFiMv/rBa6kKUNHoxgCRFxyHZadqAx0O2a42lpHAqPf7r0n3ZoqO9XzBhKn0AQFu
eOw5ybyc2oV0bHthyDaIg74HJ4UlGbCSPLxfdXpC/rBWpiUpVN75arfTeS+XP1Wa
WAmYLCKOEDCuvNkhZyw7Ah1xeXaGlMv/VejSm8ng0soKz8p6ZrFr2ldfuuBpvmRE
G22UttBRtiyZKXB1AndZWKKt8ETuLLudBqkxR+GgBh/ZptbiWbEH5hCL3SDRAHkn
NLx2qcuIe9AkWUuamMWlfE9O4+k25FO0OV9aIuNKPsC7+vG/kVac/U6jG/MvyN+s
r/B/Fr49zPzKRJgVhUzUj/++eXQQ5aT5ey5ea0edjPoLj3+FqTSkYldJjgO4Ct9T
BWObKQ+Z8ocgcA6XBg483HaK25TX21CW+zbKanHzAQtDqLoUf6WVL692vXoFy89h
9BhK1wxeg2FVR5RZ8o0KHQOzK4MbAcCx/bRI59zBXYVz4cnyRQeIw8AGHLkyf5wO
RNZo2OrVTSFjGFXZC8BL/7ISD3ACNjt+2CE5dlJ65qKsv2jfcYlbofbcNHKIKnZp
JVXjYwZEDGwmSiNBtm3Yl/qM9ZKKIy41TccKyTAYNjd00gtOqtQkCJHgFQ3opnu6
GaevAzp3F/xWfcptuZDzGmLAWatjbC2ccr42DH+bmMq5of1S2EVM7OIJ77bZ3sG8
AZAFc9B9FYbh5ppkVa3xekRKujCw2kUOIOnl0c1Bj3FxWszBQmz0ZlqyLBB8UoRk
MV/AMIXhIQC/tZ9HEtsMp0j3AGtiuxWCRcRfEC1kQMDvGK7TkAGInm+MZwwAFrdJ
yr2iIgorYTva7Y3pJnhs6rhiN+ll/oz1VInvIiNn5C+7RlN7RBB4Ggcs59+1dKGX
Wfh9jP+C/e/JNGl3t8R+4N5O1/sWHMJ5DWpwRYQgfloypAh6NWqdt4L0ewCTrDV2
8Eu9Ddc398p4Pv2yshxWkhnCbbOrHTbH3C1JD8pnJefZVfz/G+ZWTw1cKZr7yhR1
IpDXa0iwBEcn6utGdoyRRI2yV7F7F7aG/9nsDZ2wLatQuEO3JHNiEYTjJI0dSk+1
zsyzLq0PpKXgiTqeTOHmOy38I2QChFfpRDfDpzHoO1ByxKvzG9Nk9CPkMIQ6Rk4T
5nZvcipuUaLq++FSmcUdnzzPLVkxxqRwx+0m+upsam3AqeU1oYVA+umKWsgDuPTL
2oSVmiwMRELbkZ58oThIbPBbYUW1jzcbS54VKPtQ+vpEyWfsaRYPsMSaDla5v6Qc
BTioGAw6pOoQMqsjlXdAS1rZsfniczd/EeJRUVT8V5StKZNolSHfrvTU3UvJBJGB
9sM68aSlmN5RCEExcgVqpkHaewdWbgQ4Tp79CNWR8MD/LcV0kubCj0H5I6ldnMTf
i26vWluLfojoGbmbmFAqkShXBMhidiGU/0XWFf7dBusGanrh4qURGtwrWEpsLHPl
pXFa45XlCGorCOBvk4OK+bV6a7/dAyR+00RhUCwebL5hnth34l50BCrnWu/cNYfY
N8DRXB91GwVUYC5sIZk8W06FX5Lf0vvvE4xsM8IGCVAO0sydmAW2VcuQSdO9Du+5
FdpQ6hbCBsYgmezNyS7F7cpz/fnfhsKMPahXR9dbnQE8NFYIq2eklAeJSETkSD9G
e0yuywt0lxTZ5hvO5/c1EGE5kzyi67vWBbYDFbyXjHEBxusMkpOedN9b4YBNlGFz
sIHDbNFn/2qK6gCMZ20Clca8mY9rCSJCE1meLCQpX/2IgeuDBUnpGe7qIoJr2TjV
5IZ3obB4su8g0mcXX9w+RJBowtHz7wUI+mIIRx/2vBGhMadPIg972NH6f/CUsyZs
0IxRbeyft25h8qkXJvSaYaI2C/Elqd2SIJorZdlZynsrjIYrMcWRJwMih3SIODPc
I6boYWYzXfdEUAff23Wml/32CGOZjbq9FTig7LVonVBkyDzn5RflYZyFTUuDk82q
w6H+O4feYI9gav741mTUYTM72Xuo+Q8IIyG+XEEtO0BexL8TcXMSO0jL9AEJoebt
V3MvNG7R78wb/HVkJpPOpCfgzQ+2jSBRS55K8Eb1mW8OoL1sXgJtngtQrhjCYtOK
0yvSAdUCOJZEYT9swvtYkormuF2RwwbIPvdV0PaLxdzhskES//MK4WyeN9n/Qk6c
f4KnIUuh55rmLTqaTL6T6ARrvLyJfLh0yTaf0oML+6mVSOGgl0k/C38Lb2fphwjS
Gx6367EjoeSjITf+HT2uVz8D6712voMitWl6DAj5exJZ2JPW0slSxDYNoSo4Igdi
OY492PtQy7qyAsvmC/JvJEkbUUSMm9AaRDyuy4+GZUpLE/ydScsAG/PTL8R26TrT
4iE71ovjys0OqFvZd00mC32SkOEq7J0URBIgP3jSMdlG0tIGCpLa0u07wyAWtU/Z
g8Xn6vB/9hJX8SKr7fRtTkGzOodZjjfxQSFcDknOiXNvv8g8Br2vUQquYNs3VWQH
is5KnVAVD/hm71wvDD9JimLkhiJMDTdVZZijs8ZOKsqReCALjKCofCMKEppGGTp0
U3LzRC7Pcvr192/JuZkh1431piygJXyLGJQlD/a/bzQ05kBQbB3FAWawBXJ9uByz
BFLO2lgBeWkc/lko1wSuns6VE9A6h+XrhzdUTNoQgyGpzloWeFiNOBK+5FPBHZ0U
R4wSZAt7b5Uo6QMBD7L9lgZEOX3oySKp4IucPLiU+Ca6TxtWMR9gz1+NFz5NGHgz
OCq++TpiSLykAkasoFyhcoYa36tlmTL26Fk+YHnPpkZ/ltrT3WjFjQRPy7PxrxGH
157huVSYrsIMfLTXOkyp6qrD/IZB/J0fTePA6S0UWfXEhqiYBwuXXtghnjbB8hCX
Y7bz+z1YfII0e6vM1lqBADVwtRh4ED108coJOuVX7CNUyLok9pxIK5jaI/nhxdvc
1nvsNxm7I2/TU2qJC8scHCPTbsa4RP0O6rpIBc9Ut32DKW8KmEgKvMFc/Fc5vLq4
VUF5zBzhnVpCicld92oUQRIyIKM5+bMD5r+U58XC1e72cf+lwb38BmBFEWiUfWYr
6WH0i12VIuimx+GMalDE+Kw+JxD8iQ8XzHUc5d1bZbdaQ0gOb/wfCscOCcrlb8Sg
crEVaDrZfsRLgs0nfiCUCEjG3oCoTOBgNmLFWlU0X9BagcDngUe3C2a5fxzYfS9r
QZyzhzJ6JYtr2H1ZhWe+pvLtSqBxP6wOME8uTGaKch7KPJo6IDv0nTvCHkBgFiZZ
64Fk051HPpecoq2nbBhQKZLzUdQGvYP2EKgNE791+IzcbLPtOp9Yf5at5b1if8W1
BgxIpPGAKWV/seapZ2sviaBLxOJ2VwtgT4+n6ktopqDnBCK4VsI77WBjKCXd5vTZ
ydPsLUT7+aa0/oQ4GylqxoDPXIRbdAWQlfZdCxQzI9M9ZSB1hsFXhfz320bNNjFh
5UpQKbtIlC3O1uTYvJ3W0797FGMbBXaNZiIzEo16+LJA7lm05wDUqLDPr8Y5Fjox
q9s2ZOvJ3UUwqxmi/naxiBG9abEWkxAQt9K3o7zwevP/pXQO44xlCArvXIytvJff
g+WjwzBg0XK84CzJhzs2RmZJYbYzrBDIFu25fN6svPnaMbCHBy3ci4GtR51TUfEr
zfPlv3TQdNGljW6EmPReAMsu51f8e3bdPfQMphEYRCAcdySv6TH6pUw7DuEta9G1
pWt7M9F8fGWIRMTh75nCMrmo4IAi5W4r03jG9txk3t4/44CbZbnKrOv6d2/YN0oO
g+NxdJCHx9fPDusPmws8IeTfMjHhRaSYw7FAEGc2RLxG0s+szZXxQXUqqbQV5jDX
C5ecn/BoB5IkgCzzwCNCgXDuARSW9rBNw1YTmSYejMkvBImu7drvwSqT28KSdeyD
VaDuHTdEgPVMgQHZSrGV8gWLeLTg3XLlSGTHkiKm4fVP0Yytb3agzB+WnG3EtsJs
GppfdRyNpBtDJ8Ih5CfnUBzVNEg6RPSP8fr1gTxDu4U87wHNZpNwtyPACL4zJGvM
QuGgZ4pw7eRQh5cGfbkxB9Z+Er3qJHNyM6RLixPGO8jmZ+NddMxk6Pwdyljp9hPB
9u09ZqV9PncgYfHkgmd5tDmoDyxzKBA/ivN/A89UUjbuvux8+wAraUExguQsn4Rg
oVNx9DZ/UAxtlu6OLfwVylD7KzRsYOHmNbr4XynLuNrpo0PFKyswKsQFFuQOb4Ei
/TQEgNqS2RJw9JyKThKSx2TQji/KYB47P4D3g+2tvzQiWU8phq1KY1Qo4d4lM3NA
rMkayw62m86f5stS01Ubcz/kkZRTAh36qZCIzl7f6nOnrPJiiVhMMR2jwBB57mXB
h4HL7Uo/diuQPyarjhIr2YRsRIBdQ/s1stqy8vwec+aiJjOc1Vs267FTKSp0iiV0
GXGNFXE6NPwubdEjmtYBOF73PjttwlejGp7us2GN3RfEu4/56Xq4kdWT5j2u9awT
QcOCTY+26cDRNn+SAEWW5kVDI5nUbKtYwlXbE9ti7B5CasMSPzIDtJSTCf2FLaxb
WrWxpvTaF4zMw1tRn2ZLnocTjZzZBd47Caty4zJliqIlkyY/TbprKEldjZZemtl2
l4iSnxAKIEfyF2IFoIYzPuPLbSCgYHtO5gWHaKdTw69EA1q1CmRA2Jq1BMyHA6ky
NgiBRyydzlG5hGMoW8k+201m6CitUBia6Eli3LW4cxNw03mqEkCY5WkAnd/1esdZ
Q3fiN2ZhyIcY6M9JB12kCHnfqwiMr7SCnG+jCrLxiool9uS0KjXY55jS0g4rFm7L
OwqLj0CX+L+nOLcuS43BGQ/8g7SMYDFJgGNOgVZKvLm0BkA+VDHw9YT1Sdy9B4k3
9cxodsg+Ck7xpslCSApHJ2PvDeoErRKG4LVoKwE8jY/D/6W7o2HcpzuCH8iJhV4n
atqx3II1ezhL8hJi3ACD9wyIuxnK45tmVnWBJQ1CN3QT6/5jFYRSYbt7bNB7j/V6
eJoBnj+P278L8GKSagIipMLO+C918Gl9/6/y6H1pwmB0+30wdubNnkgzSzfhn6Tf
aEv3iqN7bqWNBCzPF4bB2f7HiUMl1vcNjjJ51FgQizTLP94yC2vmVTDyJgKKehrp
x7OYsCb/MrQEL9CiG9WJHfXTJaEukSAR2PRpdLRRZFV7U9KWu4nKbyo8hPvoiHuW
mJzb767Uycg+HsRDMN9eImPe9pNq4zehShKzbWVkCzsmwQPd+0qHWYfGmOqe8GNn
Jwab0IsGS3whY4qg0DJlfBIOjpqJFUutfpNqR3NRHcyei1sJS+YGuvmLf8B6Swn3
1nZjn4GAzGzBncqYyIfcZX7VQ+NDadm4j1M3L0icIrjxdPmdG6Sq3lWdu0mLi4Y1
FcWCMYr81bzHgJm26A+CbYwTBnxtZ1PyFQSsMlDip6zDqI0Yc4PpppwM5fZXrQRR
3pF5cN+L/IEVPC7SCqgqeW9+HXtForkZ2CcjXrEwox/bHyjtjYxx5FNCK+V9GSKb
AOe66LM7W7Db5Dlr79hR+x46ks/jGIyQW6APPctyehpzqbFDmK6aiyU9g3S7V5Om
NEjXj00VzUvI/JNttp7t5v/+t/AuHnZl/pkElK53euixSv5sMOci+9++46N11kHw
oKhckB2bhoKW3ss6jHUvE3DgKfWcdr6uUNeNZtxu+H5SPyFLBK1JtVTTbkQ2qDpH
50OR8okHwhOGBP09qGJzEupcswaBjA0iSPhZ31O+w2uf8ruYIQkm2FEjvsozAnX1
BeA75OakjJ8gd47b2x84DFn4Oag1bNSURP2qUIQUOpsMuIzZBIh+ilWXCDmuGhQb
r2hHdBNuK2cZZJKv6yVaBOulA/YIOJi3EVtJZMYNXMuRj78kUIZg3uklUvwsptlV
iZbjf0HtEVJgTarxtx1lOXLB1mcQhzT2ctA6vJ6dDazyhHx/pTnaFgYAVGSYkg6B
kSLB7pTdiiZBKiQrt164640xqypinP9lqI3WHcdiLaiBwhV44i/XYcOHjgr9R0y0
x3B+uYJ3FLvtNRK0w8iyC0VJXoZnC3rjkFyo4IAmzxieRLTgVId8TH/OyMFxJWBN
LdZcU4fNyA/VcU0orDJcqAu4fIA3LiHeL+VimBFPMR0LZxM0/6a8A7NiYhlAkp2Z
hLiOz/J6+86la46e9Tqx2DL+0Pe/DUupsIK0Wv4Xe2UevZyHcUlytrBscWlpTFpo
z/ylmtaD4fWQB6drgQJuWUdmz2XkQ3OaIy9Yoz8YfDAqPI9GjbbkHkNbCLyUdWeW
hY4MsjhiOmYO3gK5/DvugvxsfZfmYqXsLCJE9jzCV/T47V7SBZTnoAj1kLvoLVpa
9yeqcaR8ezKUzwgNM3FmOkz7sxwDYUzotRwpb7gNJ3Ejq+HvKdCQhzsS0sdOCFf3
QzglJP40kKWHcEn+HwdTamzQz1geAWWYx9OnbIGly4cWJSMrLZtAQ24vVGbHllvO
p7c+wUoIOet6B8y1n2alrwLrlWKBLH6XFjxNzvzoAT8l7CgG9dwim3T2hhkPpAwI
9zXNMxXPvUn76ajXvaQuS8XWU2vLSQkinAdoZytV4X5pJqevB/eVvsC3jgfiKJ71
2KzdcwvRSfo3e+V8GpoUCz/D17SIxA0B2m0DMcjVv+GFXttD/ggxNG3vjc8V57oA
Mx01MkjowAIoS4yKgJqDbU5iiRXHKYXc/1gVyl/k1qgEPSzm8dyJXvHY5IBojPgP
o9G2640JTUa3M2njMo1QWFCwH9mbFlGnRo88R8f9zhVf/PyHX/eS2F85UEhiMw+g
oBD5+eYWTfDZFKYkgog+m2H4qp/D1HKf6P50j2dTw6NcowNCgTEdDLhm0Qmk1gTU
2gDSuq9vF+Z3JzUrF9SN0+nEmrKOexUax5jijxFhxB4Gu+zIFvjPgRGY99wTCa9f
MsKRtywGir/7EoIlWvtJHifYGINh4YPdnc0WTCszxEI5NpIVkwYmT+e3+10nVTl0
ubkRUTfsojuSa6rTLvQSs0KDKZPTpNynWLqjx0GNLyN1wRKLUqC1yhYl/aJfjhOm
25TtyXtzpgusFDaEuWmHZKW9gDQP16Uk+AQ0LZZC2nnzR6T7EkheMB6N09adn+12
GynKTl+fBf26DC28rFedvwB3io2GrODIX/vT56vt/0LHrtXUZPMfUSt0JNnpgZIH
/4zFFQlpCxYxJrC4cNF5Gndk+FvdF2w626icX1TRsrCsXHgakdnScV5JQ7Wg8pjq
y3VKbaiFNGNuYfIZeHoqQoxTD+JZxlH+uZbZw2YOWYEHfbNsxlySIQS9RPWHGYuv
2gOhSjADWLYTB/5zv77UnzHJQs1SJcutcEEpxbmjbiizok9gbqvMqEQIVkaPgIBp
ZrzisXCxBrqnxnVdTxLunsqWuXvw1bipMrI/euk3sawjoCmDA1juRABP1JwYdEnJ
y6+tJDdUmlJJTY8RghkqHMKiThhL/pMahKWpacgCvunnI6q7I4Mm6qRRhLauYWYQ
EtHuPtpXdDT7AEopDnhkgMPDxgLpjcbj7dcEaWd3Wd3+qT0ADeLr0NZeULLe5Xe1
1lhQZIVSRwVoQJX7gmJ3VZ21FO0Xf4XW7okvuTOkAu1Ilx1RNzRcPAsDewrOjC9S
KvALqUcuF3iPov61WGwe+GJhtQu9yGYmHofUiId6rE4jcvr7fTJns9ttMCVDOGfu
fj46hrDLgwVrqhfki7HBmhHznf0G+syG8Uo8wmPa6ChUfpsOQXjMZ/VFTwtwoxMs
FVslTub6u7mTGtGlhNWA6MazT6EEEutKRYYB/1h9wv7UeRSdofN3wckBQ37VRk+r
t60CPAh+fFy18WXMwPmpdQoTHGeSAD+BUuhJSdmomGN32oHhx7Aa/Skiig1Jzmft
pBUq0UJE6BDqqwEiASlkF+7i9swJt11ntDVAe6nGGLNJUb43xoC4OM4RMo9VI76r
jfcco/pLtLifcTK/DWgXc430oz0VZcfYEAj6k6kT/ZcK++SYslhJooFSCCIDXTdW
gvQtdjasI8k9zgh6DbQ+eHEXUnb9z9ZRScPjrG2ehHoPxQAe89NmkcMBwmZENh6X
tCBIsHWHV0Tluc8aHgj05xX5Z9eX0zMJ0RDFeenua7yrQcK+UY9ls3dnIFk3nr95
X0NSffJWUB75yHIfhDMa4kAYtWXxqH7ebYarnLAoLoW2LqcOASM6yT17bcsY1AhW
OxRbz7wZpZWzcOZz3sToi6OgECB6tbMtp1LEoqi43N4kMF43ido74s69FesvJjNm
lyMYibr8yEm4p8/Tlurw4RiR1Yv3NrO4JpZfCRKa+eN1X1+nCqw17q0dNkA1Bfqu
YIehKHUnBsbYhfc94zqJnQADyN8uhMDWG0ZyNJ7cCtB7uw5Au646Z+1EPR+TcG/H
NnxfV/GhD8l5TBsks0afvzl0VnjzCe+5CIqEQjQ1Pq4AZhK+aJ70fuTKpxGs8baQ
bmeLHDdZKUXNX4RhT3rYhTCehhoyJbPps2xEZ/A1ltUHra9I1pqADfYXwW/DKy0v
j8Kb+aJZyjxI7LFKdoICpuSLj2/MhznlYB7NOKipdFlIjtxAt07K1P1RQ6+r2gMq
48d6JESqAfUJTJQPsKTcSVcVXLai49Eodp6cG/jaFtuWZyNgoSd/Kc/yX8JLIDdI
DBdRvufl6IgZH4Pz8bo2ufs6udVpSwv/wnVWnucrmQ59wkWjNCQ1bVv5XBhNJXwn
ujTxbg/zcu4bTHiDTc1Ib/x5KbbwiAjRX5m9PkzNjDv9dikD8w1tZpu88HznnZC8
By+A/w9LuppK/JedO5H/vYRqq1A/8ybKIIAEFZBn0zvpBa0lDUqfkY8V9al5BIFZ
AMYYmJqVuAxkv0Js6YVu+Ohq0x/H2eNtn+43NsTIJYuFrYEC8XQpJzDFXFc6PW9q
PSSSQ0XCpRo25BHhToOscq8GNfD6uQq8amzbkxxdkcUb8ytIWvhSRQ8VB0x4VqJ6
pQpRHtfGhloj2Za2qf4UW5AETRs70iORd2xuibW3VQxEUsLodAuBx1UxmFlnf5jp
DDHNPUvFzdsDE+XoDcKA4YiRnxuOK10SaO85FCpAyX7xh8LTPvJy8K073BXL/TqS
CjjJQP8vfsIaMzZdjvagLIKSo7ot+oZCOxVGn3Dc+0fV4xdExaD68jp1gTetu1e4
YJN19mzHMLsg3vm4o+KI+DDQ64NCFJlc7SVH3PufxVSdkd1WvjEGiw+tbUpaOZvD
esccm1fXpoYNJAqYe31XbrzN4JkWeoUk4eb1ilBJXKyPVwcp68N5QziDgCor35tR
d9joRqhRKFPaZVsVzLs57OYkZnAS0IWuOsapcG/6RJ+q3Ya/8rMt/5d1NsmhoPQA
JgEo03Tdr4tF8K6itQvczwSJcgtDKdGM3Qgr+g3u40YtkOjA+7M09shvlYN3+lAp
260G+GpEnSMNOnGmaFH5eVGm56NfB/2jzBAxlS9WlDl0Ii8Nh8j3NTqdxX5nieHi
T7V0DJnC5xopDCtTepD2Xlsfel+5oofikxjyMSRTR9tAsZme7mT4UVpezlcX9W0G
rNPyd97eS4XwlIIbODyI6AZLOftWW4VoJq7evTKug34S8oaU8T52DUnBlDrX6B7I
e6jBySglrMPq2jHzMR7iQwSN4rjwA6NCkhofg5fIHcMiDUaTUgVnNH01w66vQ1vB
gkr5FhCfr2Nb4TnwwGIB8anPPOSAKXtkzdm3g4KD29JiW/o4T9Px/xlw5CZuYSjm
fONmkQDiXahGTjjuaNh/YL0dxyjEt02uLnAmPQ4sFJnduVe0Ct32meEpuEi9NGZz
bkXslHDshxoV0fQISTCZR3CCTLpY7/ExVOo89rFnumRJYxDJp033NcSDUxwFcfbA
KMKh65b92CWAwJtirkiXTOZ5aBx8JnQOr4wJYirZ5ObJ6SkIaHQEJl3qB37CFnpR
uXwBpAijUcxQDeUzC1m2i9BFMSQj/UdYAePvTRY3dyQw2HhW1ZPhqdKlUr+cLTKU
srsL+ChR+qaMJhWS3+yu5nF/hcTpuitxaiQgtD8/5iKuAMOaksokvzQy9d0XhrL7
1FRgAgC3PRHaCTtTACpCdW0t31MFjLiTNvqnSkNs/IWqH/+RmRfj0AkgVylyXTpv
5L2n9l5467Yux6sGGtjvkGKauOp/TfO+ZmBSMYBrKrsQUd5e2L+8gZkc1Kxve5ja
S0cFG9gvG0Tx2CxYjEEOXSIYxt+Yua3g6oEWxUEQCHpaZE8y7LXruQIklUjsIPB0
BMcxDGSXAzvPD6ePYcXc9q1DvhMl8gxyUJaDzK+fKJg5LyzBTD1dfK0S4UQeJMZM
vqOxIZHYd77C54KoJ57SxlDyhtoeJtNwEzB3O/Z1bdgXNX4sZ5wpV764ZoA8/TPr
yy6R2fSNW3YyY6mSK667bOqjUYNumI5g3cGIPDoEyJpCOHWz/mQQaqyQwLmdRdTI
lzrckmwvQjgexH0AOd349IuBodkWSuU334qlsk3W0Fosvl4LjdUly7daIAd21peW
UTqXrEYyYa/rF2ii+xbAN/wfHPkvnmONaZvM9BSq7T1nE3tEVOra4MCXqKVCS7gh
KDBKQknJzOm21gAT43VesA/tNyEcQ0tv8+eKRAXbstpkdCDu5zQlWpFSPog3n70G
5hJ4CNqbGd772V36WDlOxBucQrujOq7iOMvGipicG644c5YG5mOvAfpmtJDExxZF
ahXwT7m8Ufd5p9YMEVz4X856a6FxsMoiOa0acPKMmqaX+94rwMAyfTMRgslrB++r
nfBNbf6Q1R4reP1Y5jJduEizQkMla/QYa4CnESxhsHFeYotKyFX36xVG2Ox+a24U
s6EKR22Aq+zoTFlNMMEeT2O/ECZsr0xbHtcdPYSZUivg5ZoLMp+/1t+zUC0hVWgo
imMaiAAjOYpdga/mYkg8Tk3WfjTouZstYHcc23xeQguxwvlqPk3TyBAHrKYhnHNN
xhO0nAgZO7dBhYeuQAGJIkjNVsWzEWmvp7RxHacXf/7FBWhaSGFRXUIpobJFWEpd
Bzn5RuDJcopk2bsG6IiHBT7KqAUv3D5PyDUag+8FQFgLqpF34CFVrY9ZQC7HlcX0
QEftxbVpwbkJcR+NKeIqB1gD6kgMd5nlGMKcEoB7qcXvTPrDirVO6qyifvltqn5V
x8SGSlvjtjolGW4dqVszYsiS4WFbVHpQSXyV6VEMqORbswlZPLv4GekNHyLpP9HS
R7wmWtqEUXmrb4hA3E2OV7vx9dsG5bRT4hTmML1K2DswdbsLlg1oC0Cf2XXwjOt4
qpaWorkxLoHBtPNAOjwxP2x7FqLpn36GEYQ23BEuA1lFPnRSRst8GudlQvhRQBDy
yaPIoaE9MS2CbS3DS0lBKlOefPXk3cMCurdru4iAIUIrEkJUAkaTwA3DfATxEYRF
YqqgQraQlb9J4Bcs4vy08D4dyod1NZTlakauPCIIDp+nn85D5q/wSeqTRX5yOuTw
nrZ2rhHWffdcZ+6Ce35t8n8XRdZwkby1Hn3WdF9D2yhy9rcrS4UrKYaIpG+Pyypk
sU1UNssOU3w1D5rtA2Piyix14JzYjlcYTFZK96nPOOIKTM4cr1rVbga/hvwhy+hp
sbc0GBa2zohS3LP6f0l+k9W2hrEyOwQ4qMLa58CrWP9i8KaBQgsbps7Q1Rc25498
sQVS2szXNOm4eBJ/BZ2yrlGKUKCrYWuYpzkUhhDC5BftDn07zxDpnYjZD4+9WvEN
vXARVkCmrKCHg/xgzCztEJX1vbgqJhD+0SWD5Fi06sXayuD8Z4cX8QaaAvCiLpfP
ctWAIWSHOwNy1sKA0adPrB2WreZKXwTLvPrR8QkcztFZU+VWoklgdhAi0c80oX2c
FhgjfpL7n7+/DPe43estI0ukNZj9uvRnA2f1GAATtg6Usr/l2aWSSHpYTz/2C8+I
xSPmNF98dSqPwBIN67bg2FzEIXvozDT++YOVMySJDnJ0IwuKyQp8i3qwtGC4OuGB
oQLtV7ukGDsDTc6fPX2KiBErxih2yTL/ds0JiZkqOJBsshnl+Pe2urd8M3oNLkKb
wNjFqnsjSnk98Vw3DA4fRMScXtIj7zwsIG/D2VMXC7l0WKexsas1GxSLBnsAjaRr
2r4bnxF+ZRvuTKN0qV0124CnZ5G6ozRjXQKgPD33x1L2A9g6s48aV2bPMsXdb26l
Hgq1cY4JWiyXagGlp2s78lQxFNxE7Y5FY4lsAPUbBB9nxaGjW47VUuLgIIixi9km
q1bQr5/G3S5dBB5GYd83qKKwkzRJPNXbnAGdygO5GGtud6vR8CvfBe+7iF2vt8BS
v158Fh+IK2QDewQuGa22pXpWWPILgfJ/Hatp60DLswCe4ipLucl/G6BETOis1T4q
J9smtP502Vp7nDFhV7CNI/IRZN+3gq++epXKFqno420ol5O6hOZ2zboZxgC787MP
dGreZ4uWMoVz3SLrNSKxjDbSsJJZdbJ5LNIlnfI16oMYHShMvAMhIYIZfvvPHzfh
hnUV+PjmRpkn0JuXCevX2MianqEqe23+qUSj+eF8JiqP2MSQ78T8jQLKpDg63XQA
cICeluIYeYunV8uXwgdFwaUjA+cP2PaTzgagLVv48ieA7lTsrww87iWRdwJfXe2D
sOa7BvZl/+DlRwyhftAQzVEImlVfu6NavSAZGSJhzhzmPquCvNziMzDGqjj7OOJM
v4WflVcS0MCiIYXmPz6riuATt3wnp4zITux2qAR/RuNffpgvrQWchkvNaLL/DJlI
4Ba3EisbasT8EQzBtD6S49l08T3PVV6ZtyKgEz9TtKbcj++TnkSXqsJPPWDm5u9S
lOgWFOmKe/oJ+36KFuKr7SFo/9/AgROvFBYSrm48o9xjfkawpV+oQP4cf+Xi1k/z
Pf357Lu7iRk4dWfE5LUt78i3vwA+1CQMgfDYz/tnigI3yEspE2DzDjrD4kIjB7CH
eg0EL2gAOI9HnPYzv41K/v1WmGQZnlGR0Cu/LhSPCn5ZxCABzljE142Qhi/J4LBm
1iZTeowItAytuTgFtFkrcs77ul3NNmxRpoP3H0DhjqHvjiHAaF5Wc4hSsafuLYmf
ryfPRW0LSxbEf7gCUBO7ePeSUsY0wHPDEpfrnGbH/Q/h8NnBPcHBmbQIDBgOtIWu
caKBzdTToN+husUhwH5ni5eLwDJYgZ4LuMAulP4QPxiTG2wzmHqfgK31nNzP7kjP
3U+Rxifp6UFfmJOXttLwnGVpI3YDFu2kTpyolgGPS8Cfcs+S0CZijw+cLA63CgKX
LeJu43Ll0QoijyiZbuh5IM72YNUky/e4afUo+P4o152XcESfGq7DKUO4k5q1zeh4
mZChnluFHN5Hr/U7hgXaZuYyMcWPUS1jmjbOCugvfXnDCHuER1oMGZG3tnOsI/39
WAit022IszkECKUO/1rP/BOWhUYbz7BNg96UXGWQklWLX4SpZXNkEdgTnJmJ60n0
R06T7VegsTOwWQfYps4LWvgUA1GLWOCu/h+2diq+GGPRY8mBCxJU5lFCAVFRhB91
etochk6B949LJlz2pB5xTB6ByAAvuzCKerfRFkSu+pVQGwJ3Sd8OPHfe8vOJg6ha
LRtl+6e0A6naIPEhonhxxC9kKSuNbEW+xKsgn8eiMG9PyFFseV7fVOMLIl1Ea6Oo
EVO5LU/W6wXWr1njxMtkYRvOfse67oUwbEVxj/Oyc61hd5ErR+dH677MvJxixRH/
PXWRdpXq9o1BgFAIsbYxmrIkE4lXMioY3A4LqhXf1/0xwZj8yr+TNi9TQ4mPik42
VnwwxoIj0xOCJ+/rvL6llkC67q/5pRAgM7YlepnGg54TS5wTTIJfTIvIjOtQyCh4
+AIxBzms1VRlPPl5N7gCE161P4bK+GT66DttJ5ztBBkqG4DZuMTW3Z8vGOrrWLu+
EKEhcp74G05Md8ZaVIKK5txFcS53kmTEYoh2sxoI9Vz+l4Squh1jDxPg9OwR9HH0
Yj/JkCfpiGXYMnQBFPv1bJbTnSZjaip6JyFcjwUctvgojGcFaDZTKzyAd6TluOjr
lojLztOZbLZsiI/CJPY9LqUneldDWco6NtLJFajDlTRIU9UEPJ5zmqs9ZOQIl63i
4Bo1/K0syQcvxAnKfP64IYzsd/c8ztTgrxlM0fyyhj8wdtdc+4q8SrpuI4fRVTC/
w3SrhVfRXXK2xN/PlUAENoZE5elc/jNjkFKy0rRhKEZDODJZHiVz4KF8MDZW5a+2
QLizAS4eMaRqpPgUHW2Cgiv5XNLF0tsQxxxRQPQYkUOx+/hpCQRxBiHbryZ930Bq
LJ2TqLviEdlmlqPAZGbeXHDpvtVmcW3LSqBdY45m2trOmnbQI/UNcvuxJQNmNCzO
TeLmO4okXkIxzJBQrRmLV2rGZh/yVm5edDwZJF3lD1HO6Jzv2bEFI5VWRDlnnxIy
yFvQpfZtuTNhh6pC0y76h9G71LND8F6A8vRdJjHwKa/mBnrQBsDx63oOmw8aS2tF
Zsb6FrW6mEUEQ5oCS5t5JuQbTUQhhGOPyHJZCa71iHZZubAmflnCsJdurwtafjqu
WQKzmtiH4UlDl8v+yxcNCfW/9wej4m43sRdS+rSze8VMNfC+CyOTSs12Hol1GsJ5
Iu6i3WPnj1AnhoFQTSnBmN2XIaANQwjx5KIucg3G4JxotjL2p44Kfr43dqpySisZ
agE9A1twyqjnW+XImOIx6iIq5gTJxKIrMDcW746PloCNRT18Odl/Udut0kB/YSsK
leQB7E/vFIbfCGn30LPV8pX39Cpty/9hStfG3t7FICYFxg0fqiPL8WvpzDiAA/9U
4tpUyEvR46W0f6lp3ahfHJf6bbl+1yigPpuk4UkhFXBTtESnW8SdIVoER3ZVc3Mt
EIP2ybvCwjgLnLKzCdqF3yttblwxbU8rUlzTMNKISQXM8nJgK0oJrN9yOp35FdOL
3YAvYDEv7KBbSG1GLjQiKK15amEBjCyh0cYT0NIyZJUKRlMhNMdxz9s+c0ZFm3pu
5Ged22Ohys+yboAODHVzzVozaMFNZJ3nzqLiXU74GyPDz+X7OjZPLDxOWj0kM1PI
MEsAds16Xr2Ujq7EfWhPBGjOkktk94Q+OqFT2N2ZwCsWYnQb7n5tQMGMt4e6CGtn
ZEIjRcFUR6dYNK9SxapDB5g/e8i+aKfd/4Gpuvi3+xz7mC9VelPlfuFh2+WyQekm
n2mrbGPh7I5WDfAV4HWrh7ihGK9XHqpFOFyfeXfFr9FAoY/IHWMOo4khDMjDAmuM
Ws+ra7aeC9cLbmsuyEHnAeg8SkethcAdriZYKBixRzPJMwkmry+bEE+b+BZlPuY7
woGERgPwdfz96mcSWJ487y/ca5PQQFHU8hOf7h2JVqnR5HxEBpirmMRTw3WcXY4V
y21i6qg5TybkmFPWV+UdC/MO1wb2nMPbqIOfF/DV9e3dZxlFZC0F2Pf1RXGNAmoC
s4qvJfvIP6ijMSAt/o/MJiLJ3kubb/CgIWFfyx0BbwgSffRgV07KAdcZ4zgl1cky
ySeExoTLn5tZiYQxY1GQ7Exx3X+VWBsGFF20A3pVo+ICZDZ58uQN1inrlGPL1AKA
KoW71CV1sGd6PC8HFYfARhzhTsz/0vBLNDFCSnlyGH08XbWVgLeU2achsPhMytLN
+ky/jThsj2deZbWGxmq22twePSf9ReWQ7/JOzh69LYga0Ta/Y0/AbKbqtW7aWGu4
HF4WtmuIfpcsJBFR1PLtH7GmnfX92gmh7D6GsFNHefmAhuPJJqYTp+6wNItwPdyW
NZsYM7eMVEW7S18xO9+kZZAHjGXa9RzZAeB0kLq3uxkuiPHsTqjyADbZDxN+WtIH
iCoU0kzH8idB9RWxH3ZBiCl+pZWNFkbF1TXiAeODPggCDKfY6UM+CP5SNOBUAdEk
Q57zxF3K9+Xj5AgJ2/Jc0b1U6qexprdYz0jMtm16z2x9Yvz2AZUrLkHswln7XQ7s
oFhDlyyv2v/QXlmxiCV2TyT5e2w9SCzmI+wOsFSHOsrPM+GWERe58C4yqiHtTmRS
jex256yaKc9UFwxIApWcSnIwMUFEtLFkcu6NpmyY241+nHJSF8IrB4N+UTXjQ3gN
FxPJgP61KnYHVpLpKJMQQ/r5aWrx5qkSy5Zdv2banlTMEL3/2nh47ZA7vBxH+Qye
hdMIypxTcjwNNM3OuN9NE2W1Z1K/vjvzO4GfTnqyzPXfhY8Ko+K4qnpmLeKd1udZ
Euyw+uIbJSlZbeLTHzldmq6koRNUy4CP7Yer5UdcCBBWr5GGSiorsFXqPwVIPoeN
UikQKUxBqcWWVgIv8wcD4m8jSbqbvjyyjqmDCgWzJo0DFrj+VmgQyk6Mw73beQEr
JdjK9Ggie5wQ5XTDhKLchj4ZhUajJ1WeMQb6atc2b1j2ApEQst62/SG/q2A3yT4Z
49e3ESoZImouyAvraxi9xKg1Ul0dQQwY5tUzqZ/YKo7mH3KhN5O4SeyQI6W9UJFG
ipJQ65Um4nJewQ+BaSZnjojW75V3tRjK59GWmSRYya3sHReNrSjC9+1RACimcKD8
T5hd+NGJZJ2yNCG8e06mgnc6hniEwIEdAkS//7ibJQXLFdZrBpG/CiZMWx1G7lIj
EiSa0z/Jt57NRl1/UjwZ6yaFOG4WwLUWK7pScp+kqwT9/dsIQ8D7/IbluMUWP6KL
51zPrP9JbuibCkNsrKO9FhRVyrk7hCiyRrVwCDygVj8eyj4aImNtmLgZQUEMi/iY
gVjTJCNnLiLnD5XS8BFt3ZmaB5zLrDkvpoxKt7Y+W9NdmYGyUVwBlkhTrDPolgyk
GM54KwxQdW1yotXO0aJRu7g7s4C018nFUDMkZC9QLrtzp7opN7gUhQBJx5oM/9Cl
szgullmwjODl/HUslgLW+pCXUMQqYyavYZ3LeshPnZI4rb9voT0hcYof50yo3syW
D8pbaPn8coTdySpE0oXYjXBAR7atUrAxAmUBVhSV1xJu8heW0MAifybuqD6cgIGA
VsBpnx70/LfJfukOSWCOS+6q/vUJA673P9NUjkyw9C2gzxd3p7LumGz8acTutS1i
pXWcxyv+bBn8X+oKfjXmXmWZfxhOdyQLokDIrzC/R4UGLRV2RmIWwGWNLhGUlnz1
3PmiehclxK5zXd9a1QoTT1Q/HFYll9oA2b9T/GzCiiwqMkzxS15230wrbmYY5IS/
7KqrzK0hXPikFeW+InNj4lmug05cX/RleaqyC0h68BfkgFs6k0mwZQf1DqVM8B3M
NBH9znl8lURJHEHF0oFurM2bDDuIerLg/wKvDshbUMv5dn+bXFailgot77hL2gs9
zUs6fE2zdurM1bTa09ZBu2Oh2aC9IN5/3cUjQVTAeB2DBHWx+7fpAKy8SjAe+NcM
3bqbHJPzIV/k11bhyK7e05Zjhtd1gHmqkm5j+aAtvYJi4EIrIANtuYGAzph7rRG4
xvFYjuIPvnQ3G2UzY0yJBv6PUlVGW696hJCEB0FbE5LUz4sc7Ij9MGRuSB9DmOVE
d7vZILtKNlTwZxYD7TG1HnG623j4jekjBBk3OU+O6RYdyp1CMY5NSCLKMINqEMl8
BUyEv8mLJLJwj3sip0HBjPaaEfh8ApALZVcU1vChGrDYArZSW+9omdSjXRYAG5tX
H/xRY9ccoSsxJ+Qu5bu27yqthqYnNmQGpC5ZGahXBAOud95SJmbRjqefAD2ekwas
5kQkVmt4NynHiCepMSYRDWFyOvOxiox3zG9L4t7rYb94DqajsEC1RPCPZA3+in+h
HS4eXG6ahwAnqD9a+qSMZgv3q8pWL/NaBEYBy4/NFARJDTwpZKOVeXCewzN6KDtn
efGN1OnIy/2cdYjYJ3WhTj0UoMEls3W2dThz50VwBT8M4UtitlNoLDA37kvAjfWZ
9w+Az3+RuhSX+OBnChqLmExovLJfT95XDF2Dww+U8x3t38qFp7QhclB3ZuPLLkv5
Yy5twUcH03rk4mJQLKPGK3q2Zg8KSIHjEKHuMME6P3eB9gqfCSAubQpFmeQF+qKz
yXeP0SMiwc594rRarqb4s8pDwaOTWs0LLsPmihJsJIGjm90DwT8OSV4F9jkio/R8
E/sSKTJjNh3tDa0M3vmACm+yC1NlN22LwecEjQy547KidUtmaizGK0bBIlEXB7o2
39z38xILcUEJsYsXUAvvuxNlc4fk35pcaa5MfVScHVYXh0U+BjvzBuKuuvHJw0Cn
clXMz09DAS2KR4PeVzYhH9JXKK8ipsZ4nEwKrEq0lhJ6BtuUcszgSG6tEO0v+S9p
d9RAx7IbJ7ro7iRexEUmPNRQ87x0VmqQnps7WhTOnleew0Sxt3uuzkzkTnmpPLjm
qKyNcFwffkp+SPhOXNOyFEWPlVnEETtw44CBGCQHTBIFyo3aV25kk4j6zmvYGyzq
qw01wF/GlBBhn93nwj74QvaIafhsi5vIGBP6difT2YIe5QVNjQsbjM7xlYmQLYky
OkeSU8aQo4Sd29lPnJHmqih5BLjRoGMdGpLTv8xpehqR44msSfMxY2S/Tdr1iSIi
KZgZEq3FgD0SA0ZtRPM+iMQ+S8OTdDe6qlIg2Gwp+l4552gEuV6cr3uFh4dCse4l
vzk9fisvl28HEMx6ByWpfLtK8ElhTdrWfFRaY+/bor5FWbLu3c+m1RTXSoOYsdCy
qtszvNd2xuHmY1LoSrEjvP5E8Q1ljt7q97u0G5I4qRIxaTmPimA+28Su/qsc0nxW
5f/d+FZxYLOUiOVQdde1uDjEwM3gnZ0sNmjw/oksVAMijoJxL8sAMZmiSeLiZqLt
k9xELqnism5rXCAabpcoO9BUvpLhp8CjfYLXbxrP7SPV0tTxjrcYmNN36NuNxNZj
mz6tp/roesqSgCNYr3BIahwi7TXLu4yECH843KSknLMl6GSHAjRUYSOo/tT6q0PY
sWszCW3y9mp+4aRePFG9zrLBjY/JtrrQcVMYtrIZVO2ILTzM6ccqM8UwJfYQSZqC
yO16VK/en52hfRgdPHDLgLd6uV9qt/zi9IU3X7yPgJyC9jl8qnA91rL09b2PuoX8
TWYi4kJGaXPj+maPsc9ABaq+dTLbLyF7OvMqvm3jYFag4iSlKycqtM5tFSY71+Yv
Gl/j/wJ0lcep4ZxphHuUxqTwFAS2dEzEZ1LYHSGOVcw3nTZfhvMjIo1LF94AiIHo
CFGY96XhEsH05ZV73KfQEQVDC48Fx3RSdF1ZiJxOICTVovSH9hEvVFKih/+Rt+qg
R3F3kTw0EB4jxGCtln9nbKIUxhCzXuQy3h0wALEO0lkGzofbbnsNuu83qgKLVE05
1QHzFJn2zTlrKTDTlUdCAPNzJvybROfYqKstoJcchpnPU4P7kXpqTtkqHCYGgJdO
SMHzmqOkV/Phl4gNCTiMbVOHMp+iuHOOb4cpEeZYZFkfIk/tx2mz9awcmSd+DajL
6+J5kfvLSUIQ6MLy2yvlCL/ZMpsFTyZlJV8n11WOD5ccrj9WT+3Op+S7z/6xLMjf
98Pyo7yebVd1WTHwUZhN1Hi/T2Owy1NUfrBEslKmYyVQpFPgsFSoepd5P1sY/syT
58hwad4mrXGQ9+aQGlPd013J1C6IuUfzM8CYjJT0X7CZDLauTcnyDpIN18jiZZ0R
NGw4ww3XQVTLGhseQNgiMgeTrmfYCJYHyHED71yeq6se1ivJ5wzmj186qzqcoyZi
QNvOEyJIRjQLqx7YPzdrOYOP0IJNsmCuswXpi/q0Zh3gYBMfs2+Bktl/xlYUg6RI
ttwa1cGm664vukydRevQ+AoxDTOsszjQOOJo2HgJDv3RMHKMBBtrEHhLabsrM6Xe
ULS4hMOtgo1FCJ7xGfjqNBde15QZ8PCuiQmmVbUJnCDVJqaKSizmM0tNS5d/RDGV
aq8Pj1rv3ai8haXdnjQenP7KhrPGLvkcoj7fdx6fPYbz/qAstoSGE59usQiDFHP8
QnJ0VxHb6Vl49/T9aQOolJ6M4BPtfJQr00cL8dxizh60zH1GBr+8DIID6QWa/DkG
iFGtkZc14qlQeXqYy9f6xWHB0rhve66hFAGvJQn8zatXeS4GhlCsEu/5qm4y6gn+
2z4dHCQskupkd0CRvKrG3K2WTsDbNuT1NgLXF5XP8A3EV+acIImFVCBHvtO5Rl1y
BjWS38bi10a+JnI42BGH0a3PybFYDN0NH6LWMPG8csO5p9mlVwe+4ouqHeQGfrBr
kTRlOsfC+7q3kSyjC2i6kYzq7AO5kWJv/MRcmWGf+/4ah35omA4tRJv7sxgRW/v7
8B96DrgN67GaPN5XpAVLgHss44ByP1sws5QCcCFwBQrs32/M46EcUWcQtM5Sp/sm
grff4SldF+qK9KjQGhR+Ygjb4yNYIg4De+2n71MDhTW3uvoK47GnX4L0Gt3joR81
1FZfYj65l/aDydi4nGULsg0C20uQmC0wVRPKN8dwGkXwqgS9CEMVgllhghy8xKI7
+UcH0NUsofAlPKXhR8JP293bk59hcymeud5k7fEL+BTpOdGIweP5CGMH+cbVzZaD
louhWDXer3kR5B5KeUstp13E3eEGfIuuSwolU13rbA9h0JXOrEljcbaA0gEfa+HR
AJtCink4LfJZ5uQTgK7ERfJbkMScltdJTCo+Tbgpp1Zi2cefj0rCBN0BIxSOLmau
wZuJdN/uKCbkfVsfJYJrnzLWht0G4mAlE/WVE9OocNtjAkLZ8G/mk/CmKZggFBvR
mrmdCQJ0uc2dA/3po9RN+PSV0YtYHkzDkotRyn9h+xGsTOsKx9sXnsDHcsyI76Uq
iERBe4Cc/T7Y5J1BFHHbPQ+rgc3ihDBk+1hS27SQ7cbxEJb0nxWJ0cArzjzCRg7D
MoaMAjPJbn9KPW3xddE91yDNLI7CUeMoUdGHEfzvMcXBBRZANq1NM7SD1OWcW8RI
BzYWhaA/f+qZIAlR69bHQr+vNKeo97LeH5NFE4IOkh30Dd/Tl7MU9ijXfWA1Hxpi
PYyIr3tQPYTIxC1djvJyIdXElgV8AAf1Pjqj5yygiFJd1vgi2HpCjKdN7xzrwlFq
N4R6A0opyx2f9BkFP8vO+JuMpyAF3remjnKQZIKxrtYQk3acouD/E6wfxk8Kin53
AFgfLK0qhCv38uGxCIh68v8raeHMETfjGnObyLD40lWBN3y9uP52NeiNCk/W3eJd
Vb4UcZJU0YR+1/iPjYQax+A6KlqloxWK/JgfWkN+t3Dozy9AiFxVENTMPDEuN/hR
o6QB6dvduTP7hE9PzQjpwsDtLZjagGikxYcetl/DvzmS9KUQU5GMmqaqBEn4mTAS
JH7lmhAKQVx01bj0vVzffF5CRHXw0XhD1jAw/JEwPFk4w91hMX9JQqNtqZC8erI8
nVXNCAGP6WBST/DYqZHPbAjRSgavzpWKZxtizHScbIKonDvor+yPNh8tzxVFztwm
DV0IXjLOgwHVYJ1bON21ZdVVsSCqgdRrcfOK2H0kG74ObBKEagAC3E5KE5b6csH1
I0zNNBf2HBlrDU8Qs98iu3e6PBRh6uo1BHjzMpvI1HOgjENuT9cxE97PmP9m/yzP
P2YUWogd2xkjukFSJq2Yil4c7JEvNWB2IpZ8fYm4czlJ5o8HttD/j8NOqpsJQjXG
dbvK9lqXRm7KH4VDJy0zPgBRB8JC/tBg7DBVE4hT1Q+003gRcs/hh8GUSpZlyCNz
7bvSfcd8o3pKJOyRh6JCly0AXwmW92rSt7O8Y6x7+SydXaVDP7+xrht27dk5JDHw
vLRmoX6ttXUspAETZ3PB/6L9obenJANCq+rbz1JB4PCftrAnDaEck9SCoo/5DYWd
DQB1mucyNeE3i1CKdit9nqzXzyHgETfpYARddJZ59+cfmGIl0P+QF2bOB2px5esT
yvQUdAQ+nrTYjxJRVJjKMEqZWQC0OcE6HRwPXNmhyBkpKD9NyaZ+xnGFNL4Z/z6f
avjt520r++pxhDh1agF9KlrEHyxC+BeFgzn9tuhg4y32RgtbmL8+LkPq6Fug2soW
Mtqyri1k8WEIC6MbP4//jNsnd7nfqbxYmgFC4b9FzVYdewqfI5Ff1jgLEbpP1gzT
zb5ZyUiR//FsT40vwndYjoRZ+sUElqPRzBcbwueCC3PtDjXSHTZgND4I3qwF0hn2
avc05gUb1GNEZhCZ0lgqTcJ9Mznf0j38qH4XKQafl04tyTyKYQkgbmSWXzHOAoq+
qpMnRKACNWPJ+K6soroLxOzz2l2vTb12BYMFygZr02tFYDB5BdWlDFsN1fP9QLle
KCatayEt1c4uWkPzFfnkbxM4RCVduyHXlRQqfG0Klgs4nrocc56oidtq9OhCv3Lk
g/bEdHVoiCtQxrtBecYh4cHkZDNNObtuGHAJ0IL6U/8ZyMTDLtTeq1u5NhuYjpE9
HakzO/1yy1fWvRCzf9lwKRPvYUZqbkgFZXoLEgxRj1Qb2mIVn6mC9YhIAaTY0JJ2
U6ub3iBaakxa22N7E3s322rFBncqg5k/RKUmIuUaIXWr3cL36Xrrz3dDHFbOkw7v
W+OwCONkRpjDU1ksQ5DSt2N/MOQGeKLd2b7v4rD/JzqAkwCkXhLS06s/0ZKn5TRw
4dMPgwkJPyMXmcfsaGAkblFYaki5sEWiceNDlF6xcwwrSgT1SnQP3TFoV/2WmG40
zB7Oeb02keenCK05aXVt3rEr2WmvZ6TA66y+LNm3xkYAwgjbEKQKUPEi10VN9n6w
8FgJgQin4W/bixerCYflXg15DEmpSG0ZxXK/ENdiyvyWgAI3Ti0lF2JwTHWtyFpO
7f8Bw93/rFz68VVU2O4GdNF+8QL0qyf0eWXjpu196a8rt14xDwJAEfEd5Q7s8x3/
XalP++ol5DSDedPH/kNwAt2y1X6FdJ5lM8MbH+bPbZ9R1YnT2oYJoX9BxUAexq0V
XZO4Jr3MyY4sRQYJIxkhJS21JUTcWuBAtRE2fmMwyZq4YyhhEgofujBboK2hWPUt
YVKZrTv4txOuT+uqm98i55OxP+rA7k+3amozc0bJO+P9YHT7TIWrfo0ClulLVQXe
qEsWwE+6S+8ZpVH/H4NX3j0x1wNk3HYfIbvHfQGvl8BZhPvsx94LM5J9sPcZQjnn
YfX8N0HG3HXYHBNn7rQ24QWtslN35A296Wsseoq6vncQPkxtZQyDr6WNZQYIKQEP
tDlujIghaJcDALLN5yIsfPwnw/ZKpsmjk48MBlG5wVRxkV8qQs2XfB93RQ7l0ErF
rBYBGw8R8jZ1QL4rhLckM1BuSrUg4ZGXi9Ycb7nF6MUT0QfFr+xCKZZqWp1rGGJF
1r+TVQhtjRPmR/zKNeQKiXjf+ACNWP18spItiQ0qwV3MKmjFr39TVLK0XfuX+2wZ
kcUgjtakoan0il/6yA1LXLIdgWsB4NDH571DvKyH1gp0BeV3Rov6qMBwywcTxURt
QGtDXg8dH4O7ocSo4pYNt+G2XeMKaeOvtJZ8bhCU0lG2bP0xa32XhWYf3Qzh0BF4
ggyuqIEOycHsUjUIpnC51UbpdxYbpmj6TapPlk12VKWwx5WXB6MOEU+hkuyK+aqh
pp+RsVbLOiS9sV1I90baPgKYI0kXzZOS2BROkYw7abzsQVy9B//lu0ILLfHIWJ7P
LJbTr68VbRwZqLjG0ilny5/eFycHxh1wAZZZlKi2OaOrmK2xa59nReUM5BOdzXwA
uhy36S1vAEJaAWiKwQlQZ9T2u7zWNntPI+D52HfoFjeygdIRnrjDEb8a1Kjeb3qC
adWKYuBrkKOw2OFHfVL+O7loib7nGX+Zy4p+4U9J4rZC8A+JlXmvQr6iWcjAyJZF
HTeQ6uZeenldBYjlLgGVhmw+EmNwCNUzy6mHt2qWKMDMXYE0tIOFBuc14eMxb0f0
9XgdWXh9KCsmAM54vKOTQ5wk0iXDOuGVOYldXHBxaFP6Mv/teYBVsKmJRowxQSms
tuo75nUGssYNgK1eYvvvhTyyHlOO7E84Cn/uUrFgnQboAt2fM4UDJ5EYAJ+GK9Rd
MUKNicaq/j0xlEegYmjYiYjrJgNnWIyVIUp1WSOpPgq0nOlb43NIu9Gz1Q19ser8
gicIa15/MEgRFcAlR7+tPbUDR+7UkY/HY5TkgAOJ93NDHb78ipwEVwqPRIK9WJFJ
/OstK3d+WzyIDsbl04Hyc29EcD47L+eR8yiqTj5Y2uMlepvVJL6JEEcmqQ9AMCsC
S0c97PiZ1qbEyoi38p2uqklnQ1oVjWUbDnou0v4P1Ro3l5XZLzt3A0zZnJycWeV+
HUPDWpNroM14GdMtHnDtvHLmVtdqCBduS75JuYeMfANG6HtrJcjcvXeWL41qx3G0
QZ7xatmcc8vtfXAHpVZXFH+a86kv2QYR9StEUXublRbxVB/RqGBZFco02RqZQFLr
yADgE94wJTe229681SvLLE8GFG3SgSRoAQymkCRdUPJ0B8KIgrsa9DyXIGz4VZOc
xqLEp2XykpzMlcUSRT0DCT60l3ZUzl292HRelkbAnpx4vWkXi5E2oKteX2vrODCy
8VU9BJaqvUlQAKdeEnZlDxxsSCU8C9jI1ohDC4mGYNbs/qmDogUQVjbO75BXJFwN
LJlMwYxFG58R8f/rAjeOU1/EqlKP1jWHNKgsMthLzrkaq3QMsnIEDVZZmZM3GZ8h
7YUNN/zxouPaRZ05e8joMOK4QRXLr7kBJ6mkcZx7KHQ7qEODfAIbIPExZqjoiJLF
WldJeoQJ7Wojau+YGjtn7/sShD2OhIEcQoIRDBCVDwoF0HCLoXSkhWGtbvZTJT75
ydbu8Fb0bpRgPyYHoxTt/FsVz/QAJYq34VwPTFOlAsdL7c+HjlCgPDNG7NLXSGpb
oox9gJhKebFdq293MR5rOL9+oNWsB3NymmUFFz6oCrtMQE0DdShpwypIbotNXyCt
Fakygh9Jmw+uKq2aQfwFRar6iHQaCMSVxPq/TXdRE/RgVa0winNgHA3jNBcFq0iP
Nx2YMGAUGF4wXQAdCqQrzeWikSGzdcKLcMw0Uns4+l+mKI6ghNLy6rU3mKkzRvr7
u2ykR9WQGDVeMRn672glfmUPbP9KOxKCL+ZuBQLqjgB2XdeNG3BBLFcCOXaUTeZL
/al+63R5STVrEweK/qb7BY5ESkDUdKF2Iyye8FRWGEmW+7Ab+7rvPD9I/djyeIr3
uS6ER9HcKXGBqbPEbKiV81yZgFZ8xmqwE7R4emdm/z/lT4K7HPeafLmtnqDJS8qs
PwqM4tgWuhdEkk/muBq8mqjfYje47FL8R266sspBaT7L7y5nVb2SnzM/8IkXp8F6
AWyDeLDClPO6vArBAcxMsMUVcn3cIqBVQKrc0pCuk/7SuR/9jJ5tkbkzI6GuAxvg
IsZlATG9tS3gYsNlhe9DgvMzXG4Qxm9hdaowD5cBCa3lW6u7FWC7pQlg+iQ+Lu6X
p+Jw3yF3LJL2Pidsl6WMQPDIsRmY2aYkZcgv1+WEP0Ge9Cf8NrSI7mffZBondDOh
uUSrgpcClcZgwEXFX6GBTUwvHCVs4ilUgeI3N1Q1KuboyVS/VOMWRr/GNsTb5GXC
meVRM2sd0JALhqWYHzOH2tuKU7VwjWGbHurdDBBlcuk5PH5sLhAVfwwv6knF9jgc
fndbx9FQLPTmZh6ihN0c5aWOOOhpoS7z1Mcf5Pa8l+F1Q+xJnEkUDVYD7smdwVRZ
`protect END_PROTECTED
