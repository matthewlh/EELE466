`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
lq4yIdKWahwS+GHmBIbcofB7iXCmPFY2fdgrJQs7PDthnXZ88q0E3OuFa+VzSs93
Ce0/s9hpihaPLXCX15MyoyQYQQ+N5oMWku+zL7xoskpyirvcZPZKUvGleUOx4BKA
Jsg+0Odm604VkpJqLk/1s47pff0UyX6JHywLarXiOSbBC+pMa0D6js15uwb8g/+2
t6prHDpwSKLSA0DQGeY8vPP1Ki6PPE75weRHlLqP5S8ZeOncRPk4vod/aIzjvKDt
72X/q/Fcoj2h/RK/AkL44ADjb+6FPs1tTbglayml9t92Mw2sYGN1wUmpkaNa4smx
PdaWtSew0IMIgy2aBDtzmf1Q+lE0Gk/Utqfg8NDT45nwOJKFvNOv1at5JUGE/UxC
NXBgHrMrIIPIBuEs2i6W/ZNokyuBBK5ntgjKOvs9Ccz1E0TSeGxvJD3rxuyFbUV+
sao7mKLN55GqIS/kXbHYzGvliTSwBqb7c2XdNcOgqOpL1DOyl6gDV9TEW046wt0y
VLeVhpP9svLxAEpFbx14OPmO3sknmbJodL/zeVmRWvPJN9j1q+h0LNTxJmVvdPt1
r0GFinTwokVo/6B/3RQqQJK+nGKlD0ejuwm+x0GpTIVNA4r2cPFJjF5Os/F8WD0n
la24mQ19VoR2ij82tsl2HchJiL3VYP7RQz0D30rXgidNq7Lcw+7boEO/Qbi3vjll
sIUljEYfyL4ttmvxlwx4Epit7sIiJnTyogaqtuvaQAk38kNt9WxO1nILWp/yNkN7
cr4Jp0SOOVUVFFKa9WXAiUB4CZbVUbhpJXo59u52uMnRoQLxo2CDnUj84Boxi2RE
vFdndeC+Rb6mYegWwkV0cQ8RwsofwJ+1kDxb3V97G2pQl9uaZ5m9AF7Sg6Zg1TPn
+Ibu2i2Ksfoi4EYfkit+vzxhHZ0QndP1zDVO/zl6qgHneP/KNwZJylazxIwzQQum
txFC7HKKzAKssOIsKfUcvm5+gH0MJUUNN4iY5yFDsA3D+JdDAb038OhcGQ8xZI1O
lYXz3aRn/jO/KmZbUdYpA2SLIbP5XL1eSLtzyfbhfL7XSL7IZsDn8UYDC9nk1PyU
6Eyonq4UxR6IhR0/7ZoUPi01PSgOd4m3kb/tnTbvxrE5tFgOOQsISmFy8zysbzWX
8EUmIzW1j9tpxip/qcPHSkSFb3q3df5F32WRrvHW0XFc7yPufZlKYdjGhAGIfICx
s5Hp1IC1fOrG6uXh5Ja0PQB0k2TuRtB6ZdHqFv5JPSjOfN/Dy2up/86NbtJq8ap0
PBDx3mA5/WxBMJ7JPW0sDgI8jAG6V292qjlBBR0RhwFxJ+TvyLm7mDbqEQT+ehiI
G3BEp1avxIBt2nqpVXPUSFXbqUCUaogDAfTTM2Mc52t5cG2XGPdM3HLA/4tq75uH
SXw1Qca/lw721ZWHLpJDaTK7jFh2f0OnFmGhgFi9XVBNOH39TQKUseignzNh269S
Zx+z5ASSCeJ5cNc1nigSASUujk4oPT6eY90ytb4ZbHUIpWVB0KrwMpTNT49UfRJQ
yX8GgdvtinBPycaXkr1U+WV6oNoUUX4lgU8Y9i78IzyNrBnb1eTcNoiiPURu2v2a
WWw687+n2AQdvb0Wst1V+HogJc9b+J3wq6UosS4z/84ZFbJeOopNyHlNydonrPxU
KoSUWAMphraNcQwo+SDd7M9616vMmatMvvKzbavtoOu0PnKsV/RjrwIEVrS6EBj6
g7BkSHAN8L9Sr1XaqSdb9Epq41nFe1QNava79+mFSfb6F9xYmj1QhNOEwEs4UA9w
DpSe5t+Cms4uelcBzLo8kXiBFTFZO/AfPr7yz0Uhvt2PN7eebvnf51gopbuRgD8H
ZoJFXSvKmIErO3g9LvS8e4HSTEee8C4yuzQ8X1QwvrqxU9dQjUnMTsLeFjyQ8mMe
sYhESZ4QIaYB1nY1R3UJjdxfVBmaCHkZsVxgvDNTagVjuXWm0SSfHWUrqRtbRyv/
xghSk4m6FsODMcMtRyjRggnfHC2pHtI3CWaS/2oTzk6gC2TWYrmBZnC9f/TP5HYU
/VjGGrFUs4T3dsJ00dFob5ul28TaWOEzeeqfZfxindYo9OWwdcM1s+vIR00WMc26
hxQ7e8taEz5b6WpofshPXftmUbYcNzpMv/pvgBqBSO27xDr9DH9ZhpcLsRCzNTEn
DMOEmfHj21rQ8La02r5CofHHedFLOwExluDI4HB0kSz0wUnouZw4bambzqAxaNZL
m4qaKJmSoRVAwGr51Vdy2A+s5mWn+7UpT0NslC0GUWmfzRZbB7vwX90XOeS+t1sD
aD+/vJ8qAQfh7DIaoopGh2krKlccyHJO7AVcjxtzkuFKg9TqdldoT99FcyVOZKHb
WBhSHyHUGbg6Uk5k679GrOy2DtYJQUNKiPryCycGcH7c8Y9ki2xwt6DgODkXTUUD
psGnZv0Wg5xNG5Mq1q+umQhT1jgSYviWJZIpMo5efH3M/W7WKP3JH8FqNz9CHz2k
tO0dDLVj0NY7MYKxYGFsL/wXU2pFjPIzL2VRjbRrdFDoP4yVGSSOcu4fJjfS+mmK
5guHXt8FUjAD/a4cHNCtTVrkfUZ0biQeYlRHptfTQMVAM5NOs1KZZxmb21JWRiyr
4wAaO/2CRgKz3GIiu0RAihpRxR3VOzMPo7XC9bUZkIuX+KlmK7cZd/7uPuztE/tY
RD/iCBIfyWceeMviRQaRFNOsrL05RiSQvjp68Fjh+kOu/nE9G1KgVFAsMvIvnq7N
s9fvNkp8JrViWsXCBXS7vFKvTHJfifjTMdFaGJ19uagK45BsDHk+lixBgf4VmTT0
rt53iRqLxjGuBwTb1K5iv7oBUDxlLuWIPzIZguwgaoUSryJYxnns9EIQP5MZD68V
PTHd7U+Ds/T+1CNmSpPlHNOv0b9d+4np/z9/m6fWk4tVF+TW4B0Rb95/x2MbOm/S
14FosnY26cxkXtjNq41CULevQdqfC4iZNWt8aSrtuquB2+e3IQBy0dZNHduA2hPX
Yj0CWREIZfjHzKB+ucl0D3xrf2/XSoGFp/VIkZCH1jlL0OSqOTLlL8ajZnPtxX7o
hMnuf337PRo6UcfmLmpmL+H51eLjMcKv7HhB1DvPPtme656AbQejf1JceIss1tQc
toQL4zM9O9J/swRxDnrdyxomz5OjqNGoKgd9cBfa3LJiQ9wCVuYh/ueqqMwGoJLC
Tv4V6F+pDf9TzAHXJIH4dizhhNkhGq9+GkBxbCpHX2OpiXEsQfzOeOo4aiMgIDOz
CL03VcyadP8bO4mYzmdwvxvEUygxrSLwbgp0wlvk+9VVKyXsl7+8fF/j/m8KLyLt
p1I2tmi8UbT9CsLSrQ4uY1sANUhPzj3r5JoHWh6F7M/rJorlaXoaZiDXdworUCzJ
8FGdejHVBKj2L0VJXlqJ6vwYUg8rurtYos+7XSTQ5YgkIQOkoYZ2TJ9pZW0CtyKE
1J5U3ZJfUobIrBAYAWVMDWjbgjCl4DccTuOuDwaAIw/dybr0wqJLQ9gCl/oVAjGN
2c+aetAOxMqp9ENqnl5n4Ee9TBHe43s4BvmCRkZSCTU5pSy1UhsAt+PJ1eFaDOWV
eiNg2yhmC5ZaisBAFSG4y6IYetk2k/RWZwo52T7cesFM6EfKOkPRUHh2sV968P0P
QHrBXrYqFEpvVgT+wfWGXM1eu9bog3M/IvJTrWGyMNialjNW8ZW+S26GmoJiwxNK
mgTi9cdvbH7Kwb9Hn+XJF0s+1a1C6AameMVzZiq6O755nQH43YT+v4ijH9CveSFQ
aM4zg3Idk9z4Ew3FA8ksnEVwQ+HVve+tV1dX6dy6bePZlDkYWzaXhjKGyXPXqI3H
oPczoYmYM6jw2odnPrzoT3jz5TSKkzQVThmPUR2o1e2r1zwf03ZcfRyTtHq5PPyU
+HGx90L7LTWf8DhdnL0Au6hDLhmJ7bjMi1e7D7wCZ+umX3PKpzvAaTEBEg/6rYbM
QX3eVlKuvHXOOSxbtkIZnIvD4Px12nRNfiGz3NBaKqRZRX3v2J1x2lwXSuJSXpDO
wAtSTYDh3Uv+hP+9k5cQxvA/0jMHg50ZgxFZtORXBaNWQannl1bIH7GFDEUKqe/8
OyfVqd3EQSY76+1X9H940txLBhDjlLmorLWdTURnSuQBps08ykHd1+9ubcygNE1S
uBvkzpXjRpdnDgULU+/f8QOh2nfQtQ8naCfnM6/Gu18ZBHw1UOpYUm1ohOK9QD9O
2J5g0DxBjsPtSamTxwhimXVEk1EAv7vwhzHtNBbUKUUiwKMYvFSBTAJ86RNqhv/r
pk/hpIVarOsmaZ4Y0UjZvByUWemBB+AzcAvm5kVWQd2NKysMq/iwnDmlgG14ol8a
UDVBWiPlNt34Ikw6KnhFR5UzUiAflnkq4ah/YvXjQ4jfdvmg1siLWzsZG9SHmdXE
6V4Te3JduFPmii1UFzma2V22KA5Rsc952anneFve2QieRfRgHhQKgiHAhyTvn/3i
SK/skE5BzpFvMd2067sTpj3xa+TtD5ZDpVHf0Wqzv/mEtkJbgQw0hEyZ8gWH5b+u
L5dXbpHFAr2xBtXfDQhlEA==
`protect END_PROTECTED
