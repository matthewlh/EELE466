`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
yPp2jAUykiLdA7O+/pR6d8binkO6uUC0SucJdOv7IS91xiNa4kBcL2ffgmI5UkBs
CWYczuPkQTy5x+S+WJiIBOWoKxrIYZYrXLcFzXTzvjqkPRRLzdLxnwTx5JPWFN2J
CWhtAP+II4QsFGvwVLuNZtML3g+wm8dmOtne3Yf6/yI2Bk1NjM9S9PgIlnjBgU9d
Eot9J3j0Z8qNQhZL6Y8FtmfGil+MCks44OMS9Nmh/U9wusphCvr1trWG038j8H1K
b6Y709IqXKfTyXCC2HAK/4K/TSGELHtaascsWM6tzT4AVQLy255t6CYuW9KdpbrX
eYIwiWaeVcVh7KLNanc0ak0EUpagKv1MGt5/0s9yUTUYIunt+1wlr+282FwB2kiU
X53eJq17BP7AeGNK9Q+87Op5cIeHY52sO7ZV7kkJu8Wyf9bbPDo0fylBVmg5sODi
K+tderf9zQN8mOWWNt0df5ZdXM5HxlyQ+DWo65DE5s1l2vUIZNIj4A99vyeoVRgc
duM5hyt8ToLTXJGUlyY59xIF+8muTI3M86GCfDRGi0wzsYBdhNJ3hW4kYuL/J27K
gemTPzaUwSIR9pQ5+u5KzuI1bAUtvh2rj9GelBUx6zUwywQ9KklyChnrUWCZ75t5
3x6O76yENTyWYf8/LlpKh3/kl6C4qtiqkpAv7Il6YXA94HTcJ6Qzvm+KpsPSwlM4
YLejH3qBJ1l9xR/r/hxuLtuavrqwQpWgIDkoUwhwiT7ELUIf4pnAG/Wh9Q6/NG3o
ZW63/sWOqHOZnHlXA8GgOZ/gHPBYGqbpLLoqXs3TaqnMWi66PJC3IBedtD2r7kEg
y2XIXmRFHRPeg3CssAD2KMh4voWePliek3a83a2q76DhMco4rax+N7kv0PS73R36
HZTZF1Dw0r1avj2k4q/xy67bHWZblg2Gf4O743Ox01DELXiUj03oKHsXm1p7xaPX
Gdy6Av7RYtvx+5lj+ZV8GAU1GhlcocKebrQz9nLVS3rXcpLvSYMlhye3Uonrlvk5
djED4S2t2bvyzHFAQCi4qnhDWR+/JQTpl9dUGzzKFmFu4k1PFdU1RnRghgklIXUZ
w0LMtomDTn66geM1yHzaGxY+66Og5Kyyxa97lTzH+QLTXGy8qTrL8sC/4oqwXXMi
bw/v8RmvHEYEAu2GFxTKIf3VYOeW0BBh2Fw6dBOPqo33JWgNq9HYpsti8x4kE7/V
XT0TYOFaY6wFZg6YoCpMNgye7Ua/zVm/L7iEPZaLfOfbY71Rf1GStDcWwMnYieAF
RE4BCNgh4QIbsiOmKi8Tjds+JF3IuJuv6ymkNIv6fdwNJpwRXEwvezK7B1faahC+
diV66EULTZiPQ7QyIlb/ZOq4WZxmadST1CSn8PPEsjWjhcKbmZKk0D3/j6srV70O
B45EtoCp5B9Ua95/pzWccbmZrqTggYSS4WQVsFqcBLgrXdcRU6a6AwBeEsWQXOnv
s13zgGfHF5grPQLKmj0nNKwmxROM679Kj8Dz/UGJHCyWH3lriY98amw3hOc8rD1b
FPiCzoDtTu0jxHv83Fhm1/U/O0Q4VFdIwjHsg16Ikood/5z5unMtmVxKFX1K1WKR
eac6kf5nK2zAv0ToRAG4GyN3rwkthPftwSK1NQMWoH2udNdNwqnX61Xlz7k7RiIB
i6amVdjBGKXxPXYHYKh/OORip6jrXueN8PNkSorIW/U7bWQJEUbffhlUnvpFzpgs
kIKG3eTPYhdFrV+Pqa/2T5qy9JA26ENWmE5nu/eqvhctYgkNBosB+sT2kjWK3k6p
CIi795WHhpBC4GZ+r/74Jc2eEf7NmbNVHrY151IQBemhaZJNu0uGrhpkpE2U1pmd
DYryYFTiGCv4eJBX11auOPH2wJKgm5ba8UghkEJ09N18vISFaRGicRYVN5m8taNc
zGDyQMYdsNynXiyx7rq6U+E+/rO9HEAeE9+lHTZr06edjN2eqyaOTA8CjMLQTJ0P
TR78dNcAEMkvke3Es9aIF72alzcC6ccj8J/IKughrjXM9dGtWHMiGumBpnuV9Ka0
CGP/m6H2wMhD6gCzj+Ji7JmE6YBDE8rqFnU/ibKYHYHq0D0hYlPchgK2XUF8b07O
ATaKlG1epftLw8+GopsFwuCzFG/nKHar/8kwPlqs00dpF6DrMk3Ca8Hcsm6qYbdi
7xEo2Fe6naJmMig0aLEvaOFEIN2fTG/wqhaKUIMFd9zsLJ9bFQilAlpW0w5fapE/
jgu4SpPrEA9K8z8/SxqsJEDHhy7O7KWjpP8H46g8miw/dDH6KW6qdjL6KjZUbCpW
sH8+KOZE+GB3XW1AuftAtKcZqmW14gZ/w4X7KEPszrkRUwmse2/+HxOMj3SDGIwq
pO7/NG0gZy0VQIqlXkDjBQD/TQInIKBcx/11OssptJCavGrQ7nKNU1cJwcU8Ik0i
RxBLEG1u94R6FLsopp7DplNvUL7NLcTHnUFHGbHoZwsJgJ4PmGx6EXP1URHChicz
mDV3Qvvfx3hFl2ODOM8AlQtNTFcGnS0q51asiO/IAkhFY+rSsTE/7YKlMkRLMHnT
AzXlosWXUY8WaCbC0jj0SNAJQk7cGzERQsWJMFba2DojiQCG2oH47N0US16DDaxw
cn03h5s4HZEpCBxeNl0om1fsBciwvepHL4kStaCyU2mAFjsAa1jnIaifpcpSSGGq
Yqnv8izboPbRUKnG1OVoftJZNH08c8bgBWoeN7wR3n+NjxZpWjDqEpcXOsq5x9bg
uv970vux+zYbvom45BsqlV1TLXlGoLn5dMcYGt1ZqChLivhe498ev9g8kVVEkBDq
g+8T9t94HppiFsmqU33LOYWH8oJC3YXiq20ycJ1Q9jKgiJETZ1r3n4/dSXcxceGJ
o0n6DMe/m6+MYvnWajHMWDYuhoJcz3M2IefvU0CyPmQ9DMyWDtcRON35rapusuLf
Ae0uEmP5i0PSpKTiAE28quoz56pF8dDKWfYzznNgWUnjb9IL6tWIe7pFu84BlPpJ
MvqAbW+mm1H8CGzbzbTeaUtySViSL4snaWlRSQf4up89daoZE1IjnQHh/ASXHrvP
Sv4IYbktAKodXV6NfKET50xoyUhLYHwOr5bFsAZ1anfudAuxJBu6h62C9agW0JRr
oqX/yxG0UgkRfqQrecwYT43dQgFV5EwNumYy8oA0HatesIkxXBmo6vFeH5q7vdLj
5rVEzjmg5SBtG9OsvXDIToEo1R8Uxdus9ZoZw9ip8GsescIacL8FFEisexlKN9gg
8QGEHuJu4AF7t8uZ2yugd/uwWcxidHU3qXngqTg3yE3hJrDGRg1c6CN9wJ+1uh6h
GYjb7fPe9gKSFCiAbjDec1uA294asN4Nw8gVaE24hHQpArzZcrFRGu+L6oTYyZPE
pzWesypvdH1WIqoXOw/ejQKJAvzJxvR3y8J47GMbDp17rWqF9XBKPwt+Pws+dS0o
1SDaXMBS0wwzJhCnKjMI8JK+6iKE/KDBc2Y7GiCo0P3D1e3ZQkMjevcz0HxdvOnE
wSWoCyEwNes0vV1I4FXLyGJeBeTaueCDXo0whKZWv9Q3yRwqivcoGr7IwstBbkPl
LiI47A6liZILB7S+weyZvyzU34jycABBFiHMrw4NOfjILUYiBGB7P0ZyGXzESVw0
XyEoNasldDlkzD1Neo0rHqOAmccqhSeoknvDNcGx8jCvBG6tYbZ0jrwwqD5x9Fxf
7rvYdLrRAkUE4v9eRFSlE2p/OkBQHIo44IdUJHHM14cu3F7x29kyg9pE0gr8tQkB
pDwoVF8FJm3yUpf/yJDSqrTKqi9kuHAVr5Sck67Mfu0vsrXRR3+dPctfqiUlUIoy
FjkORl717nwzdLqTQqe2eDPDfvG6CxGu/n13MyZmPFv7bCrrT1S9GVhLlszT7XWq
M5OJcQVVEJoFy6I9P8o5U6rRh7o2eu2OTZyW4CGjpMRYLVWNdZLfO4GCL5eg1wBK
uY4yS118fcEH2dUP3Qz6fE0kLxqIV4dik6/p1JETZh2NXaxDI9jbk3xNn/C3MP8S
mxCzMBD9RjJybQs5svF7S7CIjbLWyd8BOY4l2PAWWH+MUsX+iawJylK7He4sT78L
+jFEvfmu0OdRqrvAK7FjUfIEPlsCRyagedWqbwxivDGxT/ll6m3LZ1c32RIdC+H0
qC3J1htm8uR4Nt1gqPpQuMx4A70NeR+zd1OepfT7o5gmXQRD1iOJAzu+xK0oiYRg
`protect END_PROTECTED
