`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
g5Z3hzKPdJzgDB8tmeQnM1YUy2NwVNK6MWYu1jv5gc8HFBvuA2I2hjLnyJx80zCj
oYti2HYZNj+xBTqNPuErYUpuWWrQo9yzpUKNdBPBgmuoJlnUeGA/2TBWvAU1yKIT
jwKyw8VsJzcmfMRkkxS8+jPoWziLVHGcZaQpJil7Y4TaCMKVxF2ilLexMh9XKP8g
fyjcP5sDmLItW2Hxv3Ih+XE1RtEt9CKDV96axCnHHZokow+Fd/E/s20BFQsLdJRc
87ek01IvaR6x/TmNyfXoUBpgpcSWsumLfjHwKudizMzvB7ZEXoNVVSPRi2ZT4pBB
ajafVu3PdZFsipSr2nZTVJgS9DKoLOdEm7nbwWvpFvETTN6bMrXuWzDYRw6vLNpX
oVoQB4hWs9KqNdNbJaaBVXXOx6c6m5Pvr3Pv5sFuTNn4OVQ1WHtzyUMQJKJN3V6Z
8wEwhSdU4CrgxEW1ykB4HpXswRJzwvcERzMjTvwZuYmiUrXs8A7CPEXt2fgttlw2
ND7vWosr4ScpIkM/8rUe7JWNOou1mitEjM6DL2RtfxRJCDQsbJLr9DQpyWWedcxy
xK5m6Ny/HYEpcp7ShicTMPqdr4LTis8Q290WrrK2EgD92b4RyTwgdxE0/J5P0ZPh
u9869mOmdkbtQbqO52eX73p6xDjSGTEB1i4ZtQPFa3M/+h7Q0yNh7NrEr/s1jT5i
99D/IwaO9iU7s2+F4VjfIKyTWvRokWUrE0umlF99FSDKTV5n3XG8mYSKpil8Fd3y
Fnx4oDz0FCTYno7cnBUqJOWc2n9yu8Z7LocLkVJcverkLCdkLILZpUYIdGVxlTiS
4z7ymkdTse1GUDZSXeGX+ln5nqSwW1On2Gr0hNcYDTTvCC0p9TU9XCxlfJ9lVeez
jit6SNQBY0oVVKSDnv6q9CYnBLxgbS8UAlunaGxhzEicqkR3f4//C5P3eGajjsRw
NCuvm2vkVws6V9BPEJz/lgr+0K4of0AECNVfj2/r1aJZQGiPWme+TjfWM+OYl/MZ
REJBeXJnNMjZkqcpCxwuTEeInHIQKWoX5SN0/rdkaegKVDGUyyo8ve64TjJdZW4d
CcxGwsXGXL1GjKf5Ep4SqrYaIKvU82CmEJTwcXcwKir8fC9iCnFWwxLNRTbx0ctP
A36gYDfUdxeRkCGeaSp3p8l8QLb5Oi9k5Cy6Hv4jHUr2V0N+0klHOwslNYybTb79
/HtpAChi3LPRjGFM/jCBeBY5JXcklNlVa8EfLpCuXFPyQrhua+N12SJh4yZUT/FQ
wwb2D7gWewKNbLIH+4jscVPUNSAbsnmsJNCj3syFkbJ8FWjt37/e6o+y4hj2ViKP
lqWl1N2DQ7UY9dhTvF8XB7m13AL+t9ZJD/YLuBwB6TACKJ3ELGlFIBw+3noDEN2u
iQCBAeSlB+ZgjrjyjqZfK4NLGpKY6JGa7m90VSTDc+r6XST74Rlsr0rtrt/Bt5g6
vy1yCQOrsFtxBPKHt1R4w+WEljRdPlLop7YLND3tpVv3oxaGc3Vf3SFnsUtUQHO2
sIGwvNYiPqeM+sxPBGOWURv7qukf9kgSq4bEt7qMsVJbhJA5CjRMAtDJVrV8F+yK
N4HFWigD36fIxMfLvUxgqkcBmH+1cW+DaXdwLiCUdoXGY7z6YiXmdeSgs6so+bkG
kunnYBsczGq6KOu9XKdaH6vaSPByM3kD3z8ajc4V2qo+Zrk5pi24rmcoyyUArlQ5
lwzwJBbaU9tCeW6Xul1o83oCygIjcOwKkCFEakvkjalVbyBZn+KlAuo/REIX1KOJ
Cp0gGm9AshmqCELhpkT+nWlSO9UvqWh4oWhgKDQyebsrGuUI7I4y1YW1SLlh843B
zuXOc7SSsOhcwhBVO75uAEA9N54uelh9YhsUw7h749laPz1hAN8GyUKFIDfIOp4k
pN6p1fn9uR6tbB1IR0ox2FWb1+h5/UNOq/qY5iFLDi4kdd/MUKnWbB+9LBcdS7MQ
e7DFD0ayuCBjayWPF1OQoLikgGHPDTUp+2PhId3aQ9UsAKmniQ4ZvpRwHUm4Fndw
hJ3sM4lSUFXF6Wm7Lj+lPoE3+jL7HmAKQ5g5WlsWECnWhTUu0W9qd/vk3su3yyjB
VpIZ5anrARMH9mMB2FFNTT5uGrdiMtk+mK3ePuFRHaixOcf7n0TaGG5CPypy9z6E
lGKl0aA6jdxLBf+CeoeRJ27FBU1arwFY5OYhhYcN5CY/WA6y4WtHCt+HjJpL0LW/
hU7+meCR/jdJHfVZCMm6nJSYIuj24aNkE19hjoKhYwxepQWyFe8iNPVs/MJJUTyh
+ZGF/UNXr/5RLINpxXq/+hx4hHdiNmY2szlGTQnSC+ASPUzwYF643atjcV7rdeu2
7hjGQCgJ9Fm/zOt6s6bYq3IX2BRgDYCQkEPjAeVMYRxL0l+5QHqLdTWAg5yh5fFZ
hDyZSbXEhYuQsKAzHOQAg3uOk+WKJWX8hw6wTBq53pJr7cp704UwT6rdT7J23tqV
OJ3SFqwLjLdRj4uciz8W9P95JUoq3NVVWMTrBw1KIJXr2oIRYJie0qRX84hTVSs3
CgFzmH+IdRG3dMGYAicSZhENfiGyVUF23BC3PrQ5yXFpspWKDgcCGBlKEMMWDchz
qPz1nzwCN+z585yaU1P0wVW+D/4y4R0SF1tOaXCzX0QFQYzUrwcPdGxi+UEn5ETg
fQwyc9moFwqXPWMGUDqGKquogIvrzOF3p8BszoqNLWngx3kqSGUxqhfJ3JpCptUc
bGC9fnZCuqoteMP6k99rD1Kzcz60/hDncywNkwkjNYw3A/YH53otPTfbtaCFCGjC
R8P6FoZlokOZhVeK0F0PTGyCClMX4Rn6kb5QxzpAt8aBRj50BSeN5FaZMl7tKABZ
xaVbk0/nWlPzyGCnVFddI6VFLKOdlzGElWwc9sK9ZPCuMj3WC1k4uHEgc1KBHPQn
jHEBTvVRgtKTFCXTVymooGk4oPTwNRYoaAqUvK9Ezom/YXH74s+jDvO8HPFR321C
0e+qgqeBRIqfws+MWhFdN9V/DGj838O9mHMm5qzwynEvZVBao546waWl//d59lwY
ZAClqmmgDDMzXLMMmS57Cr7zt/MjaDf41+xuK6T82UpXKKA///L1hYpmIKCwdY5K
3Cklg1cGx63jv2HKkcvkLWwP+Qm1MekbI0DkFPa+TBorYXLu/8nFoZU4vUuvx8so
RZ3oBXlErvBE9XU8RQ8f24qI5ALOplLhQfKZURwlxhWC/lIDel8KHGAPYbm+3m+L
eQNAkut6BJzjqqoJZNAsos1EqjIXZGkt620vQusg1WPpOKpyod+C7dBCydNKb0Xr
P0ad8SUE1GpjctdZEGpimTZ5Z03ebhh5QS7OnKvIR3tFTIbrpyBLVATNBSo1S8/e
fLB7fAwvAVrjWlPNf/mlGgXYZt/T5VaSjQeLqIWQjKPpR8Bf512b/RH7NREDMxXZ
uadkduVzVOlZ/hpVp0QGKcX47lAWJZ0xjRSDepRipCkpT1/Cfx5Oo0QbAPXaC1nK
Mjq/CoZ1TQZGT7kTTziVLgsXGPOcLJW+NjKFvgMMsKIuQC/Om0Aq8bFvPNGl1+F7
FhM68w2AVw1hZjcjn0Tdd+EshHX3SLqJ+v9l0Qi3Yg8byZfZhBFUfaI/pGIjC0dS
0cKqibK+NwM1ZXresfFhRYTDsidec6DLQdScmufFAR46zyeEbLzskV+3e7yyIlDH
2+2i6Jf4DZYgBmN0mHaQiS42jVoz3pqcddx4mAP0/RzTMNaOZiN8z5vH/2ELGqzf
9YlNxj+NJcZFdl6pGpfqsB5ye/nMAEbLWDiIcxOPGTtPSVSwMNIrTnOsrKtSk4F3
YTJgVtFMfPjh9wLt7lPIjgs9Ee6h6akegUt8uEF3NRGe8bS14pLdhsg6P8uHwjI1
brYB6EC2mdd8l47dpPvn4E0ExfnlJrCTPC8dIUgBxvlfPBfoQ1tM+hEBhdAa6Zzf
rUMtkgLXH5A6MSN0AWG2rWLWgVZ9bQKNmCRIQHLR3dKSeXyvm/+rlqM4iBr5LVZ4
QJoGn6AyrmwYzGBl2MjJ6iDm56lG6er4BSYVdVrvIq/dV+pKcD7YlVkBgPBuZy6r
3U/IVR2lfpCnEtoLt/ze5cbEC3lZgPl09lB9ghRPf4wHHWAqQf0xuLcCSwokXPf3
uEJoCVYyNgFj7ZNL1Wu2r+kqx50UZvNWNalczJ6CH2vLXhU+J09Ckv6U0Jp2RZki
BoqYhbJmrYwlqIquDNNhxVQAZsCcSFzIBHF9TMGxTzYEaEPLLPwoC11YFY1uhAB/
GGHAkVTGlkrrwR9OnJrv1tDH8uXUSkl5gQtJM5Wo37uJ6/xKmO5RlJ+tzSWPMP5l
W6xks7CvlZxKkn2fhzn4a7tp0SpLDlFvvKYcDw4qHjg=
`protect END_PROTECTED
