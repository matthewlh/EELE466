`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
ulDVi4gYizh4NiMJ2jI3xjK+Y2cpZSJh/Yk0eIvWrW+P5u4/GIDAYEeNtuM+tzM1
ACMSV59tTN5q41ehsMzF4Fs3CgaQ0fbaPOcG+lZRGtMSSWe9KJhRe/SoqzVIK1ez
g9JSSiazMz8eJmrvuqNyFORk2qq6r3GfLySOZ1LZ3DbeaFOLFdr+sPl4rCcH881P
MnTllnlcVrbP4gJZJpNmCfYcQE/WcxFbt3FgFV6e/hjq2xbdO1fdZR/c02Tfwj7/
RZ4igYiU38R3/QCE+I0GJTxc9apU/VpeahZ+CBKgiq3FHEpqOOiS3Hkox4TH4G0o
hqSCaYvsSAXkxtgPUMDiCX6r0Gv27h8IyeHRsVWUcz7Q9aWX3Lxvi0woWA94g/Km
ztLQas163qIIu713vIm84BianSzfiYhiT3mfj4CPc1LP+3TIQoiHYcSmmP7IYt9b
Yqa97SwuAGTrZ0pTl/aBydNj/04RfCUSik8ohhOIs/IL5rWI4p4ael7c5rnXHFGt
IoDDq2iMcz1NtH4UsC+ux30KGqqCuYQOsgUm7Kk/7qVsT0V2qgVKoDJREXPmFBS9
77Qtw3iNiDxa/fBuV3BL0iOXv2xR+NqaaD3vxCtDiBK5fTOCAH2QZrDYwD0fkdEv
9rAlVEh1xx36NruR9ghal1OdWDnc1KeBryY5cjmSyDNCShCNr+s1DTHPL8vs3Lje
l/QtfUppHOAKCxLYQ761iSP5jQwJiTXB4hMcUJtjiNM2DFUlg81kua9w4hNvu3EC
n6lJGjybpXhW/MDURqI6+Zr/PYeckYuMAfa/1MQq49eQi4roaPfH786Mt4kBmDba
8tp+DSwSMhmKG+nNCMzEVkAuB3+mXisxLfUXJfINzKHlhswPd970/3UV0j1zz02G
BR2NCvLbR8tWJpV/TH97t19Xozozc/eH4kcTXcqtqA8FSAPXo3iEMQi2Hvs+KUdk
xeykOBdkKkRk9sIIGlk/M9H/mx/zgUlQXVi3bywI72dNGXI2WepMYTHxVf26KVhC
Exq/qr9dIR8Tjzg7LsOmdpPhAd5mnWTJYgcpa1qAVX+1CeE9I4yrO+ophmnaJGc9
AtZk+RNC+tSVgWuCb8Ab7PSP9LgGyl0xKWQIYHLtT35bb/kAhRqn0hrAiHwwki9W
v4o/Y2mj0andrF6J2q/sQBhRTqtXvUc1uEGwkX5QsoGjRuPnzJ3lybkGq82GtdEy
AvYmhvidCsLW/gVNCkU0hWkKH7ja7fNG7l45a8147OC8Kk48O4P+ydr8s4hBgitk
n5ZTSz9nXLOthZGfwMWVIxd+A84HBq6iDkR1BzLWlxqvVbIaKjcPEdBjQ41q/zVR
bkvAdHh/TJXNT/vKtaMXireQqWJ9KgniOADv3nlytgqzKEJWTUjGwdkbPZcVneke
HjWQTVrXS5C7/Kbc4dWjQOel7RClo22FzMjmy7ym0DikLjOUn2rDdXCvGYU3F+AG
M9duH/kPNZOjqZVM0UuGpp6NwkzDGHXiAW++KEPpW/2SrbQEgnkLmm/mH6zoU0Eh
ye2X1m6r5ED/fwkwTX5alK8o1sEvNWxmhXwY8ge2VJiURaa5OPxVup14Hn5wUAOR
vYiC1/Wzgj9KbiwNagWbxEK0bD3jtvalsH/p9XM46dI/EOopy7ZTmY/xVHikCKU1
KvHuD8RVbGrUcVcAEOXDeMF1Attas3mT3QyUEAjsz0K8mWeN++rsK4Te3lclge4T
EU9ebGT/OBqz4GEDVLP7FwRzpJG/JuVs/LTudA7HR2FJscDdEmmKJDoOtA17Xhg8
Pf8+aQY5uEoJOM402rzR5tsEmBSmJKXc17xY6mth1RV5sCosACGXuVuMJ6HSZOBc
r7tBlXmdJvFRDU8YEdQsTNJKTkoK+/kZe4M4vQojyXmZCOkPth65bfLmXAzu01rd
FQ+5zcPzJU8en4scvbQ0TV9BdSY/nMKhK0mrTKM5S5ZQ5Mhp9Hf1pajshlHaxDKm
1EUX/rDaRXPFeM8i+Hg209cM+woBh1L21BxItErlK3y8/J0iF0bR0PmcuK6FXVvL
c+9OjHuuXTJOwYwhNj+KpHOIb0+w0HPjpfHmKKsbi84G+m3y2dxyGyZ2EGASxJxn
5nSqfvvP7O/m1GeJYrrCdvj4SGY/w7/L/I/TKe0elc8oHLTKqLAmFdqSG+/FLTtX
3ZC7TmV9NWVP1WUNi9vIkZz9MZ+qD6z4wPecDkDfXSMtrXi3h4qlv3+cigMdGrY9
p4Nq6nmh15nGzc6XVZG9OWYsnd6CyK8Le4VuZ1JFf0y3H5BMiF5yoO5JGbdTuJMK
h+89ZvItOlezA2zjS1OzjQ+hkib4DaqRMDoU9PYoOxv0lNEO9yHT3Z4NyUuJkjBk
IhwsCuMT80NcOxuk/y2nHXByKzS0p7ybVwpDSQ9MHvAJOKA8bEx/IAHkaxi2Zcd0
eORRz2+xc77esfHkUVouSeE8n4mTc2aFKsvlFLEB6MSr7rd97TebPatGSGWjuaKn
M9/cTVWQ8vCYKR3SZHFRGNVOe6n4xUVEDjJFmoOJ3j0QyvyjpG9zCjxPCH9lrh/l
zzlGlyThqi6uTjZIct37hfEDg4bCKfUwGYPKH9a1qs5ntbUPu5RNPfz+rAevRqJe
nicTiFX5SkxOqdXSnL4tPiyQ6g3j45xgGVJl+hciWvulx2gd1pjk6SWhNAb19Voy
K7n0+RgXM2dzA32g1AuWDpG7q5hEWPbP5i4GH/A+KbGwgd3LCcvkjLshS0/KlzAz
NLHGIk8qigNl/3aurZJULOsy/g+VoJ8bQQEzT587diM9KbqVyYwUA7C6eMFfYqi2
g5T/8/v5Uo74Pslv1lHbhUnyZHbOF5SmqGONX1MGRwF9vszgoJsKzrEl3lTKlRVh
t1Zoho7Jdg7eP/FzT7A0/X1+wRrIQfGSxVinG5DixvlfrR/eWFN3o9C1gbd+HVk+
af4po2Eb5kyMFQusyv+TaR3bF7aqmStvsJvKCZaqUxvQUI8FtHntrpA4RGda4TzG
n0DwQTFpeZ6bDZogvbYJBPlIcJg/ZX006r1tnJjxK7fKisp20dVZJsXaz7UrA5fF
nZFyLBsK9vZ0paFkZh5T4CKWcQ7iZG6PB3pU9otaC7osN3mCACwXADzDVm2Ifq+V
TVDkhaArSxKkh5kUGh4qENWanz5f0U1Y24hRaT4YCElE36/atmu9snDZazaAQxIi
fuphxukg8alfG+LuuuBZUSpKKxm1IvgijAcBGcSBL7ahEbxUm9VROIOn8BJ6TMvm
qKiCBqc6YKxh5peTWE8UfcDT/mJ50GH9LsAe0DtzPMF3WSgS/dbrZP0SU/5KapkT
4Uk/qp9oRrUg0cPjjeR8Hs+DDUuDHFQu2EpF8jD4TcQKcRzbsN2nqueyecusRZ3c
PuS/v60/krgPN1oJuiPDKjibczOVoejVjLs836uqKyc06hoZ8mmQYxeWgSrQPWHM
yvBEPIx51MXemKnaXEzidUvvWVegvEJpeSAewR2ITd7pFHtVyJryoCy+vqAi6VfA
BNZ/5PUIU5X3k1e+NGvTDEBtkyARFshTesnM6Rx+KgKqYSH/AWU7CUz/Ln7DGs0k
xMDvrz6RpoNw/V3YD9g2Qm2EqODAT7DyvfPGBwvXiIRHGS1I5mNWCyBlObjgApsL
4l/B/h9Uo/eIl0wQHnzepLrpTh3iKM7/6lWgpReKO60w7ZqDqVuOqQyVSA03xzKx
oewvkQnZfM/+o0GF+FV+fA==
`protect END_PROTECTED
