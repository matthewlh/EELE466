`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
+fkGItdn8Wx7ZLltbjdLfAW4baoQr4RsSZG20rWwRVMMZ0nmHK1tNDBEcqBUVvIJ
VYecGK6Mfsz3rCXr+fz5kP1V1CpKgEJ/SbYsCBwqJ8Am73q4OXbFZXD76M9M9R55
onJd8+eouEpxo0vtz8b7/b/qtp+iaUjLa3mqkn28nkVg78Nbc6dpNPwbuJKMgjGX
X7J90KqO1Idmx4vs0S//Z8p0ynlaempk1q5jPff+NEndVwU4WXpwayxmVmX+KF9B
83xEdhqyO34E/6KJamorbkxOD6dCL9fPMnEpaBs86OXUhix+Bcy8mRtI7cbhwOrc
/sQRFM/4cPNnFl27Ym5fta8Mydp514mhuOLtNFyjZNeAyLAqJ56A+uSeWeoMH/QO
p5e3ysyRaSTNQOPZnVULYOG/PoLeSqPkmYELadduPq40yb1LDZ/iHj9iQq73/5KZ
kH5jJCK60jt9+6WpmwjlLn06FCqXPfoAN0Qk++TwSvL/K7zbduCkE6nkD4wvCQFP
59iqz1RyMVDBO74XkX4kzJUDoa4CoVmGMli68iGXIPdS8avas6jQqCUBQqBOhZ61
s5718eZCouLn+SkUUBzsIN1p3fstkKlXUeibqWXZBgFru9aloHFBMSKY+VRG4GL9
88mzrgcSunboMZJq3NFbB+S+JdFCr0rcFGcNvCzMhXCDhF4YEjHP9NpSWugRGQsg
LiJgcz/Y55KY0WHIAColHmiAZXCVKKuEuS0jRSnF5lrk0RpthRKQ4rhFrfz+p/Su
1JhhZF6/YmgazZ5aS1oHsAFguDDZdf8rZLoi0qud28w1o3uyXih+Mx6cXs2mYSV+
AFiDGwS8llvGYVaZAY4qC0GXMmj/puNwrGdccV+8sxj8Kpl/HtRDd5EOTPEkGpr5
8PbL15gjjkk8Cnkqfa0piL91yA1YmHzxQ1ZaoNhfu7hNiVo0GfCVSCps8HLIBsxg
fcAIQrOYpOZjuyKpn4tV1UqmGLUEYQvKNx8RNA/V8neLzX9gxqGWPp06waZzhf4v
fu2/hHChOWxODZANYSpiFxZkocE8KUH3CqZGWiq6uW6cLaeRQBAgfxDi0RjkDFB/
U62W6FAH3On5G4ZBvW/GCl85TrkvnCf+mG1VU7hyPKhNtp+ZifxR979p03bcvZTk
vGHbXDyKn9LIT8hDHeqTif/Pyq+HFC6xrRk5X77P2+i3f2ssl4unljfj5Ral9+wH
DekW8ZFOGCeOlK2rN611iSvvMGW7QqgEN4LyvITNKGBcqRAZHkc7ZW/93L8csY7g
dWmgloI1PslWLifDV6vdsL5I+afh7xvQFQhT0FvIGDHmbTctNhyRHjR7hh6n31eY
dIevHkk1sQkE6SLWDaHtYL0BjxPb0wsgbeYEHqXAizSrmCcA3r0YjicFGhcqybE/
0cAiA1iHgK6MfEiS5QMR5IiOU2BrnwzPwzEwySfyAehEDFfqoeeep88d1x3KxnVp
Hdot9uVjZRD9xJTecEGit6y3w7nHKGNdR5t01D9ZpYhKJvIODWSxCY1DA2EoE3gP
ZP2TjM8qOsaFDR3ZwoZ+aSjqottbhBY8FG5cD4cNk0LEX/l2vnIes/+eLcbjyZHH
pdhBCIIqQsELGFPUqiG4I4GzjMWfrqBM9Oy4F//yzXxxVY/dDbncgMhbp7S584KE
oQbcQaTrPGpFfqTnH8aU/W7NgupNUE55FSFaeDqdQfWzV10i6rw8XNutGNDNYNGm
r+BdVEAOjGFadsmd+Z1imiVU1z8R+Qcru+xti0k0frvV5JEZAxypo0wq7gNP0j82
fACArnhak7lvtqoivGk/BLYceHUjxIOd1lSEtewy3g2TmnSnfctnnLaE2FOyp+rf
rF1QmLYO0XPL3GfgXlwPAi8S7PR5yoKuMse9A6FH+07vUAF8OicczXS4I8MCSQV6
x8CU4KIdTv2p7aK6giNXH15Fwdt4E+iA18DwnyemZoA4QpG2xqh9YH4qffzqFmbl
170ff2Jg0LK77zBB5Bv5sA3K7/c/1kwyEH9EwGmNeVv2LAmFTjlJhTZX8iLCVE8R
JMLfwZ6wIziaEP8KRWmLN/MZOWM8KIL/XTysaJkOBTdhpqj4ilMx8yZwRMXTGM8M
BZxODeKfW1JYWhhnWjA8kiXcOsdGk/Y/Pd6q0SqPLKUT8UDMuTLue9fproNuRkAS
z2K9Ib0+6YfD6AbQhO8jwGtDJLHIbD5sK3E7BS8YM7X0S+cv0RF4mh46iNVkrGGl
HTZ/BMj4g8br0bVZvlMKHSIsIZyoD/7+P7SvhLLiGCCfdEGxKTC2vslKkvFz36qo
3rw4qUWCaDY/nmoVogY86bqzokP3MEfnzrIkNRflSXg5Gqz0LuqLSj8FThKkA5Dz
CrMiPfuumm83SC9Lrg1o5IY9erhOY5xxi25rnq4/cS+WZzKFiWWA+78dAyZQvNjL
/A/1EV7BaohZVF1lm/0PouGJxZpUOfmqArz5/G4vc9Hv/Lgp1zlKMK9cgnhJkD7R
LP0CgimMclnNIdx7VqNTTF6TCl9YGfKt1Cn4b/bG5nEjAgIjrxfPkaP0xKVC44dL
qIeVYdSHBnniCdpXcrZBlz7El1TvIZMdpdir0weHTnL6xWFX8mSVS2Rmtee/NCyN
qOQf5+YbaXBWDVxMfRfnjEKClc/eZskBYeajmXbDHIzmjUF6kdINZZUaLAllHFUI
t/RrjYSskgqKAgjVe4YsbPaPkO5nPbsJN2IMMOnzRR1QiG2optmUcEuUPe0IHxQ9
R5XQs3IYqShjUbYp5quhQbuWQ5YCBeDr7xnoVJy3N/CD+N1BEXZT6ePmLoOk3GQR
8U6ZblkBvi7E5X7Anh3mRr6ddS4jGYdcJPS1AmP4HACIjpJ8oyPUPE6bpgszrQWv
ctztgLy/vOB39qF63TSLucpfx6l3hry5i3ijEowgWXvXeH5ZBqXSpYIuzdjhntDL
bDztWoIMXOPUIp8RBKN3j6jkk71bAPhRewRSoTJl/wSgeaKTyph2UaZJUWkSYtlC
RoVJi/LXNH1IeYCKP1az8ACi8uOCNiHf2LiOXo/+jir0zmeqMI3W67/H1GCObvZ2
ppWN1LuBq7c9x3lBVnzA1CQx6MB3yCVGBz8QvU19ar02AH0k9+5xl6/BywhgwEN8
eiGgxx4RSA1Jd9vyssACoh6cB92E3IJENof2sPIDknYcjTHMmOwxCBGRhjqdKavb
ODDnHEnpGC5PogLh8idbmdt71usPRVV5tOUj2Y9Gb4THqevqtIEWXk3VHezhXY+h
ZgX6uVBalHF+81VXte+Er1qqea91xSBMtTI2vg/XxduDWVk7kSeJZ+K4YgG8e/VC
qzox7J0V6hsYpCwcsb2lrKoTp/9Chkfn+dEGidOR5ZaQEBcdhfEuWp+Lez7cObQ7
teSm9LQF+cZHgBhPiXlRBTwwuVZB52SdHQRQpR9FXrE9y3KjpXy9P1RdWAXmNZWO
TD7VKx01m7H3VzDg9xcL2DplG7bnwGx4yHRXspfy5rrwWeqwZy1flhWzSu/DFfPg
tLKD+DD7YGqEKkudW38dA+og2qUhYkngTRFzwvUQqHXiotXTbx0AcdxCUblyBBJK
2+rf4F0p2qNVB3yoSCk+cK1/QBm9bdoeuji24SkW5cDTenJpBvUIZDTWTmWoU+E/
PTuTOi65Upm1n1wfTTlx1KW809GwaRz0wIVpcM58ott0ePh9XQZ0ia7h3VaeGPRt
1hkOJnmz9MBvFjKEIMxGya1BW3WbMV7oYufPzM9R5N25M+GiKRRlFH/jRXh+Gyo5
2GZd5Cs4NbLWkvTJhEfOdjGLT+L/rzzGgwknXSO60hFZhv7QwsflqPWhQbcCwBGw
auIHu2CYGrDA+PnjaDAnueffOJIWouGrK96x0v7El6wbXiTZbB6GFYvGe5WqRO1G
Sps8NDaDHHKfE6dddVInWf5m/bTItwyaOFjKBGNy7KQwIbTTHwsWp+I4sINra5Um
ss+zK2At+FdsgPhiXEihMWhbo0eJ1j9eHI4FE0meJVS7IwRnJHxah9sodYDoLqvW
lyJp1CQE9oS0+CgNicotxgheSeZyhn5kdgE9g+ajq6TAg6umSo5IKv1fvc5PYJql
BRV5ppyhQ4VUkiMt6iSqd2NyFL1vUzGc+6aA23T1Dfk0E/M/ZLPK5To3lyAQokKt
UQ0Qq9IqxyCz6Xu5LeOETrjDPhUtg5RIRA14AyvCxgp9i1hlT9X6E1HEw0aS5Crv
TZlCtztp2c9o++LqIrPco6z+Qz2sPtqu9mynkTRRJawxV0DzaRnh3DYVrxUO8qX2
9v0D0BzTWpDsK0S2kZN1yxFbTjZ/abo5qX4+6vmx76f8P93msSnXsKJo7XUwcTR8
TNyrkvJtc+Vk2nsG+nDzN8R5ea2AdigRHSuOQajL8M+8Bq7JkKu3GhompHkXSF3v
1wUvlC32PxQRkQXK/TgN12+RpkttrJOyUaU1hw6Kgz42bb3tvy3AICxvUghIvIs5
aAtR+6TMgKvufBZXxuZNPzYlsuV3g48mCrEjW1gx+piFlAJFjO1+Ybg4Z8ZH5MW9
keeQEJ+XDcg1J54hJHU7LwS8rS9zSZ8tV2+duNtgHdej6cZspleEtxkQ/rNBa8nW
tGAqxLrXZne1byl1ytwZ7FhSFd82ZWkU0vQRdoM7VzW3UMKslLD5MJrysc2v46Ai
3ieJxQibP62NvKKoTl+oZOAeekhAQuV1cRMkuHKw3zdx42mSwu247scDNi3XjZdZ
4LXQ99D252102I5n+lIUl+vByqUg9QDM+DHHTTquXg/ulc5Y0yiyrjMOmfGZZZ+x
a/6BDilOivzUMbY2obwK2Rkn4W9BQuC0aPtZkSiiNLXa1yzxL7oHTmVlmd78BX5p
2Js1FHI3qIwY91RHvOwS8dLeLVtP6bUkoj2ifB3vl7zerzJ3kAsAJw5kFaVo0zx1
nz9Bwujptv1pUvyfJAd23B3xI/aTLr1xN7+MMkxTtMUUjCRNu1sentg+wbk/AWYz
AeWevhflNSP9mLD7XloL5Mb36Sx0YdfHSNaXV04v6IDPGWXQsj1fa0Hp+x/pyG71
8jtNyCgJvLxb8Od+72PBpLYfIbHSIB0Rr2C/Db1UKOdpPqu8XEDwKvMCuYQQA6aT
3Q2slyFKnwWkSb8N2NJSW4n0+0AzKCo4CNkvmV7H/tVbrkkKJTIEVuKXAhp8fxQV
8OzMbRjIyNq316VBxGhe64FzcE8APTePTcXcKdsD6m1rVIvMX8SELYti9+q0bimC
wIsbSh142i9ncahMFtTlFVatBrbevQgQLXwlvYlB+w2B8mKsA+oz5hyX/IMCwK/n
v1XVX/wT1wdz2vNohtzrCdkCh5ZanpdqHn9Y3ZEsoW3u2WLlLlDmwOyKyB2wnBGF
5E7U7FMR1Lk487tP9pgEXBRQo4aw66r92zh7Dkh/O9wYEitHlinuO5TXElgXFBPk
aFCy/uSrXNBzNqdZNWxAMUtJETQp404MOabqizZVVpE28vAAsyHvjqY11IxpQBE9
marCaFKxhdeZ0BTF5TI/LxzI4JxIAX7hAkx6UfWiEl5uwYFNtorVPMBxAQK8fUiN
d2pqVKXUksRw+O6oHeWeNoZCR+bqh3/OpzAW55v8T8KKA7Qv/wvSHxTtIgdUYlkV
riE0Ag2thIrCGeWW5bEI9CTtFEadf/uEps/2LYM4OoB9DxXj+i2dcE8cVKoSERyt
H/izvVUPRQ1W4tLqwBrlvX876+J2jgFhXT+Mz6KdOhvOZ4ERHytOQSz2sI1bLn1h
yvV6BVIEiIt7lcOAlS0T37Ydp3PXO04g5RRRTXUvSTyTfaWkL0tjHBUkWFa9zMWl
UHd9B+qkDV2KZiH/bUUDmqR2OcaktZuYf9XtJJjIHOWSnk15TosX0XE8ik6n7NSN
SzfZnvKlBWbOgck0iMBVjiSPyVo4zPWNv4GiCbIECpfJOfiUD9WAlYIDK1EFi7hX
rTHo2SaQ6WHb8wZBweUOEte6Aonth5HlhJPE5hKe3a1SxwVKQTPcOfo3puHHgVyU
om++vYvGA8Vlwr06176PVZu5OnozJxU7orFToJ5aie7f/PnjlYLVnhTGElr2a1gb
VmHCOOQLfTQZ3y8kFz+nsU+0DjTqHKhDKvnVPzku1sDwRDhkx9h4gVMHNE8G5gcJ
SjjnhhuQCkt6BZs6FlJ4DUJiJllnWNjP6XYiuD1kTE51gHh9Y4gel9/7/Ldy+gHT
Io+cAjpaIKw6ff/1Gwa2zmKkF3eCyvaW40jSXD8yxEjYJpZtfzvhasD/J20LNLye
nQvK/b7chr1I1mmwPIUYUrZkTlgaNPYR+u8NZS28eeliOUM+zjQayiz5clab1i5o
chJkwlgq9jy2BBCkiQhsxd6o5ntt+aKZQ2tWsAUG4LPEI2NArPAmYBhZFllkuo88
nkiGTwsJ5LSzcpPRTQof4TwgZeJhDgf8dALjhfmuePm1hT/2CfsPtpJy4kQxAHE9
MnoflO86h639xNEfOMXS9QbOTGPvj++/xL4odT7lJOJvc6jXhQ0V9goJKJ4O/0Sx
wF00SAxDAku+j+bg/j5I0cUR9Sq82HXefiz1lV8VbDAfJtg5xbk+RbHX+jcBXtth
QcGnO+cCoNM14XRk+7jMAtCc5bAcG6QRLZs7ce5yhnTMjxVlERdf+DF+SF+RH4wg
ghT9VR2BWxZ5sxbLeyurH0/w/aAxrRl3XB77Sn+UPrlM5FV+Ld245gf2rzuiCI76
JAxHEJtoNl0e5ek7pnobbLs34O8PDaNElpDkbuEKgnePjVAYORnGVMWDw3rzbqhF
UDsG8KYD3eQruLD7OnPDOiu+NUa7CNAKvirKWngS4xIy4Qp5B4jU4qOUQAzjlpO0
s91SsjCNcIDz0JSMRMd5Rsk75JyWbur7vnsrTmTd8jxfbEphJTj5kukKduhFUBmu
OyKNUTFBs0JAn9iKIQS8I0bA9gKMr0U6Uv4ArGtpuJ/P/tKZu4GOUnZx/Ngtw/1T
wTNwjaAxwVnu9gWb/GRXQNVdrMUlUZNwi7N/+btk90Sgu6S/ja9BF4Lqj7Vj2J4J
NUHNnA/+lw1PrJFodeN/NCaD2duDvW0Kc5KyG0OtPBKdnQZImguCBJTRV6zu4Pkt
vbzgxrc0JKG5gCYTYUcz1VMn1et0dgz1VLD+wExfKNyZ12iTZR6TtBrmHvpbkQo6
n9PfvjbDHILskw9dRfcf3KQIyfD4i+UERg4uZ7hBYgOiSR/2IgJQ9CdFFWGDELrj
eWg/6iWEAFIQOPqSt+VOz6sTBQQSbQLRet64dcNSDY3hy4tP1HGHh9uCabmiWfUv
ayQy3wrrgqOXZ+67YiVBDhIkGF1iJl8IiNafF6QIVWWD2gS8Fu+LV6loVKXREnYz
/0BhdnjVOIQx4Fx17rgTd5w+KJ5sOxvKyiSShvUYPta5FVG71BljyMBu5G5AAkdu
8Fi+OggXowAwSJsnpBp4YhzMKWgd+2e8rRHMSw7AcnEAK0Q34NUMmBoznt1JdOjI
unZrTojeSQwA/fbjjG7tIcACm3ACUNEzMXAKziM8RkKGg0SbZ6t80MRVoOxmFCI7
idz1L6PLJSEfpOnl+/g/MZmN9nC2jCMzihrzZNdjVOYarq5ExN+EaMEM2lLMKp7K
tSLvHQvQaoK168u1O5wPwvG/0PMli9+NcGvYQ8iIGFWUOnuFQ9NO5UfIq5KnGCfC
zrLedsvbCVE6DSNOJABgt4iP+egtQ4gGr5Hoi2OuBmKk4qi913jLtajE/M4Ytwe6
zsnK5abWil9aEL3UeY06YJAcp2X9LmFTKjhhE33sUYUhkoGYyNcLcgLOiog5FOzj
HVHoiRs6EGBHoN0C5AvEHB4xEXTs1HkjaAKaPzeKJoREcE6ti15h1R3SXU2JRwCI
nxuLu/JIQrmfgYDJCfoEYkil7rRo6jBtP9ZTw7TlV+8VHpw8oYJSigHXhOlj54fR
IsJ8Nhdu5NmxjS4sdViPm2ZWoAH1wZXJtHjfvGmy8frp75Dghas6UlGUILCQDUhT
UDoDz1DzSIQqDCLOc3uFB9bcxNwhKVCrotZw3HZszpZxHmEIRdLKBUpSRccOERA2
ANCL4hlBqwLSaLfZYn7S5d92NPpzVqZF2N3pIbegZNPXXl/BW3hVehoXT6UKrVEw
o7f4mTD1AyOfH7AEWzy0FnmnND6L3VdOrNgilmnOUM1W4tPJ6FTwX2VAg89RMKeZ
zFrl41PY8CZNJwTIH8ijFTdiSlu0Zk5/ROaMohyWjOotMA236c+CtzkQ7r6J7+sH
uRcYDFiMFI8+jix+QxDe/1eKpBBQw5jXTF8+En9kaE0CF22F/+9jGZp0aRMX+E7S
jHV8ZF+BQa8N6ALJ8bpGAFw18aV0CLThkpb+QdvQ4vieYXlVuKEGKSH1U//Ga1Xs
hya6zjUVgnS8FFw5b6WR1AGsGfmkTG1bxfwr0/vOR2IVHMMlvTzNuf+I80R5Kucu
wHe7j+YkP1GPT5Wc9pG9l84xMnOOnaptjzrTdqN+RTFP5ogFgbo5UVMfI4xFTgWZ
XbJ1KWZN9EqaCo1sNNTfvtXkB1QvVnxsjRRM/VPh+wVpdCsCM7WtFfC9M/CEsloA
M0m+glFJ5Q04MTCtSuUJtyUfP/Q/G2wci3GUHzsjGLWz9GASXOp6SKQz4cYoL226
QgYCInFhxcp5eRQoCyhcnpc/Jahtwg2FUXft894SLndyJBIsTn5Dg8MOYr4dVIK5
8FB6Tf/aIs6vxPJ2fYgfOCqGVsis6PMpywm85kA6obhRI6dCuRAqxQJyPB1CVEVL
+9tKR/ZqensVPl0KDDR5Pzmp1QQ6sv1Iagp33GWmmwDCSHco4QyEjs67yVahmhc0
tQL4T03spsPqr+WQnXt9RT9kpYCRCBq0W4Yr6uwjuefd7s/wPQ7WuvuGJLP7CSE1
yRNHvmkTMzXfH8SkQmITN8bdoKc9nrbNW5V2Vpp5N00MhdxD8mClZbRbxLBhveDJ
8iYyzO5tym8ujBCHyhrhBe8OrZ6OFQoklfAQpf+7GDpZ09CV5QV/N8D9yGJEsTiN
ed5qhQokMZrggTI/vi2oK4/83RwjwKGmbvJFnAUHeXRZOMx8Cxgm3ROjKjGZwWmx
1uUtbIa9IWr4feBNaquHUJM/nBbxmpokeW4py5tb2Xkxjqedgd5GCfG5WUcwIwjY
KGOsDzp+DLUcnN0ofMjBGArzjMuAvDm+9Lg5W1emEC9I42Q4xzI5cQjI5LS+SHd3
e+29/sRkPGtNhosBE3yVI1zZ6QmqiRiK4IOJzSE+1yoRTReG36rvKVd9tDKUd52s
e7LQdLfhqpE0IV5xArEfnzAqjmfHgulY1Hkq9eTBODZEz4AaWcuUVV0aPWPkU8AT
MzIzwHIcQcVfGVZtnaenRJzpADrq9+apZxWhsKQdhV16dhvKFO1bsRHJ4MTvsbEB
aykEFWvGaxAnViOZ6rCJEa5anqALsU7/s+vnEAImijVoPdN2XeSsPUQT4gbeRbVs
O6Z8USR0CJOREUepbYZdUdU0N4PtAlctyKsMoScGUrlBhmdX9kjgR2jqq/yhswcL
y0p6sEIde17BgL9AvumpEQVT78K4B/17pzB0MQpRRBBIxjcyR1q/NrbZXyDK+q6U
/gAREsV6fpf0dS0vqFKULJePbrF0BDZ+wopWhB5mwsnbmiSJhtdY2rJuyjUMigHs
Bia64716Vl3MR1UZgqw1EGn+H6+HJLl/an0YaK7cy938GIqfydK/UIEf/hg6NRPl
aluXv8Ingz6wJ8+ffLmMOv00qWpn5La7aVt9SELndfZ+Ga+pmzH3UQaxEqqeO9hW
YoSGec067cv16e1DDXCE1sDu6/381QKKPgjEfr9P1Hi5IrTf5fABaBaIZS9+ZOpz
iXc7AU7Nv6Y2tQ7KXxMJdySddND1greTnZr3+pAD/Q7LQkwGik+HVO+H1NNLzvOy
ReKTjx9fXaCcnSmss3lACNJFgcvCG4FSNdtsVA/QD3R+C0XkySV6bppd9mEbisg5
KK1WiX9fD6Oa1x2x1O2p2kOEoQFSGg8OgLlXbB2LHOZfZgKXs/s9qs3OQBdgODt9
ycqNtMrU7Qb1q6uWGXnfU7Oadoc17gPoUgr+8lSSUKF2gMFIXesISM/gaKVfo7Oj
iDNFdoXUeZT6zAVPikisj55cVFkNdf9o2MAwrch3GsiRBneMOaX9H9nBbFRwz055
xI+vmBOGjp1HzpGvs+q12g7b3gnAx4sf01dd8OS4Ht/RFxv3uSnu3uP3a2MF0C0H
lLHrur223G0OA4Ek5OK1hYnDdUDYPlGepdrrKd+OBxu9IBJwR0Xg8fwU0CeWu55j
5zKrwduOymXO6Cc4NTrltP2IOHNdLkc1hGCLp5vXYTu+LQKjgrZevIhQhIbDjBSH
K6BxSJ02PxYIiaol5HAWc08T1SnvLlDhaULNJXOhR18xFLirBvqFAtw2FY4D3aEC
EcllX1N/mCLpi6CAHm24XNLMVnSDgp4+lH7a7WfVaXVudROPKuO3j+1DhjmLM+dx
k0cXZRDP93q99muSENIh38XGo5DpSQ6BDekw9kjvJAxrIPCv9zD2qBonKBbpkb1l
KwGcjvAP7SOjtjWHqC3k8FQWaFeRPXKAeEK4tqBdf0vUvMSP98KF0KB0rq6jGa1G
faau2zvT8iMgEEZVoAyeJgGtCThGdLZaEpVxwi9HmeaQw6qXn2H6oxhLV+TcBRWL
StCQ0dlZmvPU7g+fh94K8gzFgSiH9In/rjhfPc7w3Tskrop8zKJ1UCMQ3VGp0wix
CgtkiGxLdPXEYveXLVrrKJqsXCUfrNGxKJGAnS2J4Qb0bKkF5EEQJab1SkZYkyd8
ViWqFMoAjLYBFXrND3eS/ZWsI1UiLHjF+VhBW7OWan0qfnWz2iOr3GfaImdLzuwi
X6uEvwjYMLW5gQgclDDGHhgTzYzu7t5nf+QYLuZ8ha3g9Ge2QdmuMcfXWyaq0FKP
2lr7FPJsR/xhkjQqPTjUFToWr6LZQ0NX/mK/9gGnYWIQojt3k4oO2Rdgr2wl0Oqv
jicm9SCqTHWaspVZxy0h2ZIm/7kSZ97cHVtatzmROT0gyOjSFH9MqbQjy6XtxVS2
3mxS0aS2f2oa1BeYDdNHrFi6yTf8tET65iCTVg8nPsZ7BykL3De5JdSZuTc1FXRH
33rqh0bo6EKjkGsi6RQV/ZfimTncxEJsf1HprIKdbSCE3lkyHTVMiQjSQm0JY5Lm
UcYNK8U1dU0MBWmTAkqmWiu39+49uSO7LA6jDYOuFHAG8M52J4Kne9EH19Y4CWdI
S+Kmcv8tJpXVx1ouG/BO649TEANlRMz2C/94TwlxzG5DN++gnB9ITT6cF94YgYUF
7iQkZMnRxv5mQ+6/BZiiq+npD6EMkspzA80Ahs2NMwXg2SjO7j56ijxh52yYoplh
WUsSRBeI6DYOAhuGYXOsTPn0pm6t6J9vO1RUx+tW+l2kA4JaqVwWB/OkfPHEb6JM
qwnmE9wXQ7exjSnI+tL7cvUDEvOrMjBRCOXjPI3rSKj5aSNtGAywifu8HV+S80am
UYCvbfI0toVPz5IQuNyKH+MKoN3aWTCPj4sbiE6xFP/N23x8Gag+rAUL1ZWv6+gp
3aYMltC8nc6sRzXzHnC+Ix2y/5JWYJKAsjkZt46QF5O5drpdYGZfO98rCw2ayqyS
AYGTptuonpuBle7yG5Jbh1d+aDHpwaePf5xnKAEBIblecWUn1MRraIW2KWZzdAav
DgjB0xKawW4OIJxVI88YjPx21TeXN+FT7xwBh4xTavaQZbEHE4+iS7TZKSF6WQyU
5qi9lehx2mSukIalEgOEMZQHdOO2iE5znW0Ow4hhbJTFUI1PMDkgalnw+Zw1Qkk3
+aMDfkR22ZLzYFkIgDRj4vtkhlN7nbO1l9r1SUMSuynsNpJtpG4qK82M6nMHCX3e
C9m48cNIkESUzv6xoMhNIk8OaAo8KXbX6xnw6qNDeyoZ+3VqKaMPfwSY694j6aHK
Tx3HtaSVu3kiFXAZuEDMFgf1r1Vucsi9QSZ0bqnyF34Sk+uGcAx3HVLD7Hm2qMYC
4uKuaUiMxREUENfuHWRJLU+scTT17gVgq//9++71GwTW7H9/y+QW7R+p/8CE78ol
Sp9FAi85tac/AhfOnZJ4b1DoPKRnaVsJLPSMriVzYUwZfO5ilRWUYES+SjAlJL0d
NzpJ7o6S8wM/gM08o6ZcXcGkRmIgJL0oX1nRvl8SWFOQo9MtDiMFgxTn0TqA/SsS
/W2+AB6JCI09Kme0a99bIgK/2CWPsbIM/JRuU0+m82r2tBiysEyUAugVg+qPFklO
u/u7660XVSbIUiuKPIM2BJP6ecv8jvB7F6WzfE1KpfjWK+RTABd7QTPjkyXnpp7M
+vvQ5uEY0FqkDm56sdMgPzyJSTb+3FmbP+USxxhrfLRxFQ8gje86u2bry44DZGwB
7X7gjkkYeX6e2SxEFZ5pHvhZQg4uJvFPwYgluTXtSojWScYCEilEwqDpqqlLbu11
Iz1MZgyfTeasePbcQB2iy4Ex32GAQqEFzPK5b1rbU+h9yzUM/Wb29odAuWIJcKEt
4HJXdlVhGy8rONZYu0s8pcJLCuG835JM70zWpLKLjF3IqjksykeXOMJ509Lp/aA0
Sc4n6kZigxqi5mFmoBBrS9GwAA4JLyQOU2PecmOO2BgF05YYYWB7qlisNmyLBbog
W/vi9Zl/pEMGS4BDCqaiW3tozSgNCJn+e48AGKHLvyb4amqabsimFILh1QaHJXC4
BM60VRDri6KY/H1HkSHYsMbPbqYmz/dHNXkqaiIy2pxjjNXZ/wRSaSA5DI8Up4n7
itx67XqbjQbEFM/Lw9QIXGM8/CcLjvmyWyPBGC9/bUmezs/UUbQPUJ6ELANlLfIJ
QW/jewyqnn6lM4OlSNKMp2/M5Pft/7brdXTfzsN+NgyRxCsI6S1VpTzSvi8RM7Lm
QIuw22p9+/MRLczHwvXjjJUgQfaojFcxGP9IU0FZKTt27S3Tw938akEi8xMiUOSH
5qeaxETYT1ay8ovr+xXbgKfZLANY8g6O1N1wLxMiN2y5bJabRwuDZOQkxf5IXn2A
fiJZT3DoIvH/z/8mdiCwHQI7g7tWLgrS8mwnJ1accpeX5n6FeMXxrao/CRAQcexp
H/RYlioB+WLwuXEe8uLbnYYVDfrmuGB8kVqwEQlzaGHRyLDj/1Y9D4IxuawYIoUA
vaymqgssGlGnnTzo8VH9DtenDeT8ZT4IlZI4Fiq1WPj0uZctLLchXRKo9jGtWi+Q
8SE2WL4SkOB4qTkYTN8ymbr+ktUj6Sx/qmGTuQyBBR/IosGWml+4UocIf4dxCRp5
YchL1uVKTBXnROpiJK9Qr5JVvrihdRQ2qexhyyepT/etOA1XLSIIJJ+LLp73SC0N
K/sFAc4E0z6klt4pUlC1bNVU7tW8awAn/Bw22Ww9enN9yJ0qGIY8UpK2IKaHmslC
DZeWPm0vzC61e8+ArJUw9g8316vpLw1wrJgQ0+R2SqPPWu5marB3z/EgKKGcxVgQ
HJNbLsQOOFFOGhns+dws8jXYGintOjGD2Hpb4t3TEkdeID2Nq3YgLOk77dO0tSSw
lN97qj/JtI1HgM6EqFhxVNgPH0k84EbGfHBXrLN49y9EKoaw0P1FN6OdTsP6b+DV
0CGH/GaEBacp5PVrRLAfzeJK5OhhMo6bLq4yikMsguHbKUGLiSH08qA0GxfiUUEQ
sXMwpyGucJ833q5GLEHKpzMmPGwlZLLCsr5E9GQPfc7wbmXCeRnqmszpHTFFllN3
NNp9IT0cw0ejmp5m8IN2hn5SPKUAJuJ9T9E3Fy8SeKU6sAHLs/IKS7O7YX1MPZ5f
q+vpJ76ojezYVDMfkYxV/kzF37ceM30RKIBgdODw5iXDq66Xl36Zy0D99WXm7Z8r
611yWRvy4H2D2Pro3R+ZtbX/Bn+f5SHzVNSlS8MLfapSUaurfaaU2y2xzYxff2a3
a5QStaucEAfKtBpB91nqedOLPLHlPlNk0B5D4nh0pOy3bnhBfNG6pSeL+kfdBiGp
xvKdb9zBbCeuqRVCGlR6K7UTgIpJna9BO/UD9SdfbZVKlwdPkq1/dZMlBMfIrbpK
u0VzZJH71MH8lUTse2BKsjMzKKb4/H3mT0n7w+OIMM3qhKC9XTWJ7eseIWpmHN3Y
+sWhK6B3Ngq5CIBLAru4uDh6+O0rP8AmzbKL9jQ0qETdmDUHs4B8YxzrN+J8Svsq
lB9Yr/BJnULJTcx+Kg3xSpXP7nuCRKjmMhfCBd5ZFG4dLBDr+WX64oy3ICrqopLm
uGqRnHZlynITSObGNSa+HCw/qA35nqYJ3qS3Zq9P1lTFbkkPfbrLBWpi8oVRxo8B
6qYQPgHzKpvpK7Od+mEgBYKWiycoTJuJcY20tTl9XGpXvGj3YDTJnwEZCUEB7PoO
OFMsOpgTrDxPrLqhGWhd+oYTqr8VsQSWd1MAGa2t8cdVtt8sri+5WgejNaYxAz0s
q3jjhUEkgNQDg6QS/ayedj24WghzYo3CodyeQgey0tw93h8hgTy/NND8T8kByD7S
ZkoGKz3YBn93KLw/i4Kj2TMMOZPLvoDSOjvb6V/P+ysrkqPpGnXiEruuOQ3nbUio
LpyB3Jb9gyhxVXSZt7I+lEi+M7g4KD74o/VWVtx6qXvHGD3DsVjeGH1jRwtJblNx
/NsDf7L8RME3v4NZlQKZCUd1K7DvJRjR3N/2MUS5HA5vMlqf9Y9UzXwixv5UUHgc
/3AD298XfLDMC0mvBxTscTZT9vLjn/Z2r5HcCVjhbcVsJZKQ++E039CJt2wzsaws
Cixguq+nI/NhSQAeCFJ6NGZ817PulwY5qNdd5qLQUDF0vnSN9z1PiPMRnBpHP0vx
nHtotLnRREDO4aW+GkDprH2zq3bt3zH11RwG4q/kt5/9OinJ3E93paFZWGp21bqg
N99uA/gCKL5Us37PJK/BzdINpNLVY2x3l66+wvnGJ4uAQ9bCGFuY287Zuqu3mG6R
lKmAkAIlv2fyZHCbpJSyDEsW+QVq17aWUl7kEv3VW5ZQOkOyGcwCOFViOq/AR4oq
I2VmIKgZQbdbZG/mMCrNGS1d9DDKXuZDWe+C0LDjbd0Zv97vioPlEKqrkv+y34fj
7RKXeCmUqT7CgwsLkGXLlKfWbn8GR3hRSkpKmJYSJklZFI2z6xB3BhypRi13K1cT
CumfhB8/w7luEWh2ldSKnkgUU9RMPo3h7reMbvH3091eKxwWtO9tygy3bzca2rNx
qNYfkS0VEfdTSRqCYhxQnHUccwEtJBCyKfHfKSITQUDfA9j49zGC2DHwbrAq9ASh
aE20TJi9gHyz1xGMPmRE7V/VGJCBH1bXLuqYasVTYi5zE05YrYxx6FoYz/rENweP
BwvD7cgCHYstM5TEPSUzq9wpaEuwoXmUQY76s/8rXsLLm8Em9HWKsACmImaAV3D4
NLQ/yYucyS3uvJ9T2uX3UOF9n8W0EJc2tZDyCDx2Vu2TryIdn26zgKPOf91yOcXR
H3GZQeMB1n/+g2XCOM4fl3liFtqFo9zV8BzNlgvc9pGx1mVXndotmRy6QLGROrCJ
lU2j/WAg42/BJ/gJJN0R3KYBUUbBJkl9cd04jC3up4mcYfS9wc/vxTxxVUczjeJI
dgVDHt6HnambElrsBN91xa6EExJKQRHlqjXqu4oZXDURzX9HzYeQPYg+c8wRKgGi
fzIEfEIggHzniaeErcSMrZ5giyXW27B4m7y5xtHYH3+b+SFysNZYmq4ZdZmJOeDs
06dDQdQNCmQvD3y6ZwKaK0+7m0zch6W6o4zX5QgdJR/xQyNVr5oQnXjJhgMM+x19
0U+fAGYAAWmbo5QYb96dUNb5GO0EmgvfDN6g8bmD7KHIKWcAoiJpQ/IPRsmJBttH
eEtDpF0/u1UvNiR41KLtXwCgW2qwYDN39O4NagQrM4dtcemLZCN13LkSumcownaQ
NksZmah4/WOcppGCiHs7RNxRrAC1beFVPcA5IrY5iZ772HFocP1eqOO3fui0fWKG
5Je4GaGVN1tneOtq7QegUTEa+EY6KDOrWutsIav/plp1tHy8pZLvshMqkucR5EaN
bjjBigPxGD3J20T+FTKV2jCXh6kXYc+O1yuH1gxAjf3o6284GTVhlpdn4NHUV6Ut
mL6t2F1KPmdpJTiIfjR9EfxbVLJOH8gizULcTBQWXEbID0va5HZ+p3X2OLQ+mb2T
eXdknAEyzpE3dYK91B6nknTSfaOhkXZ/qgmtv0ozR5KnK5MqiKGX5LIsYi3d9Nj/
UvgzRoR9+L/4uSh84L+oMZoRzzX+2PM9tKPkkrXsLJ6pCP5jbIlZrGxJ9xTBUuYr
DmdeNYBRXRq4izPCN+DHsKObNNoqs70xhNWJd54+UkOSwIiX6Uns1//WduCAkXZJ
LhzlS/SGctZsK2WZ8R0bkHDpq+BvfzIYCWA3+xgOMZkujpq8sNOX/vtkD+6V9xu4
hJs6GtV1ozYYNaTGShhMWNxALDMrbCtTD42fwN5HmpGE/QZOQSzlrM+OtfzbPSKt
nPpeKqfSLLIy6eM0HJAOl0tMUSgSOO9Sld4S6zvq0h75qQg36zovoofTXF+Mmp02
ZzMA9sUReyfl+sTgfR4nihJHZ6bZnHYKEZBb2mxX0tocGyKYiFRmhUOSlY01V/3z
id/CSq2yq96dwL7rEhH/BJCTVpiWn6eOQl5XQKwPFQP+q4DjA6VdK+Buo4C6k9ik
Vu5W/CV6Vlj9D1gnyTXBVHe3qX9W0xDP9Tqy7sljQNuYyosZX8RdYiZe8K6nX1lv
AWAhTvKgvkw3KjkPxN1Ui6U4H3foOfCtBDJlS+xFIizZxkOhwv/q55IcqlDez/Cv
UMyrE/NOcjAAT3yVgEGc7aU2q+Wyli8hPv71lyw+0YwjCrnybQnkqXjbWG6xdmna
nUjgBvKaFS0OxcIej0Tpi17xyKbd2oyrTdnwECTQSW89Uwo/DjRfGF23bx3OePMt
d6WkS2tVrCY614A33LszkuTRimENVCzclRPd2FfL660+rdKkXsIGCzbbdNQL8HWB
ezq0NAtS2dskX88qkMPZ5hkcsXStSq+9bTn/f7MLocGyg2KIFdTgxAQiwKKoxA6S
od/vjUicIEqjKx32Txl7PcYexh13I0yX4damHFISU/S28J8qOwoeom5WM4zRqwbZ
gVoBQdbvjf42plKa0JYWs42sp+1RrQRnrBxNOdO4rM6k/7WHZ7WLbMasoXjUq12X
QyOfcpGr8aSxBPP0DFXFYM0bgGyV/vdqLWkIgZ4KIND9tRk27M3zw+7SY+nRZpWb
GR6iykXPuLmG7LSCcSSuIRdj19j7CLGKpzpIon2oUtdCVxmAekIJVz7RxEGnLxvl
ATnA5US02zQ1aae+YzlYwUlqhD6jLgqAXLPvuYLoNH4Uj1euPtBVLn8uLQfqwqXE
paHwIpTJsoLOur4pNLYu+x/CYz8C7PNjDdYw8Zl2BWlluBpRApSbMeQpw/7s5zHb
ytqH3AkA9qs/otVDW/Mgab+rICQv/6f5Yw/dCFmgZY/H6cHFQxNQBvfW2c3ciO7Y
FFkCRNUwSfn/zmyRBS3QVDux6MRs0SJfNGvAbz6RikhvpVt7kJYSc+UYy66B5jCw
nko+aq8CHwhOxfFP4ohW+QM/pEkczIIxLq0Z4piQnjHnfAcCib4dzYaIJ37rZqBH
Y9b8EZb8dXxdGjlEZUNf9Y4u6X9fQ+1I6iuEUnsYWCTRPcwQ33GKkbtlMoZOCVf7
3WnIxWr2b7TvSRIIliPz7psDbDGEHFSBAs8OFvlecz3remlMtd/vRHROauqNS/9R
+wHlqFjO12q6gCRg22ANXL4QN9WRz9gi/pvjRSHAWrkj8Z4YtXv4o8K7QWlCQwWS
/u120C/aVzDZd292y2FYariiZWnQrjyDhSEDKvpduPjWgqARo6/e/W6neeSJg5wH
1yldz/7rBzxnBJKNh9btzESomord4g4IH3Zalz70jW1OOL0/AYjr+1VLzndOVI7V
VYdg1zh/YnOb/AlM8465qXrtTpSM7lnfMU4RxrMWPqR291uambfabZL/Ig8HAHG5
3Jxy1ohn/MA4lxmWIPVAC9jPy1CiBds4WMJWPscyfgt6TRhcNy/kKu5HxlRLCKGa
4cgG3F+GnvZBw1ZDffGpHbGKkYYltFMUh/aO7DXTObiYSf3P1EauzjAraoIed3JU
x/jvskIm5pjQsAFRzLBlrKoreJiEOGPmeA74I+lc+RxV3XJBCnOMBwThF10R5kyt
pHExxv2r3fGiY6BmQQAWlu5qmF6GPdqXR4zYEaYdXDr6fTJCrlkQh7YMPpc9p7JN
2zG8Cd/WRjn5Qi1WhCnHJrZ3YxIYQQsCdkXVZrdQPBgR2qMcnMlUFqFL2w7JgfAK
XG4aY6Hk4eEzyhNRrFCHFoLbuRTW1hPHr5MyDn2fSMwts0uWlGQbpOB117mxtIh+
tnhLxpM7QWVH3/XNYoDPnduCF11ioNiJURPEzlDVaXg5yxdSdlrfhAZ2zehgLpyo
z7eJbU/TMHuHhxAA/cnAYtIvKfYF309EVju5jYIrEQiZmRIMZQ5sVCRIEVHjCqa4
h9NqSCNa6jC0qF4j7agdM2I+TYTwgP1ErpAx8vPU5No2GbN8vibwajXeU2vBgRzG
kBmOpKHRMYdUMXUP06wsMaaqrj0xEHHdWOQXxvhSUtjwkUM8qDMHm/K/ia5PCz61
k+5CJCamKAqEE2E8obVtTUS59HKKzawKLUoYPmq+gn5YJnjrYupW+RuQsxHA9w+W
LsydY/keg7Eohwmi0Qc9c0HGJNdC18tDSc2cuhF52WZvAm16BQRqXapbhn1C/7va
b5NpfUs+R2VHZpwzGfwHtjUmMVGJuFCloSGVaLAFHAaeWjWtER4wmSNKj57J4zho
vPZ1cepRqC3DtZFi5UN02AQfOfpfJkbdbcjPYaTNu1tN1aZG9euT8pk6uFsNJ4MX
1IAjZgB1ysuA62kCDGiq9yjMXVMXUAYuT/p5JyL+ycjNDRl4pkOYyMGCPv05X3f1
8w3rUF2YZqZY0ax2BUU59DFHV37kvMe/+abLtcyZBnFxSdlni3yWmrkzY1zqzD5I
lw6ySYV7HZLcCoDRAgeU9n9Krl/R7TdWXcrU9UbTceZbvINuypOdYc0JGYMIfhuH
QrgJRczyz31OdDsLW+xT9s6uLP340hXfCyPHid8TvFHxOjySGZCMT8V05M7WPGmg
0oB3PkeXR4H6HIJpgJ9XtgxgNH6LyVCCKxo2tUa124i+rGt0Y7TPKE0K4ik1jAhs
otUJ6l/ktnZDX9uKwYN6BZbxDDm9aDAhpBLvz92ok8HqcUVKnDQ4zkvt4IJOpMTT
JcseWQKLYG2/2HvOnH9cImMPY3lyhF3T9DhhTyCgEo6iMJfRhVNIK17wJ1EgpHPi
xt90yR5rIX/Joy4ECSnzk10fbGjKA/4hTRLvrexNsTN9/oVGaTW2IHrZ2spBLWMb
mS+GL3d2fwpHiz3u/QwH8EzXvrCAOLLgY4QL9Z/o2zNvnqyt0Jz/1gW70Hw80a5a
bXxnETgDhSUE46zpLfcdrbc5vkxm5Wy8mWzNgJNOqPi66e9qFr005J6vyaem5TUf
nScO52mf2sxBjJiievgS2AkzBBjCxY0bwbXebi4lnJ81WbFC3vidIwpN6nu7ihQ6
KQQXJ/VCO5+crbfOinA95gSVBczTbLxPknSC/RK3JrMP+0ugJ2eT9YED1tNlSHVJ
9xmHC3fj9El2/5laZUkq1ujtuoqmUsVSl60Pj9mt5zqaZeij9zsH72nNfOESsmMm
8t9SfI5/0py4vxNQnXHtbjICTZuuA4gkWd+gI9wxFl9ifYQFwRyF333QcqBmgpZ+
4GHxpkEZJ/UgizEgPa8H8QzW9gjIjsYZnYDlWc6nz3SzCRVCNo98CddpJemht6Ad
CqssLJWwdfpV2oORqceBrPjLxpXwsyKog84DNdDmyKxqNOgplEIA+hERJjHIXc4W
iIjIqufjAtED4/MHwC1oOJABgQZS6KvL3DfRzoo7rREx/BtQramWW9XbnbCVcgU0
kZ/jYjQoQSq8Z5vBMoyPutw1zkGIyzHaJSoa5Y954nb3jlNYX7IHveA/W2YBIDkd
tXl3k6YwZFua+iV51VtFBCO0ir9Pa0vXr0o7BxI+3v5e1SGowtVIBgbLKckDevt1
+r+vhrEY55CJdCysruAhmkc7UW/YviJ7WeLvpDRq/5z8OG3FDNGlFGty0VknjeK2
GITJ2QxgbRmGB+qcjnucyctOjg+M7dHx/tsAkTvDZV/goOdI3UY1+gMn/3H52LTx
u38fBw2BZOAvxSu4BHt5YHcuBwgjpZU2g7N5fV80YYG1S1DPgbJvxvQBUfL0TcKn
FWDxZGEg7S6XDt/9E54xhvsSLiNlfDWlec3CAc+Iz23clLNeYGOmyALBiyRNx0zV
NT1ZkJtaa7NBRcaii8j52SR0KgO9n57wFSsz2Dsy/Fi4GpheXsy4FSP1/n3IWlB3
J0TgxY6N2pKnOVTirymIzrVHl8MKW2brxrIqnIYkTKzJ1qmV+bpQ9IC5keWP0KmW
j/EyB0TFUuWvrTpL6wkxzf1W0HP4xSiJMc3b+Nh+tEez9B5crS9A4fxvDD37yk5Q
uowUxqSHThJqMs6bxMcl9ZTiwKXdAO35y0Itncv8emcfy1xTsukIjZdkCSfcuD5r
2WEoa1zNg7A3S7lWPkQKt5b3+DCLGkfZh/rD3ho8l0VE/MUhXmYiWHL2IiSuvA0I
TgRBkoJgiVRyIkaQpypahTTph+2tpHzCK3VMyYXn672kKz4I+7ot5tRAxrP/X5Vh
+AGnd8SjrOinMA4CG587tfA1CERRVK44xuNdeb9F+eOtr8Z9PpDlszKEIRvZ+ZlK
4ZABzKGfDxO0TVcWEW/TkhYx8JXxF7AinUD8B6OXYnxoBceCDG25Z2MbKW6aHKo2
qyM/eFc5poZ2M7iqSTmc4gmJOds8HjGF1DJONNwrnF8CKv822FujTfyzmsd6Dc6A
DlRQ8a9PNHFVfQo30TWXfsBRXBUY3pnSWXmuzhEemBCs0jcqaKEwRioxpsgq8ons
BzPbAAr3CCf21ON3m+VqYFwQxJ0ZLX8yhgbI0DUtpD/vYNsPAy8nd65+bXk1AGG5
j5JrNPXy1/W4aUeXAxdPY9/0UEe5W7twUzEYlE0bdNddKVuXpoKw12aomK2KQjvG
Bh9S18LqIFKPDdIEAOoTIjlZNk0IooYQRqt+dBzX7JjP0DUl4CfsBc/9H3tED3Yx
+IkRRB3msK3Tuy2NI0a8P2sxAdVGVSz9z60snR7rAJz+F9eg8KY17LaNvdYyEQ4j
2Gb127EP6o2FfML4fPkpLPGv2jJM5xYAgF6XGkzi7i0XgFYVCvABvNP1vGTvGayX
McOlvlWNnnVB6qQbBBXP4eGJpAt+twpuL7O3WOtMQFh4Zz4ao+ZlnaxFMHPjgOHV
JhTohsmoe+qUmTMjVAMtIi8BQN6xiZ1lbtcOpxYbhSPJymItd3xbNvV/0oOgMJvA
ROwhcvMLSrHKoFMNxJsP7FVEZD7DmkVHPYamkruCczxVJeSfJgrUaqrstgk9f9lX
Xil2l8SSZrkDX6MNZgEt6nPLgk/BIrmuINKo2kO8xwy19gPiSor/UsLPQe0szzKl
57RkUoV2pvCrE2wH0wv4WIv0gzgNBdUxmjpYPwfRcsNq+CcRfgU/UlyFR38DKphR
WuCP58ZjaZxJ5afAlf9utR0ZP4JkQBLhSlL9uquBychz4VH6QYABj8x/o9+Rw+No
8EE21OdWGGRkND2DcU4CT1At/IL/ZTpyCU/xeZ91BjtNY07zSG0Zy4xgUbywKthN
qlWoVc3cS/w1nxYloBxgqw4eE9rM6nrGx2Q5eOyf3FzSUMCVPukU6J4RGC89h+ZS
cr8fxFla5sKd3whOXfnVhTzKQyhGNZc3wSaokoRHvIQczNPiSMwPOUi+H21YyTk7
IiJx/qUV10hPtub5vAufvuQK+rIggl3xjQi1XLBbUwda1V2JbRYS/2nqAvjoVxpV
bSJ67OOV6PJbRUuywhmG9pM03eM1eWZhkXpQsJNnieaHdwSZJkCChYhZ2LfRA5bL
t5LBOqhw0AbmXyerdMEKzwzF9PvEMH5QnPLUIT9FuiLYHxoJZFoqyoLEYQ7EIRgW
+FUuSPtHlQT0Lh8B1RKrqEnmTJeDt+4MDG2961K9m7Ppz0eWeM8LcuD1l/ThOenI
00P/engLS6s+qfD0IpFcDArVmvReHseZxxMYCjuXxiyKag8Fy12N2vaAv5dP4mI4
vn8Rs6X81DJnhDPxrs6bO/kJanIzbZjPq20/ZBxtu1bfxsGJRsWtil/UxPw8JZ6N
pi0s7nrHmgP1gwygAgiQo3pE/eiHBofT/39zqqkTKansGNbrQuGk/SJHQ7gggVw2
L83o7+NYdMgQleO6I3lQRc0bij50i6AMNwJqb7nyN79PS78S9rZHWB+qs3/KtQXz
aQ7+m4UV5WKmt8nwKKHVlASP9qxT6HzFb53LLci+hivr6SNrIy1jd3nd+IbH6t4s
FskAEKrFe7/uFhBTIvX7wbSOrzAcegoU71Ukl6ZLGTBdePynEJZakeR94XyaFpgW
RKgzByq4bTtcFPFgEBdJWQ9jXJh7ZFSohYNdbZSDnjIWUfLbfo/ZOLAVV45bZ5cc
IemmkwUDjdbt4q9/EC0IfumoOkKkNHEg9Nm6B8RX3K21wKsIrQwoaaHnMF67PVgY
X9NxyRZI3ykAIaNFkDPpENtrOyD8Hd3SSIjRLf4fjY3Wshrcv9xXm3wFCKKgC80H
YDo6xxGRU7uTQYFdJcOriYgjSNw6Y290+a6ILDjmux287kU2fCA5BylV4g7aBm2y
KzVspZcrH1RHqPbj7pTxm/fNZvYkFkLQ4uNEXcEEUp0CXeKREFZzc8Cey9T/mDnJ
1pOPWZi+fUP920vmYe+aZn9+mRFk+B1tGbdf0f+mEUokK+uZrOizTaUOZY7+JLuu
xkBcuqlWFsJnWrA6o/GloHBs1QIErMzKImvS/VhMF73fLmKfzTriZK02iFQSMmUw
W7wzWnbxU2ugOSlU0EKBD9UWfIbrXqnT8hfhYuR8Z8qfyUdPHa04iAG3EtFAKX5Q
OlF0gI0ph2OXg8/P0aTtTMl45SrLPUHnGr6eRVLw/Z0a98ZJb47EudvdiUn4tTvT
vw4U58XeFxShEhXCmfzdiQZHFt2CKhXrCN8k2KL1vIOjULPp2StiaTbQjO4iOw6h
cc68JhxqOD+bpI6ZqRU4BNeff4QtrZvxPYnFv5Q8BX+yjpo8PlRog/Sa3pv8Dre5
oKwfNnHCDZYexiHlxqoNk4GZ0y48wDHtVPasoVojdFb/gPQynPAJP4HFEMDK0PwN
C+ak38JuBu71ZHrIy9q9FYxozK2wMyKeCKPexOtttDizMlfFTE1HgJHynZpTARtP
UVAuUsHABOobNq2RldS1SlZ5818UEvOCrbbjCCDSUYOPzKARjOfMQMPUYLLEUHeS
IyH6i5A5vCmyMeahkQZeOdp331eA6P6LFJVyqWYKTSnD7z/wMECoKRsJdQXI8xQw
whGn95am1zWlLUCk9kaWvY0TGtL1hMEsY6RmVXSpXbPjPBpheBqoVlHudznJNdkp
u8m4qHn1/9VDA74RthsofapBvyFFhLFZXcgZyXUm0f2vSygwoRe2HZODiDuNLfpr
Zdcb+Ml3Hr6s78IE/hIYLyLl095q5AKLyM4Q/lrpZ5JyK7LUb5ZUbTOHEpxys6GD
GZKNlo35asyPLtfZmLy9Uslk5NfcQloZcgyOBWnvJNpoPPsE1kbSXe4yNlWWCCgn
sBELMnx7dqC7jYnm90zO54LFdG4ccF11rBiiw14KV+/DEsBYIvzfHVLeGWXXmWtq
9r5ItNEHKOtkwCY7ps+yXKHnMZMJq8xwJ00uh6fG+8OJ4JaMM/hD07CbkInGk+U+
4C1bKZ6QmCWijV7JrhRKoQ0D2uHpwxqxAP9K6SrPN5t+C882zUFSm6dKqR4FMYx6
4qP0BCWuPPm3QiF2tO1c5orWn4jGgXWQN8Hu8V6mBNG6sBvUIZXC/Kjyu6ATAI3e
zB+Gs/34nZHzrAASHnkL+3xb5gE1kys88jor5qnGtG5TQJ2VZ/RqGNa7Dy0l+Kqe
sNFmUy3618Y0VEMht/pQrB3mOPB4+CeedNUHHDuPoz135mbviMMY1ZiNdCE5BRlV
bitEuCfm2fzK4k+p3HduXj3QSXDibDtdF7qwa4ZQD4Ha/LbP+AhiWYRuZPXZKYwR
E1ZJ2GNjUkdmRfgRMHLtfUkKyY6SmCcYYHSlNvcpvgvtlFIg2Nj08iwXNUGbnlrA
FNks3g3TniM89ZQsvYkElmZnh9SAVYAmSt81KcPOLWQG0tTNwFl5HrfpA8y0t8/w
Qlsf0Btbh6M/3EZXIDjgIOJUDVome7gnageLanhh7ce7N3e670WsfZUwQ5CPTH9O
y0SzFUtAvxIXAzto1aOQvC6dSAnqV6V5dH2ITFL8pY4ATBnG47bR4lYZohuPMXc4
8caofZvgZTzxBszlzStEmALRowEAa5DxbCajlmVB2Tpo1cWwHM/eFYpGnpwIikhA
Qf1OzrJSG/GfYf3h48ohf4rzkmImUpr54cauvp3pu7Rap8kHE454z2cegIuzDVD9
W8RlaoI4X4t3oHzNasI2YSXZzQrlPgf0hhWj5ZmpurtOKFT8yofblk4gYAwVchk6
nkp2S2p8qrjQ8cwiStmdrMI6/MQ0b7lriubArbXT5LjVeiMGFmWkjfUX7Gua6inE
e0dqsEJhTkODym1Va1Fgdx1/3z9Q4pi2okxjDakrH0gsRVqwkSKWVCEpDFUXqtcf
mjGGe+kO1wB/I5Ua0ZDraDy7fkzH+32T7vfPAOXV9g5xPKizhEq2rNo/Jl5hVQbY
fdsLepoiEoxLaCFa6mMQqG6HgIYgrP4GoRNWDO/5HoKjwVGQpG3QrwmtwmiKVook
BvaltMzqgp2oOkkTagimseZvsM0I5DaNzDJLAt0WLVVry/LgFAthUd5fedAaCrA2
BRD07SjkqrJ6VFpQW+aDqJ+EAvFmiQGLr3NKLOCJQL0zA3/EtYvf1agECA6YHE/6
NI/yLsfU1GJrfhjXieOV60vRNWj6bOQi+d9EpXlG6hzHWVp7D76DmiNVrymmhZwz
RGO5mE4BfmAMlIoTOo143QRH91B0caSk7CsaQoKhi+5vWR3MesdNIv8cYAd2Wrcr
zoRVALm57B8/MYcCQ+28CskOxO7zEaIps32ydE7rnlga/qY8hFNIYW2TTczwmLco
kpFrWLXbBCm7eKsW0VFkBzATBPbqWhAw7sZQlZlUlaOVzpy0c9Z6BXE5PelrxR9Q
VZdOykv9a6cNfTLWcVwUv/Be6w13zR64moThQMw5mGQmf2b/LKk3D20HuzWfRcZq
G0Jf0lSmZxuEuW3RzDMQmBGsW/Ob79lD1tEVZUGOCHN8n63tHVyUtf4FWuynShw4
040Oq4cxpC3g228WP2Mjff81zxpfuAa8Ft5tBrlkWve48OPrUFQndaDfFpVpuB32
HG0gB6XFsa8laprOzd9jdNKiEwH9zds89vM6kc3Iygtxo1LRBvTLgKVTt2gG+VQ9
PbxloKCzo2DQh/+kiWsi/SCUOaTVt9K9MyURHuvZozCcHwuH+P/7E4CAYYLMpCJx
x7QfpRGql09ErMX1trppLV3eairRTRBHj28sM0KQGYPGaMPwySBabr0/Iaxt8/lP
a2n16wj32N4XNIfrgp17FQ5xkBTahAGxFacywRl0ul9CLhgM9o32ZwatN1foa1uq
SujcqxQDRuNpZldYc+Vzj1CBc+CBaUjSIkoOZLk8ypv8ZqqFU360PS97wEXfFd6+
opjKmMZNd5vb5SoSTlVKYKY9Yrs1ElFlxaEtMcAWlaowy/+WBRODyy22t0Q8cV1Q
gbPAkHg6Zm5XpCl5Xyd5OwWd/Fl2LFHsUML07z3fUuiaLBLgqD/3OWov1EdoAUGg
itbX7Rxw95FCe+cM9CTpwHmRvNQbL4ahV0oZyYSM0ZGOE8IfZwqO/2TFbRBmjVbm
HftAZq+FynXrqyXPaeyEZmmKxXTvvKBsQlaSSzuF7fu7nHF0yDHJizZia5ReHZ6l
4Seuq8lnuMbBeuZKdS0oDilaVRsGo1U25dnps0RGMit2ySQAfory1HmUQSpZjAtH
maIYqzAMXFzu/QtbmGlJxY8LD5t28/IAhhez5iq9XD3b7nXt4v9cSrBIPAtb0aAb
nFYb+zR+v1cEc9werKgM5riEuA05Zp6f7v9ETPKLcHxzPEql2u48Psg8FLtjNW9O
3nupwWJJ8ec2CqQBFKVGzUrOWqNlOK15Ygdsa+3tNaNCK7rSdZaDykNhPOJoD/Ze
M0lMD+5eSRG7tyIOfG+G22NhVSGaCwGDVEK+FjnCEAYHwoE8df7FmR+Eg/Nzj//n
qmvbda6zEA8ZQVlBBXBkOhlvNvfL/LfjqZLUaFMCbvDnsXTj8p+kmHpyHCXixu+w
rvigvuhkevoIPHiDL32+cNlp7/FC3OFRHGZP46GvHmjG5oAxbYSIIf8uLtVTzsLZ
XRgfcCPp93oV9gvSOy9FJNSD3ufHXYgKCxmjdq+oB+Gud3ZGq8X/QFF/IaNfjmK8
VzXSw+xQ4Rumsug/Y8Yvwo7ctsDCTARZKBDqs1HciFE5PWFr/PPGuCYvt36Ozs2N
abeMeCBNLO9vKrtgd2xZPyDsBr+dRUNzsjNBFM1mz0v6PpZG0/vbu9i7pBvf6j+y
F3M9l55joe8Y+2IjM8z3vS1RUnpKIfLpc30uWsDnAkycyHPdxKGJNo2A1LWa4/HQ
fSxZEksT9nVII9cfbsuLMwoIsfSSrBePvnspYMW76QlWaO6mAKt9CWfxVoHmsCwY
towuttVBA2G5oV8sRpLi+BX8NxKEiUolTEq4NI+C5FcHOrCTZd1Kmy1rQZtS4v9k
kJpZTaICaJ/jQZaX+Lx4HrsKxMygM4H4oo1oxi6aaADUgGywo/CXEjBRCYJPT1bF
CCdKR28xuqmuT+RhZR7EkxDnCcOJOgqKxNy48QSF3AIyPXVm3OW+uSxZLSzeq2CZ
YcwGGYMo5YS0KEAADPtDw2enmC5hoDsZQnQQv/Bx70Hv+zOIRomcD028QjkWnaz4
HYd/HxQMSxwOXxRQR+BKFIGITerHMBC1jvJV5DsATDNNTk7SS5wk/kCjjXSOewV9
f/AI2ffUsmp2WSlcA4Y5y/a5RJAVIavzPLTyWcxqwTYsmS8/I2trSYChizmXwDJl
RKgWi73nDI+ZNYRfQO1X74Hh8wVlFfL9k5Owmb8+4fc648uEG4PxNOS1t9qWiXgw
on5jI72160wqW7i0gHiZ723zeh+OtdDSL+bgIUupxhUbApeQ+kfaGPjLMPCQ8liO
t6iwrZAfUR4cpMWqeo7BkGeIUki7PudyBOIRIMu9z8DtcYyAmLNEjgYtBp39+NDk
stzsoJFTNQ5vzzj7gQ8f34D+tX0N+dkYwv4phsLulUCtmZI5xrie0LRdGc1w9X5y
t+rDoGDkyUgvnwKhYb/ZTuZXZVOwVqBDOdUSUyWdQiXZlJFP2GhJbc3ZCIv7gFK5
wp9QimH+vmokwePTt7QusjAoEeRqJ28xHb2lVzYLkS74zGD3gXH12jmJMWuuJtv1
FRg59DqELRtFL6axWs9IqHD6E5cUzFLRA3+xOT4AM9YRkEih1Uihe8Dun1h6jueH
dh239bmbY7bAaCYVOpWNWW/W0qF7PzKU9bG2zCU05yVu6wqoTxvpWeemaHhN00OR
mJanrg2MW7YLNSKIox5TUu0oAf1JfTdL/xqLSUxpTlvFBKz+makCPTpKwjS8q5MS
fjdbirmRzkIjWVxv5HtcyN8rJz53tU54X0vnATH8lUgg2GJ+r0N2r1M6WOcffGOv
KteAVC4V/PQimOEe5iL6ZBO00KEHV12u8WjQqrv7Blppai3Oou+exG2E3Ks+Knlr
40aFd9kkVriL2K4nCLM3bA6qhe3PLOZZ6QArGMdi9sBQTKuyemhGLcqxtDeSXG3t
d+ZgNX1zUS1y1DGWaTONJK7Hqw87nRrCSItMdWym8WIJcK8eEbtUafkWFxJLXLEB
dHB1IyeY0JbZ7AlH22QZLOsvCsWKINf/b9etNLTht5stp0/V3k8dV/9De4o17CJo
UwOXonURnwU7jx4o7vdsp7N4CiifUCtdB7Rk4y9Z9euWUbgvJ/KbLIu1l8jVDhHO
9q4ZY+PDCMZCSHRwXwXn0IXjQsa+FhUHGHsKIGaoQSArA8FVILJj9ee4ANbgLub0
2ZZDR+0D60qhPY/TTZ0W+V25ILSSX3mV1lpa4aBpqnSGuN9jmmEKm5NSYsSQCXq6
tlSelVCh0kG03MGaLLwlUs6U2ZXwpldwHkgPym1cU1+I/we8lyF2tpCE7KGJ2qFn
O+sLmpyqQv2n62dbKT9CW69wf+6sbqUntDBHjol15nbCQLcmjiTDjyxOUEq2Zejk
SO9QaTcaY0X4IvHdV/QR/TqVCb8bSr8aDgq8JnyqwwWZNUTt75VE6I5qwJd4oute
2knUj4ojGj9h9lAuV9zmz8UFWZ/G34T8IZK1Q30Th6ZM6BWi3PkdG9+gUY2MTje5
w52/Umk1w2PuwtzdG8ZlNG9661ydHiR0pgdzTQMneUh4i81kONEUnXGAGUklfLLc
U3RgcmDxpKQ2+kQmQTx54kgpXBCVx9kh2nMeQTdBHCbDf2HDebZB93yXAD3OibCL
kycOU4cEiMxlMAJHo8iqcyn1DevxxTL51OQKZnDidjOuyb0uW8IuAcaDRbMkkDGn
EJvkQxiG4cl+n5tn3nsDr+8uy09SdzIInKg8GJ/KAUVJv7ApBRbZtWZ0Y79/uZ1R
8ZPFMd+3KgYnXA3K6k5fw0bBAXHnNtXRTPjgsMzOpxi1X2onmi6bm5Z2R86woSOF
an7Qfxx0kQoBgJCE03AuDUCF3NnrcYAxAmMrlO624F3ZTrFQftzPoHQs6GoJLGC0
hhjtQIYPeoTwJy+nZvKHj/GiUbfyqCnuaq02WrMa/2cjMno32FQaKI8HX7paaXKt
2b6q5YRIj5iMTUqAdOdomH1a3jMyy7WkD+gi6GAZBO95k1/0nNKrWpuVS0SGlUXv
n6skP0Cd8X4BlumE5Zi7NL3X3OM5Umhd11bjKFlUE6djErYPEzM1iXjw6BdsIQpB
7ZMQhzXlZBqmL1vpGL8YXv765e5Mhk+Kj8Tt5Aj1jCq/Qnvj1572X6JeTrxnTeMz
oJvuR5kY039R+k9gc95rrqBAS+Pf8q6Vhd/RYdHe/ha5xl5VvNuZzd4vYyvf9VHF
Ib+GicSYDuJQ1i87r1OfSRS7sOcLN1ekdZ4ZYSnXkds5iwD6t98BhXH5od2qsFHQ
9MmjlYncwqtjwUVTf2llXAH0fmNJ00LEHgVmoUUGJP2Yf1Ncg6eIy8NChw6Y8+E/
VlHUlPVd2Vda3F0iUUrxpdcwhrh2od6q52yWkNt0YZv9uMu9TWkZAKaFpuhDXpwb
9lTX53coanfmQkRsbD2qpPhEzrB18yHve9A5iho7RiZ4YiW00L5qVIUVyOLGuJI5
YwZRaHRYh8dsUf/HbBqGoO0TKUc9afeqmvkxAPsynmC/U+z9Z3SHa9CUoCrk5Qwg
yZwyyqyaZ9Ei+LhDIw7ZgTnCGki+yaePnXUXCaH8aKrpXDOcd83EoZfGeGEjNn9E
IPWtL+me++RyHHD9XBTcYctY5sM4lb8kM9dpW6zOwgZ1xhjvBFXoGizkvziytLfZ
E/Pv+MZc4oMi6xO7peOh810iWSwpaJTcO+awhr4U71Cs7PXpV+WowwIFwjc+02n5
u0p/m9bnJjE0cVQar0D8j0p64TUPjaEwnLOkPXIXfGqszDFphtmF9oWGYm5r2G3Q
yFYLiaHB0VS/5iviwmtue9nusswXGBtVq8gv/b7p+GR8uBlv8w4m0hVq62JQkb1I
bhyNa3W9IgZ75aJtiZp1Fp8zOup7Kz7Yqe+KDlwskbcGn2RTLOR5Wp5WO3RTT4QI
wOzSXBFZAI3xAy+IttBTqIvc874X4mFuIIT6QUO8qGlf4+pvhS7szjQSsxdiBQk3
qNQpPnOFZVc8iP5/C4zddwrdqSWX2Q8pRChJwFv3RKq/mOYSBjto5jYNpuhcj0hP
WlPvuyaBZyr0f7AIjQcTe8r+YP8EWK1qUWsUrwbI/53WzBR94Ni7YFhRN0SCJVD+
UDxNtgvK2AX5rlC6CoSP4qZvKh1oNtT81Sh3LmcXJm7AP8402xkb7OdPm29w9Unm
6GqqMi99elKj9hSxmQ+Ay1x7XTlOsDeZ1BL0Ygmh/yZQlY56EJbjgqvFy5BLd4iI
QcXTwdO6CV7v/43TywV9yJrSsSOz9e88gN5tekn5UCKZH5qsblHbH/4Tl3nZMmyL
K7di72yIC3Mg2gtiFBkMvXV5AjC3nVUUMJb6bReIEG4+ksZWHWKBSeAFbI1VMgga
dObOKhy8rd/RpOPzUevS+yOOOwTdouWCWVO16TMNRjZfJ9eRpiPm0b+sOwTiMqqV
H6G4L6q5MfBAbNabEjIAV6jCR6Oa8PP6cl7ZlOfEQVzKj1a4EfiTntHbd/VgmNc+
Xa4X68S/A5ddlJ/pnzOT7C5HC1kLJ6kfSp/vPpXbHTUwPsmZZvYGU9A8D3vOK/er
fMhRlNSGpVfFi5Wt2vhlzg19CMxa3WYRQ/vg5p/SkvBIL29CYu+0fMDmIb6E95+x
c2N/El8yv77BqY9Zpb6MIMNrNmbFwj00sHknVG69UZwUNLRn3ilC49+rwlBRBBek
djpIE0mWPr+XDyVtFn6SWKv8IaVkbrNa8q/x2z1s906iafV7MkdmmsB9iio7/9Dd
NY805xRqb2fBxYI22BZyNLuxlB139NyQl/7pHkElvScIEUj0o/8gUBWDB8I4v+v+
M8NIeymG5nsFM9peqWj0ErADYDDgGJPH0ZO9JfuGXGKT+LiqMprrOz03oGbP0dPF
N/CBe/OyRSjnUF0fGNd7ro7d/u0NOJtnordAULMzvamcGKkgdZO0c6KgYF4T30EF
iNqnlORN02Fhd7ub5KGBOU1K1hv+2bAcxMoxHh15mUmfZhb1rsk9y/3CJ8ggiRtW
PoLXn4iaRIUMNCOaK+ciphgoXZJtCi0vrLuV61N801T1Pnlo6mEfu0xN+D0c2/oC
hrjei8+96acZIyDe419LnvEFOs9fxcikF9hSucduMgaFNYfAZw7FkZgBp0RRkt/K
n4jYWrdYE9Yam7hRD/E72lprWV0vtazHZDkXFcR1cg+RwCV1NE+7x+dsuC9KF+QW
6sOFF3UQVAiFVtERYC1L4IUTuD0h6zfOmzmd3DQSxHFRgjrbZbxyVSzaVMj1ENr8
vyqTb9+gq5hSCd0JkN1c2zjJaP7UoVyTnHr8haZUVgUuHodYWVpuQuyYJneKGC9r
/n52tzUNjAFR+Osb554leBiwwTyyLH/yTTh7+iSQiSBP0GYMMvdJkpBZRXJCWjwo
lt/j1MSigj7v0jihKnHhCLLoGwo3d8CuC1bMK+LCWKbOzVN06HVuibSSDAcTx/bw
x0hXw8AA2lf+PN341ZpPlKhQW6kzztfiIIhsHPwuChArwdIkhw/qZHgAwA1k8lFN
j8XJDbMhsjovjoay2+K6UtOlA+LLnrDz5JVnMNYxUhAMZ65KtISkX5b2UBcRot+T
vDS+WL3jl1SUMYhTHzWiC/qsMWkKy56f/JQW2+iTsQwyVIucsibINRxoQtt8VAFB
d/YMVJCcgXRtEg2jXQTESyuvidSn6CZpWcJsywJtHVF4uuraWusqNXUHLWlwar7C
fSYOwMhC+HHSp9zwdVQthWMpWUgNWIFMp6gdIAztYCozyN31E7lR23owDJi6s+PU
gOVgOz6G6c0Sw/aGWBcL5op/UZFXNN6SkSAUe0pkxTR0Co+wbhpPYuao1n1irS+4
kjdmdSp5dpkIhOQJwvH46UMb7+qpuC4ONjz/2/r7AzxpJbUtpxyuoi8VnxXpmIG6
p6TYbXApUh0gYRCoJr7a9CmDRdvimCavvaBCH8kL7Ex7s3lv9hmJW8aSBrI4LwHg
Ot9QMTxt0FDOpcZbPh7/Au1aMnmvSlxtfVu49gRZk/6iqDFTcUlgmDC1aMl/IkLX
Evc9NMAyZ7hv8s8RWfk1a7om+FFo+eu5G2jpgupkzwKahwW6C7OnDFwQsuIef4M/
bKJR8OES+L9rI9krjZhm9KF6RdHQPSEahgHudu6k+HvI11dcn5dy0WqbYGhL/9yw
/jQNZdj71f9kHNPl34TKIsrEuul9FTTPum0DuB8Q5b8PEPDViiuhnxGbgzlS+EGx
szx8+ERTZo9uWPAbWlv3d6BdUYix/l+8nvvFMNC6uWvfNhtVr56WXkR4wH3ucKqk
rGKWzmwLWUn4hjt34fcK/TCyVVJ+iRQgkGx+gIwp5qS27tQCdexe5aJ1jYfs0WUO
qhrqH0J8CzuT1+ImDpo3jmV7ODuP1/FkSVKATJwgcBebYZKiB+WD3jitJNIG4zD3
GkFLK+/vLBre0YAHCm50B1a/lQp2DrM7ML5hy9LTrSEmkXHMlCy78ZpRWKX3AISb
6AYW+ilK6TtLa6muWCeQzC4H0TpRVfnNLh6tWVW7PTVUq272Q23bW+qn4xHLWjiV
thDuGqTiUe9zLfKag+fjUuMnPe7dbZmkdk0MLAZRi6m4FbUqR/m6iE9oq04moUmS
+6QaLfXiEXG3ag3DrzgbFJOxQ7uFhQcS0WBRI6yPwm//50+J+T9E1fKJtWoIfUan
KqjjuKGBgrnpse6adyftPmNi2asxc+ysmMPEBHbsqRSeng/0OtH/PJ9ynKYVuIn6
19JSfor1CYNNUXjbHatTj2BVSYyxIBSIakxvulEYTu6HsKwTB3raE2T9AlfyJsRF
FirVWsRC5LIvIuJ5mEFPsOvVWJGl8hpqX3F89nbruwDW2Fz7F8V6CCcoq8HlsiNo
u8Lu/5gfGOElpSAJAX9OoW6X1AQR0jVDRMlhQuqcFgglJulaMkBGVo3p20HRRil8
Pi8kiLUGBWnPTRR8Ra+GTnSY1dAeqbuYBBn+a5G2VR6rr8ddK37LTmorJd4YAno2
V2ozj8YZ+iUokpOZJR1jp5HDUrAaCdf9FnL4dxAeS3Syxu8c2n8dp5wgDYVgTKCS
EUAvnPCARhpinPnquykW3rS26lbdmu4Qcp8bCtKKQjo6ljJMmIqESIssrgJgTbtI
QlA16K0UwMkU1Z228Td/5gZAVDO0N9SC+goxRBhLoCygJnc+8JBXkQJeteWrdSZ2
tu994ZNg8P5Y51rzwrvBmb2ddvsbVNbGVaRvUu1wRv/4H7oEYolXFyn7eRx1KnUV
oB8ekJuzNACG5GS7glsW2Q8irLLW/K03yAflt37DRlTZ1Bi/0cAyulFVwcKBhzqG
gl3u6fu4dlSYx13IInHx4c03QoQ+8LNkiRt/FByNroAug1cDMkHkhDabNLcssnSV
GNsr/l/UnjxWBoT2oO9/PpvTmIWuazj98Ay/voZZLkO2/PD5Q40EQEyDXfIeSXmF
bxV+ShcHIq/zt0YZ1Eujp8HrNdatsVznl9JVKwxjgx1hiaNyyCBXqMhPjTXZj6Pj
irAp3CJ5FR3ZNnTfjDgsHKcd89opphrRhnfA6DWT3eHjH4VOL500aLGx6JKz1KaW
ZEetsldtemLTccYoIQCOhra61ZIElQZgjdvcsfMx/DyntejYXSGdZ2iJcjlAYyhB
2DfSVUF5I/jRaVn41dClKkuC+sbgLX0ied0XLoQwVim7pRsPZmbq3sPohSXXvs1q
xOrHDuyMqXQh4z9V34A4+uojNs/sOaiIZcnkor/+Xco2EZr818Ox9lkqpbVLgBKA
s0c8MgL5uCma5z10D+KWr5Oxe2mDOyCIk287YQjfN96Fxa2aRYVWSIFmrpQJAf02
zK2mn1Lk9IOZwSwPBJ3f/KqYQ3V9Zwu7W8W1feCFPDexGlMgmfAYunpxphhZ+Jez
sjMrpSOToi4mmHJIAQvFNXSnjldAegiHyA3XmHZtlLyod9+KgV818FDgTnoOX1LI
T+toTc8LVqjFoTuumRV8rGulRYg2VsJaBNEcV7GBYFsYVEQ/qaCaly5bnWXXUxLy
jXhcKPekLHsahSWUZHqqVPG4AFsggHkY2nS4yOjSPVlRYk+wot+Kos9Py3cSDZ/R
d3HTGQGyndU0Hgziazwe0shMWDvPV+UtbVb3PbdRrcpOJj9j1LQTkR89a3kd0Eu5
sSiwwaPfmK0ApKr0xSmXB1iurCjtZOMfoANj33KsGuMrwlH+bzrtY9odUhnJSHKd
jYtbYBApnwiY1de5105xdl30+mQOZzDRC483/Gyz6hO4af8R9zlyKVIYjyAMg3vF
AUAsXLX1HoWg7PB4Z67JRgiw0vcEP2Wd6JpAJz8OJ0fsCtDUxfikpM05jyT5IHAq
TtB/HCemnBYd2KXMa0xO+oPvXc87FCONV7W2xtgPvgHAF1IQpachmVtTMqhMp2Lt
wnVgU+DA+3Yc0NkIzBQMDmy3o34xaEkesfPcXC0F8FMRnXsCuSjTNYc5qddJNf56
Rl8X7jRIwYCm+Y4Z7tnUwdNC4c/IL1wHJIZouPMtHHT14K0KWAtLAALPOJsR4Yso
TYu+GLf+h5P1zA7OoOth850FpXTEu781biqevZeH/YVBxlp1NvtYd8Gb/qHuktnz
zlXvg75N/SRy2AOnwycX5zKa/+XwDMHJX+uGJ3GcFj4WK8KpbUnKzsF+5hsIPXKt
CFIbppmT3X0sUudxFgu7y9duXEEtGMyzNdqZtxmGFjHHgqA7OP2pKLP+exYBb0rN
qJmBR3cZprws/k0K9ePdvpWJNmcLz68tkOP9y7cDo/VSGEmkhW5Ctz3B95bhYQ+a
7EEn/6wMj02USXAvVhmRuhSHt6794ON6dhzNPnSu5fzBuYQd1AAjuTg8r232K5Au
1CEQFdelsP2chBaKjM1fCX97jP/9JwE7h51FseV7GwPiKKbU1S7Q8tUluzS+CySZ
NHelI/Q8bmYO4R24Rf5Q2t/l2goXEz7pFLYgMb4TqMjQcuCKF+NJTLVTrrs4ikVD
XNYy2xdJPX+yXzclU/Vb3u0GpRw0x4d6Ii2/NJI104ef20SQC3PjZkpim7eIIb3+
DWddZZW/ECfGIg6oyS/yc6E9ecGXur6aOU7QQ1adGkgVCjfgfq1WBacObvx7sle0
Dxz3D3ZKUYZmHSGNVBBe6CDeep4eI2aeqoHcByv8mlj4e0OuEnc4FmDsW7q2V58S
KSOdIFUCEAGyurJKKVRMM+5Bwck2rpal4yJ+S9uInRLvxbbv0o0iqueMrLFNs25n
jWmUOrFz9Xi+FJHCnTO58vm5rxkQ5Bg/1PfG09QVNCR3Q6YfrKMo8Apj+1leKqlX
Urm8a7tTRkJegCZav6jjwMYHVpsoA9YxnZ4NPL66VJe/J7YdI7RixPQwTlA2Jot3
/0GuwpK0wjsdbfs9ZgeThpVaxDPt+M/tUoc/vZ2jMZF5WYD49JyvslTJZ8dWCBu9
ONV7tlqsa95iU2QkAvb/PKRgGK1Ajqfz6qyQ/8M718Ag+ieQou19+lsHVtSxW2dz
9aLHzLkTw384V68qn46PZsx0jb+mzyI3TnNVEbZsvke5zKBuBycpmHfFonFioOTS
vY69bYF/T0syPZTbG66PsQy6mSkS+uU8yqbDZOYYKHaVHntxYJuNP4CDBR8t97x6
rlOicPie9A5LQRirdbB7iAqCnppvVuDgPgGa2niCzTD9D9mQSXxSaEHJasp1J4l/
yiSKHisfgNQs7KbcrldaqpfxUn8hxSMFzM8sLp2S8QUma3o8wcoIAGP6ULIMBP0d
BHOUSAqjmJpa8RKh2A9uZqdk8nrprx+9SC0fJofqrOryuBqxxNAgo1LLpKaEKP+U
jrXeLoZYLjBUK32i23gfh8xbf+LSy4g3B2Puk3DJVdrlLGHW0auwwb9faZfXIROG
E+ECECfMvywOolHDIQWil2e9H5zri/r607BEUADXTwJr7CG4XjquCgTPMfgkVtV6
zx9toCjGHA98TzJ7I8MdphNwt5oEhfaHlx7/y91pXuBokdpAwGuT1+WXDt4AvRCf
R0NHotPH0YTc/5TCxnNan2OSGclKY3U3+l1287ZfzlRs8a5MBFkqMC7TXGjOz+Ko
k37HxC6J4mrlxW1x6hdeV3QkfguzxhMve1XPYGMa8bgzJOwqDtn0R+Ru7Of/tLtH
KpBGl+NZV0LKYjgbGI9oR197Y7q10x4FzeaB9pdqhdT0d+COxmXB7inT9pveTlo8
eHrT6r0kkXWgJJBbOoYd6I1QacxuT35n6NbjJd7yxUSV4eRFbEX36nXcZnPmUC7b
Ot/bmCQAiCM2zCHBz9EFX2y4PIPHPg1Mwm5kkJB85AhzUJSMWsAugMcXVd2Q/7ZA
YuKAB3loHWJU2MHZR7zawjk5/o1Q2oDjQAoYJhafpgdbQdGaOfWdcWZ9l9Sy6otd
XjIY4rdq9V+JaesPae/ImDTbDuSsa412dy6dcpY/nOOVR/E4sRSjdRWmEh0Li39t
7N3XhIV7DxWRhZUpmPr39ZjY88md7U9EdHgKK1s42b6UGYN82n7EJtmS6B57PXsS
hfOxGF0uSIh/gUceZhpmb1JRRfHLttDSXO0QaCl+XElhdP4ii5FjWEZo1nmhywCL
81HYmbTXxXN52lTlXY6PNHMcB085kDKztdnn7Z0bEsUKfK4HsKnm+UJFqboEItDR
1uEgCZqH0ylQP2Eqm7z7nQ2V9L21Q+5Ia4cWjsysGnCZEnnKCQrU7tDW8iq4nTWZ
E0sy7+em6j3mVmCr/3AO6rKeprHwQW5M2cenZiUHX1w9BTrYCteCRJnvWYHh5onm
0H7E3T3zzezRyO/KII6oOJ/jgkjiOYrD55aJhFqxwphoAAG4TBhuhItMKoswi1sv
kn3vHJpeJ0Q3HnAObhRjefKs3O3jNpH/aTX3sgyqIoCFQe5blgr5WO9QFX50VzVU
Oi+OXlQhTgmYQvb2p6dJ51wM2ueHXHISY9vO8YgbiO7SGN+fWzYrQluD/dlc0MkS
jo8GO+y02EhTm6ptYDnvXqEehgF1DvG/8w/qvBCIWjkKMhOtmey/0hzKaCiZhLjH
DCuld8OHn5coPXbR+u7AIzM2PjwUiPuOe/nyVXtxqoAnrt53WdFCwNPonWt0v5nt
vgs1wZoKcjaU7IJ5D6HoOmJtZ9hYKceDJ8X68IIeDerD6JRpx0yj6ShhpwVKHazM
RZkxV2fZWQk49FxaxMFeeQjsPXvE+fTFseWUzNjvFfJWxQdVcHNMVXFkBNiBq2FK
HM52ZIfc49lzztO0rb/a4w8KZaZz5hNBtsI3pGmp8/H3QlbnTSV0CuvBwvOwNvMi
kGsXEd5bc1KixOKUSMO+wt1w9SsQi2kQBMy0jYabhV1qQv/VxE0q691GfGkwQSGR
252A71Erw7tLUyydjCRef7tyquFDobucH9KzB9Kd5PxvpkWZo0QSjsQ979Yvg2oi
XOLOReqN0O9CjRCIdzC6IhRS8zbCVuj5Zz0haFzKT4AZzsonRQxcAGJ+UoD+AerZ
gfW+iOD+bQJdOIBuYimO4D7GNiXq5pl2+9HjMqFf2pGNqlp/PbniDYVJySXH1L2P
ddxfuHJuX0SRqx6eOO66HcpfME3eAFA/LJzH20QUZKT02jiMlaixnpOmMALLAvFX
BERD+oGF5cPxAC3yCfdjPtXHtyNT3k9LtL4rO1CXqoZ2HvjwgyqP2tBu5EtGBK2s
Gnr9b2dOysUCyXWsmR7WZ0fSYLaj9NJcSmqI+CuXHy3lNknn/ZjATAV+tBDIH+8v
lMfRZwtOXZArUioU9qYorKWhBk2lDVXeVEAkGhyPNjeZA9hC9u4w5bqAduF5RWZP
LaSD9jtkL0PxZrhafRtEjEEQ0UCeNuN0AqjjNCjcxKiQwZjw3P954OGD/yvG6d2x
Dhqb06TxUoFy7q4Ew4nC6B8s8dozgj5hALI3XV/FsEp3OSil7YuRbiTp9D0RMyrS
Dts0opEYDdQFkxgQOc6I9yVAErzo6k3x3xuFjCycLpdA9YZGZX3oKjc+DiBwfyNK
TOawGxVlfmF6124j6WaTjN9WJG1w5uXAvgtE8R9pWhRSl4O4oKmNyFBYJ4SQcA+J
eO7zN537G5J77Ziwr0+WmyQIfXfR1VsDayJD++q1G8GLNLCLGwJ7Tbikt0vvIEza
zUlxG10tMkTirMpVfCGVP/Ut9w+5mQ92roIyHfcqa7tZ6X4GU+rP01OmPsGn4Neh
kdZKXjKxXcpteZQh+yLWt8gkkhJmWZ6G1ktgy5IZHNu9dZNtpzA2vodbguCQ2+Jr
Oo/L4asM5/VGThNjqtZsaqRL1dAIx6TW13JwKNUqdA8Mt/T32x5axFnt5CF8FEFl
JZPJI2/XHGsLDQKfY59mNZ3TpBxukwg0g+SyePq9p+R+4mEKFN+bu0nNHU6ojrH8
y+VNJFQKwwXlYLcFMbOSbEegGZWm7EANSzCs1jiyugiscJE1oXNp5tbohSGrnC3f
YaE9dsxF+7pqpbPbwOd4scj8zo7bLHHx29i9nJXPyWPy59AGormfBZULy9wSoWjz
HZvhOvhVrpxBS1dYESMZBrntCMra5JgLLajYJwRQahWTcfnU6FBKvyuJiIPAXgq2
aEXRLKYauDOf5P7PfIKeEVx7XDzvDlt0O9AZYr8tJ2t2zAW8mDf0SX/zbjOIdrqm
36+TG9oiZ/gfPh6YNukbzxjyqYwouax4GyYc3GVn2Xvsr+DUlD11yO2MuQO7vQkz
2vUKndecTTz8N6Wy+FNUOtHYJiNob80AgPcf48Kg44cDKQVM1+yXjU1ecCMfV6x0
oN40AuS23JkPLXZ/Pu+JgmS0dYeTQKR/OG5BpM7CMBudOy8DKG3jaHfic8R5pKUY
4zRaNowqLnQe3fUqDoiwRkUSFyLwU9iKDyrWoHcPMvQRSJI/DEjcrveHFlCdyf8e
DXozD5OqEH4ygtSJ2ZIucmiwxHF1KI00V0d437cZanOHRIT5jxUI3yZt+R085TsL
GU5YAueZ6/7J/rH0qaaxjPnv7e1JKAjRmybcLIfOYPIPd1CJPJ3QG3Cha07MxAPP
FSHfNU4P6a1YG82PGBm8JOWyF/tgz9ka08F8ifJbJRMz6SfIHbnkpsHt0Ef4JJN+
ICrc56rqa8d86eWTxoPseA3h2al4SIM1hl4MEYnJDXi0eD0l0gIn9lXGFqTxFfiv
Ulu4WZ3wOs2Ht6pmEtWv1P99MpCCa1/pt62LvxGdjBVw2U5ryimaRCzuX6DS2MZB
VJxz1LHiHiDe0Tpweh5lMCkK0GIw6I2GRdaHgIvnsfg0QHeYFEpQt93dlIBB4zbP
88Aafsx2eI//h4h//EnjdrgrHps9aAFMFsjFml7lpZvbIRLuVUpe/PztoSKerpH/
n0mvu8noImgXIRpfTfkURRu0ZvHvAdfon4vAtnYv/pP2qubQZpdroHSY86qETHkw
7dZ/4v2K6v3YdIO4NymWTvx1iyOrzmDD3dnOGBeKuU0gk0vJ5iENTuD/yyJRGKBP
4xRvmnQxsA3ch7YQH8c9a4Qc2RuWa9kQ8EW9kxuIc8U84uXMUHMxfLwjm1i7bss/
5g6U3lD4BgkU8gUQr/EO9QwsDfChjmHyF6J8kiOq6M+3+dSYNc5hKvIBq1Wru69n
QqUsSdlDZTawu4GEB3mW1YIVzPSpILLC0HrzQ0nJ19u1tEPT+kuSbPqKH32lSDsp
5ITJqhFk39S+IeoKrJYL9mbEk4k2Cq2RdKd+4VDal0V9fnjX3EQphSOCnhQWGSuA
/nbaNKQvT4ts0TH03hXf1ux3jP6GJqBT0X2Is/e0eaQYacCYtieHRbDeNzktvysL
oXauRJQBWobwVXq0xvTFBOuX+BmLMjdWs0QoUzL6IktOrfA6WZvamYUnQT/Ap6oA
c0u8YWOK+EaI7apPHwExofgFEaTU4EHUVYRi9R520v8z9ERIZZS1dcOAwluIHfMJ
2wILY7pM1pG41+DavWNyznq/6d7Blcf9km4r0ebUONOHwKKeOWRvA13AuNL+an+J
ffIlLOn3HCN5Su2yFpxeevsAJXjgm09A8OhZoKmmFjcoBmXX4S86Lnkd+//2hrzl
BhjlSEn5JpRwGLyVF/u1qCDUkx1Um3n9s9am726WKxZCB6Yu+rAO+dZNqfMRZPE2
cZxpvoQC6yz2dr94JHLqIcCNF8yl7rGQ88oswvQ7l/x+w/XKKxkWG9nfJhQxOKKw
aAy0su1+zSaPKYNIeZMuNoMZm5lLdCQcMWC/YDYUhfqcgPphfMV1q6Yxj1i0IiD1
hyLX7TLZAf/zm93KyDyS66nPoiR9ozk8cspnlth2c5ixX7tRrpT2gsfbjBklKZ0z
5+Va5xeulnuYRC5+1vDUKzmG9dlNuvjswIQ7vwu1L9lo22Q04ECur6OFaJWDjwP1
dT5l4nolrJkPLVrrGaaaoeUkKhO/hgPX+NzTNm3q3Dm2GIOgsrdLl4uy23A6dtIo
9J2qScoJp5Ev+WAIGwEXiAWNlECoh9l6Bo0UPAL21mZFZgthkidN9/3YRjB5xQPL
X3cKiHv8Fk5DWSoFKyEST/Kx8xbewSqKc5p2DvKHxfzfjp1wu8qEZAwgxY66PFjL
QJZBRBImZwkNIFRcai1cWCcyZkfbpn6B8LvTzd9+3pkbmKS9ogVILkbDMDVF4HKa
LeZZGGLar0c9qP5ARBubyqJN1s0+dHYUeyRquS9W8+Sjk9xBPiccIC66lAIuUGQt
7PoJZgrOKc4ruiyLbz6bbKLI4IXv0zfqYqGFsa3zNRo3F4vTOKSHeaCS5riRvOGt
1as3T/OU5wBMd5Q3a3UT37ZhGFb0KrU9U1akRl/ucFwjOg5fDE/j/iwPijz1L4kK
2boHXCN3d9bbA9K5t2YZgmk2w0esUQE4wiklT6jPfDzssSGSoNgCpwZWfNUwXKdm
+ECi/rtmZjjbkyZia03uH7tl5+bOdO4abwE+FyKP2ubvKb5wbGBQmhKGbM6XAb0T
v3gp69CYpJ/QEE9wBl24UaZ2ptPSggeYTeEYYBYim0LLCgQR090KSyurO3XBf3aH
fzt5xP3KNHlD30FRmWYngjLljPr++qZvag6zw9k5SXg5m2owoOU4XTGulzCl47Dk
laOmtxpoku6W0+MNVpjdrGado/YuBjWVMSc7/nvVURIMRcumjOPuRcKoghRcW7c8
mC8e3gBIsxZV7i8vPG8HJTb3L0VD5Wf/evmazFkv0aD3PQf7q5uPnB6cvs/wDK6P
Pn8YlEd24MQ55u2c8VtBBeoz3I8opFFeBTadXHL5/T9jFgmi7Wj5jrsJf0ciWoYR
rI2HcDpkSgfxjKFmPSOxTQodtsmoiy1X6DGDSNV2oPiUxsSvqe0No2joifI2SB8m
lLPanqjp4NyxfH/F3sPYUuFsuShqhs5ubnLzN+Wbf6n11EqdAcWKZUzla8R/eN5C
KRwjzAH6shQeDQP/YEDSEuTw8i4zytNmtHeRHrpeBexLW/t0RNH3Ov+macp8Fdws
0/ctWBNqfMLtkZX8K8SuLPcAV92J0zH08N+5XfbsKjsuvoizvm9jBAsSLVIXP7lz
ZsZpD8BPITlB1+XrTPalsKbp/iiN9409wwfHkNkieDV/AydNI6jeysPuWqbgjwqk
3nBKxkkVWHQpKjeZ9iUuYkO1QpwmK+qPHEb5iVKoTFtB3QkXvm8qpcekWRcGo527
2HpQDcCCn+ekqZsZ/LrBlOA0DtFHZLWDWtMwIDxMN1RGIWQzrqOx6PSYDU08kr36
TCn9aipio+nHqcGouMv0kR+hbogX13p1qhrYXqkfcVf4O9WKoovDJBo2iNOS++IY
GGLpC7qPaLRbOC+om4Wrzfl/ZtDGlsgv7XSp5eA0KUpZb30SCxWXW3A3m9JyFRIA
6dZqrvKlfqaN+xfZKZf83322XE0iB88V0NCZR6iXIohu7mOX+Yho4zdqmK6M/iY2
1sWgV3MXISHjJnKFhOuuQbktfnT8OC7dqTqXlUlxlYYMfW0pbsiKFhlTWl/6WRz7
uuJ6oFY5o/gC51i0ZPsivicdlwLMYEO+Wv8dZ00olO/dZdWN0ZCc8N7HDV6PwsF+
1bIjlB14y7KjOvW83qG4DIrahXk+psuvEW4ckWnPhW1uS+MobEVr8ZKe3PJSuv/u
4Guuwx1JzfjjTwqhQXSazgjN5tRScc3b2e0hS1BoagCmU8sO1UJO43r7ba5sQtRZ
fdNXrFIb+Lfm71/vVFIVzBNOr0JDYacrF5obQPzGfbiAJdc5dykOTlljhe1dhZGQ
58nSoBRDKMXwCY2WiJ8253mvSb8qx+2ZsJHVC+MVjdvtsFNJ0lH3MgjnvBwtotbJ
Npk0oBlT7ySvLB1Zir7oI6SZsOSfD0F+s3vixXL+CIX8zZOKzyLTbu0/axF6OeQx
djaVlLgb5enGOTjRjAjR1DPv5Udu52fWvjonpBYX9uEtaMaZk5SUdQn8y/gVJKNG
7Zxf/OgdQoKVV3WUzhccsJvd3H3tmyH0O4HuU0KnhzB82bFCAzhuhUlZ3t2A0Txq
oZ5Zd0ObyxjHknnxu2kh4cXtOmagEZKymoP06SeXbPSUlwBTsP2Pz7FaTpGkBr7i
rMRLLy0A74qDaitsfJ58WBS4JxLuKQ3WLpxrL0HK5p/Bf9XfGQkv5kwqYk9Cx9C3
7xwVxjfKrilR8wBpOYxseI0nb6tYV5AvWZG/xwZGHiSxBIcPP9eyGfJki1zFrWqW
W4CIZHiUNjLLphb4RWzXAgvNSWaycJGTnQxB1SHSxipzZsum7T/bFZJ1b9+qXruF
f1DKiwueGQIWE5OoJz5DOqhKoLYy+c7zXFImK8lw3rl0fzX+ElytsjedTHEZPH0j
1MJnbUq8sSn48yir7MJTwy7rLcfH+w4RAdcgrb3B9Kp9eDFpigcrh6U3OSUECxrB
GI+d/D9Ga4KTEsRW313a1OIMVtX/Mea+96SrezB5HzGYN3wLMXRw5mp8OdJwp7v1
HJgBM+WwwFabslz1x82S2Y/gWDSGlIPmYlEDhwx+aqJZpoHxbO+NwrLbVRzci6Ko
Sy+A75/dB/NB6qnEYOPZS0rcc+zFytIetEoM1COP39ZzGCnL2uY7HkmnJ34fngiK
qGGYKvQXzA0FrpTWP7J7OPCXrHMsnLG6riypo+6aGSISAu4rMgSqDOXc+scfukuO
W3Rj/bgBLvyYgFo/iexsA4b45nnk+iqN9QznsKDHqfcr+tIx7b53bmEtOUU+sUtQ
ukkQMfM1nxO8YzXzda91XMt6rksr7w2/9s9wRHVJsh69e5XuC3g738e4Yw8RoOiw
EP/jUZzP9RSwP7HEw3PfF6/6VYvKppn0vlc8HCrqa51QBulaknQIfHgrJwm8YaZ0
CM0FKcF77YXI5cBYWQRTXCM2Oc7DbuHi+B4hfKlJbAi1jntYy/dda5UIzv24HdCE
iB1KK/dN8Dn4sPwRFPDvCWmf9IxXeSEFgmA4Tgc9wKFXj/ueYoo1U1jWZWUUsciU
D2mbxleEKyxB//V972HmTPiF50sFNAVq6db0yI4Udg/fvmWpSNptqeSLAqqaeZrB
YsuvKZxBmjuKaGwlN5WaifIQL+7piWNLaFhX3tdOOkAqnf6ECuPK6ADI4jlTuAnj
UeesHfbT+wo3XLe6lIfm1x1b2YIZeqmmznh1S2BAPEGxmiUXe4hu6UEbRZV03GEp
UAu1t7sDFDJQKmUorrc1uBrvANesLW2Y6K3BZbWkcLeU8uIneP6MIToHJta7H5uH
o7lCQluwb5niFaKB25vxxhA0EFA78/g4IriaLMot05pToer2Azqb04nY+8KPy4s3
yJ8H49+AS2037Mz5GAi0DgZ4lh/Br/5tm5JKiWJHkJXws5F5szB7FNxVKseJbV0Z
iZyDu9UKV7vrUwemMZPPEYfujoMSm5y0DHqvCh0WkO+ZGGNKcJuocHL1wC4uPXgB
aV9wOVT1dDH9OX/0excfw5FrKB0UMzv4WLIqDW1LAdzBpVzlN3HX4tp0GbsHSI+p
+iZIzzfjUZXoAo6P2sKFs6FCaZYenrUe9vUY38lf1w+qK4j48sIke+8xQ7MURyt9
j7hnp4Q9VtL+GPTnUhijuNNTZm6KYCNMlWuenBxcw0WN4zab2ydFqf9987D2pz7p
bFI0NQHZ0TXDbpiYpazi7d/cs2x97h3JjfNU05l2bhoL70TV7nlcG1rcFLy5Pd9Z
1ex3TB2Z0zn1e0l3jvYdzPxtiuMCX2zEOeBPtj6d3bSWf84AsPSvrFSTHQ0p+f8C
IVv2SSLVS7F9YSdSz8QeoWgdGybywX9+sc+F4a1nLHldON0OlOClUT/hhGY+SDRo
3ytvJ/9VO/v81pLEOsCfqA/d1iK21Y/0ypIbD348I5kOJIzuG5kKuhdxeCFjD/RC
0qyoOinfBe5Wrd/fHFB+F1UHvk1aYxahRZRJ6AZhsFP3OzdnBFgpPEqZeqgLZz3C
IAP5OAIYShttNVMTuQ1nAyyLE8sd0CJjZsq05Jd2BHfAQApAcuUCN5ocTQgsrOhR
U865NyLvpdim8YZBuYfTEl+16WdOEKHDw50GBVT2715QhuWpsjpl4+6BdXxCFqVZ
SZgwgdU+mUGqVl4nNWR7tYQ6FRKLdJUAw2/XbkdyH3uEjPiN0tm7zccCN6muyW5H
ykSccBG60o8KIp1FUqd9g6fbO2qlptrrz0P+0HeIKc2oToN6fJ/pojzm2HAVtGi9
Ww3KBQ97SXSYPGyvVT90YUtOJQJXApk+D1KBjuUX2f+TCioSKimPKLoR7nxgNCC/
bbKa1ZP6AyjvsQIsPx/7+aXWdaV+PJjQEDl+pxw46eTKM+odWWNS/pb+172/dSGt
lch4XX6TjkCnlF9ZNeMgxKikoi9gs1NcYNX4WsnGK5uViOMHW+qxplWoo7MspOUw
e3mbyeR4ADVoC4OPKl1pc3tfHJ7pEZKNvTjIdsYXBKndtr9FjaNOOyeSvM3F81gJ
dMUg0FoqmNQooZU96V9irKdZIpcgnjMAPROybbuuNp47zWNNYUHYJupCsr7F824X
MMuS7PsBTDwdBE6hZh7sHFD6xExSlNMpcChdLumKi9C8vjCYXenTFYp9iVWRwX8u
nZ5kYz8mwwrFXIv7jltGMnur9x2eS/HMlvdlPUw7XRAcoUg1COAphrX+UZl+HqAB
7GbyJXShTGWXswKwY0AdRH78VpyMWIMKV13JsH+G+BpuNIvGqRdDkjRm9BTFur/d
ZHeyBW3Dd1eWTcY9jcQfBnXIiIVE8/Z2QH07aDQ2Olq3dksjdUrq9gzwi/ZA7vVO
HbjRxDp3ri+EWBWbjue1Xepj3Y9BPRn03yuWFDcy5nrPzN54vbFh+wP4RjLFjxEv
xBs0lQf/xDQOL0rtmgvmop4Bb9i0JN+J69kXp1cwLdQ/T6XE+lDspvMlFvAW7r/Z
rOZz8GGWPP8vCtF+e7f4+KeK3jKfONOyEltyjZafcp3vBmzsa55M+YBWOwdqq2d+
cg7f+XMuhe2PbV6Hw1mMK6VKKI9taiERhbTlyHCIT0pWnsAFiAjB/z6BkvQ2lhSi
w8zq43vlZV013DKDBmZwzQAIvzFWIHaE5vDZkmoRz3iD+2AI6ENhRsI2hVyJ5KKA
vfIkAgf2sS6GzWA8q5V0FGqBzAgonRwfnlIimZ/OCJSitQMSP2XeFo6h6seSLKht
EIL0r33+eCMZzzkq5bK+jQzkRP76ISQHUZV7RRvqONIuimiY6BdOQa2yXWOHtGRm
VnxIEZOTPu2GPsI0zh7YHZlIXTWC7XqyMXniLNFjDm0fPz3Xt/lvhJFzdnvXHGFi
niToUilAoeP4Ev/gLBqsFQ1w/pD/1FMxX59sS3GnGzhMqxkxA1zbTboPg/sjR7k+
sqCKaePapU1jKHXofJcAzTpjbiqC4teleJPslTixGKJ+EF+3FPHGszWmNtXusERs
NDHxNaclUXJQxjQhPig9GDJFZBPWIa8iocGbXs0DlfbcHMm/nEwBxnWwgABrRXSx
mr4LtcPgIYLBnIVjIrIugL4NVR5YyDHSsEDqTrR375kGk6UiFkNO/pAogylndrvL
1gsQsV01Fy9xct6Whzy72zZ9667XRsK6L1HGCNMsQ0hZs8jQmhO4xBFTvuAX7AVK
ZtPNYj9ltsm2C4VDhlYGbsmbSAu2sZ1ktguDEm5Wu0TQhXdoBy3jQE41HTZrcQhK
k+nVLEy/Nvicw48efGZeKOxQ79jrL2qrzShEFagH+pzmzuiPyxgu2fXPewi4HqBF
5kMlquqdyfrf1IPyvcywvtQGBEeI57R+Hgqfg6PqiXfkvjiUZCKJ8f+bjqfDwFoe
uCmRoNIUPP3WZIJam+pwhGwuZDOcFxX9+nUaWdqZwUinEaQ4bO/fNbzW3xkJAz2+
sfw6rWR8eHx4staNma86uThC/hH1qT25GUKFCKlHasiKroVxeiyGyy4Xp3tFDRmE
C+2/+bTH4mc3+rZ0Le9BmSlmhAV3kCisnV3iXOlzbCAWFhMG9nrj7X37XDdwphIe
JmIO7HuYKGd1ZPzU38SOjOROrQd089kcNYmjxgWn31YCITOReBmzenSsnIVKni5Y
K1QkavutUkLNQ719ZZn2pEZA6dOWlDbIjVqFU4KX2FlOoeCRFgt0Gbw0L7WhK4xO
Z8gAk8pc8alW9GEmuCUOuE1dmUggJQc7yrgJb+4wLLqsX/TyYzBruFGwPuKNFKtV
isZub+9VopQ3sLMGF2/cZVpocKEhHjM9Uk61jxgutvyFsrofw9D9d4Cmu/6ZZOk4
vgP37oKrTblVfHm7qDvL2N7zfPaT4WThDYk+hWQFtX/O6ZKsi5xpA/R/M4a/ObOM
7ACzXn/xT+DpgJJPXKA+h6DcQppEeI0nb18klyE3nrvlro67ObHUb0/C2122Ck0k
5U4DkMbtKCU0oSS8wLhGLx6Z3EBGz8pK+Xy08P/ZSkWq1b4QyYBWgLLc5tk1K+gv
NKUlyzXZiUk+bDAk1cKAy2KhinVMXSg0dJrJkpj3cQm4X0Ad/sKRUyZsIrAImLlC
rBOlaqEH2YJZG2TEbsIE30oL8RtviqsuoIRWmkzQbi477mMzJm5Q+gWfPLogy0E1
ZOThyJJiqhGRHg3h6zqv6kKhZoYGFLmQtPwDyb0CjVwPncXZnraPJH/cZIpK+HtF
Bm7LI5d+Tw1XTwdqX/LKigYCJQXhiVvu4Die70CntYxVVvdnwpL9vWS3nKez41NU
yimlUHLfjyEDpsfaK/QiBBHFZAN6b+fDY9GHHdEpMVy2W23Flid965aP8zyU6BFf
q/C1S8bxpMMYVqerYBNKXLaB0xfKouuQK6kFqggaBdFh2CWwVLdPRq/oxMIauSDk
ABexlDXcilhKN/WrAbA2Rtdvf3XJDbpElTxDjYsu2ITmGdP6CRJjtbmJDzXta+qX
a5VurRooeAb8vx2PL7u1KGU/TDLgxh6X50OE9Lkv72u9elCfGHWEzj8BfmkDtug4
usSoQWGvwKCmLp9t+yPV34YM3xCEmgQTi0A5pw8/GLkTlkoP6h2t1nVDR2JFjXDa
30ZTIKxLlUpazFcRXqeeE/hM8iKpL9oZ0Gm/NbYeL1EUAIw6sSz0qtOHCSpDmdGA
7hTySSwNgr1tLnvSb9NAfYA1Tni1FUkUYX11flxyzT/gpZYnTOaf0b29uup6qiNK
uZQal9j3KqqNWpZL/difFUNLcKxdPqs6IN2Vih0zh/LRsxcjSRu2Oc0OENIwguSd
nt0pgIOCyQuTxSnU7KOuCc0hKsGbqAZPNsupbDhHL1TZK5u6xwfhu581BxbNHde7
70aQSZ2BlpIqqYT3pDU4xB6jotOGbaky68+Xoh/SqpZLGEYYaXK37DPs4KZtUS7n
Zgucpl8OBWtDy4I2xVPW+ZpoLahyZfhZLxPnW8u0duHuGeSabMhMWdaa0CYkoYYc
tyZR0fcneqsevPJxhW5KJhzqQhhIShu8h6n0YBgpTkgRhQs5t6H6wux2KHsS7F0V
h+hpCyH5XqWoEgVNXIAVjeV/1T5MFA1xl2dfWTax7bt07ns57+QpHo7qjCkjN5eZ
x3BY/TnQ/3t8+2RSLfXEQfCL192X3x5oZ+KBvZ+CZCUO3hrGtlazWjqeJ/lRlEuE
4cXYuYgNc6kpK5UUVf5D1wBDcopHU6UcXcy0rkWzVphUW5o8bGLNy+qutySIHAYc
12xc9ZgMbd4YjcEATt2dQgzB56q+jRiSwawTbWLr0L2QxXvS4ktxS3/USz1jUfVG
tqc89fcAVh3uOEfzeVV5pA+voMMDwCrTmSs/x9cnaDxGAhh3IzrhwH+nQJFGkq87
t8L8aQoTbfWSKzcHP4WdXRgQRlglfhFdMmev7clenvq82I8mkcjcbDaJXbiKje6k
xJ4pNOqq6kJ+yxUxvQbp8pukvErYAOEnUd9YuAJDJ+czwAw1SgmsD3hUqUbn6UV2
oae00sSz0w4HLw4kJwL2pMdtU0A6hxmpgEmHo6hMnFoElwthzTVw2DxZu0463i3V
LGCI1aWLq1ztjkVx5KCyTJS53PYddEJwqGXjVsoD22bRiSk6sSDn5mOL2woMbwh8
D2cBCNwBJ0/6Elj51sfb6D+4fuuVqI6ue031rn+ApggoCJhxLwVMaQQPaByHB++Q
zAb8Lso6sjXVVM64crWIysOXqXVPefpkKo0WO4fW1Vu9FV/p6l3wj7Tz//uVngM6
iJMT9kGdhZKHTysXl8SNQLAn5WS+ZCqZfGZTwLMb9LZXOh02yYauOISwbL3GXPsT
nFym+bexh5K2gBccDVztgBwO3gBcjjlbz+IbUpOMtY8PTUA5klHfKub+nJTQVGKI
JL+0NsbezHF03UmQ6ykOupqBXfJDQ+gOa3+Acl3EXJrfzfzucuoH2tY1DW4wcJ11
pBozEmdEQq9bPP5yRxFW4bwEJMgmMJpsfGlSIlX+C9R51BTH2gF1tb0K9GjTcWrN
NDLTxaAf1fdJ4tTwCfZX2SPQOZCYFXbvlJ351pY+nqCRgDLtOwVLnyt2JolppYOZ
is+ITjt6GoV6/trHXkKQqMOEIYnSxAJgKN5Qoqf7WIWuNz6kuU8WJ62l6dGeLZfx
7jXVl1AKQNKpWzqbDlC5UXotL9DHkV5iJFuwcBByotNbdGgM91AvoLNc1a9WJSvb
sE24bcnRLozIHij58ROZgINhRavSiru2KcUWPVSLm8lx8ebx40bSeGXQKsA4DdVM
VIRfxofbynFneRTMHS3ifEg/VQXIfmr0xcb/AIV++KrPmrE5zdm9vO5uR837iaAf
6PiwxfRS1/T3b9ws81BX+HedbNw85zoZZGR5Ak30N3xz7aDctJrxsljXA7bNw7aZ
GiDUpsIqtr4r2o/jPL/jXMIXiiSXe9/XWaqjy/fcE0Ro3NevH10Yi2qtEHOQ4o+c
/OI0Bz5qOaRfYj5pEsWy88/Gqy2J66MTmyDUAY5xXXUOI1XCfzpHR+0ZHjl10pjU
tOLkGCfRUiybHw6kWv1xuuDjOtOYepKrRSumL8AJ7vZCLFm2wdajoQN9L1oy9EWb
bFtfULtbGTEJ4IPd2mjvtCLei529n8qNKsUoSh5dMk5HetyjljjfHbCO5M88sue1
ymxd3WrhDBs3YXZjiTXHjioPaK0plCcG0zynuOTgPfDDf9ks6fuiQS4eWAS8mBBx
zX4cww72N62YfXaI6EBU2NZ+6AbS5VaD057DaonVkKA+QDM4M75vCZcCnJIEq/ts
nQNhjBYXy+hknQUKLJ9ylZ31UHXtFE0qrxmOzpQYpxAo/Hi0fjgBoAQiPae7aman
mfejBaTXGLh20aiuj66ajSNnMVtwuScke2y+mczxzrv2R8UhYHFLYCpT3lHi0+w8
bfvO/RSdxo+Dry1H+i4xPqF91LvuNrAHIQIF1JJtuoz7sp3cUoVL5Y33JfG7kzlB
w1Ee268uLAIyQW52Sp3l+Do4kpXK9x64q3vrN1QfF9YeugzuX2tGvMQa05y982aD
hEq2/KlaxDZt7st0jhbLukn6vyzmPfEikB/60zbUa8PMwXHvP3z0tFMOWEWKMFd9
spKlb7pThAIVepV7dqzmWtXDMCk42wsoukv+NHzAjSj27R3DfuVRHrv2a1V9Wa9S
NQiFStrIs++EzDGqJdYaYzxlWRJj6UADZ7uXb8MYqvHCn2+Ru5585nT4fVqKan+R
7fQj5u69XivBpc3X67qwUTXQuPheBPtGwi41v3Z2CVdETh/vLyw+5VbwXz0MSR8A
+ORsKww/nLL1zgXi0lk1Yx5x+2665pXyD6dYh6urY3xFXv8MS6UZaCGzGhS+WdrP
MXhqIKmpG74YlSWP1a20oM0RsE22oBq9FOpotDkOhsXVqMSXC76Ab03he0b16R1i
CMc1PzfWKuv1nnPvb+0bPPeQQU/4u6ek2piz1aieEGgiUj0zwBzUsoYgV5Z0isyu
/GBvtIgMORATBqsJDVKQukrWyp83IDeIbwF30enzLV6/wrjsObCbKAtO+7xDYcZj
N/Dlg9GbdnIENqaOW3hRmKuOoUIiMoGsI8s59HPKq6MBzfFW9a+JUvcOt3smOUQj
CUI86sg0qt9799YjDejhbteES5CbkZIt82pn37d8QNnJTIupFPQ2uEVypvgVLE8q
R9GpWE4gZp+PjL3BBLkZF3Vkxm+mbFvS9HdKW32OGJA6yCkvFweAI/5Z0KR1ZHnk
vEjfLaYQsJNksIlV31ue0RrbURpDWAFX8c93ljJ4ckCP+y5g9tmdDRwcM9egtTli
zj+lA0Hwkxki8fL5/lb2YXNlnu895/qAtWfZTd9wtCQ3jgWpVHkQI5sRTI6kcNfO
m5jX1/xYExGeAEUawzRs/tK6sJTw+6G9k6NRSwOUBqZc595G7ue6kilOzjNScQMT
6AlGWSF42+WdwNaJpPeRalxauVq5+zTk6TiF4xB1rUXbmXLFhnIrBDCMbcTjTAVe
9HljPixHpuioai7+HVMdV7Wnpm6XnLV5DeUQRwUMkE164/Uo90pOrYni/7VyjEoe
XBN2kkmSVHGzA5kAPrdp7Gyz1dkj6zFOmy8P3c4C8soreqqKRydrV4jfFZSr/L4r
CNqDbk+Mkz9BM7cY6rILEHO/+jOir2Zn2Tv0bdGfFtrrrF8j4QRVtq29uIKnCnmX
eM53jBZ8L3AoUEcEVHqMonfPr+PRKhGjZZFjivxs1MFbd6M0T775iIVMHo59aHd2
mEahpCqPlMMu9M+3lwndl4uLsuf7UgnJXpH9x0ZSOXsqi/TJcy9uRBx+U1788F1Q
+AIwz9JNSQDYgu7mLhhJNPiwnXrt0cFwulYBTyyY1O238/688g+wNZxD36GD3G08
W6FdC+Ql38czIh80+hzOjM/3r7qXVz9CXfWOAfPcUilBtlFEcY8DlvAStNxVQz1q
KRHRpQux9RIC8EI3IDrO3d1OVbmPLdAOW3rqueC56f2XGNwr+Xn1Y8RbhJGPK8hY
lCc7WnW4izYtWCVsl8hxOvMq9Ma1efco0sFF1Djhl8fe/l9UL4h890l/7WniU7z0
EDv+8KUm7mme6fDhhKN6s+opT6MIZnhCoA9SUvkttzh9Aa5VZ3zJSMhP12losUuy
27TCC5TFd+ivDyknQQzcNfBOnqyoBLwCgBszdR04DMDzVLCZQ8N+6z2I9hsLcOAY
ih5NvFyFejDgopm3KdtRGMmpRsW9mm0L24Xvk/vmtfG5DmHr9G/Knwpk3vKCcqQp
3z8GwbfdYc9Ir5C60fSXDAlXQX2c9J+Kubtb7moYjd9lfjVknnI37Q0H67MaWl5w
jui3gYgW/fxYSOB6RchBXhBt4D7sYOJwRdfysuAaHTnVM4Da82aqkvuOsi7cD86c
/D8RDq3j2hPP4icoXsyqjHwNbCzxaFsn/Yj4TUzK+WwjEZHFa2JXn86j4s7Yk1mH
/CmiFq4EVrr5n8qwJODThrZdxUWJT2Z2/P6yKVUrXG8yxVSvvWlSAqmnVWJqYBOq
rtvrJWikqns1qJb2dBUqFVwHy0Qu8Sdma9k353YEg7th7PK84Kxk+UD6hIeJrYov
Op3sKSNkumNCRWB7U3PS9qxllkdGRleV4VugNSAa9jv7rXLlq2Vyo0x5G186Sd5o
CMOfAcbekCCz6nSvLF16RvPEyi6+CtHR74nMeWeWDdTfvXIxi1R9Sq5cJzKrJQ4W
qiM/dAcaQLhyeiaDuyw+Miq8zOjnXfLRhs+bNJ5h9c5piBYMVQfxLJi+59v17pH+
FCr0OkcJ0m5TCTFT+qo2Rf18dOdqz2jQTecTb3rivaoYJLXgpNOMaecWk5xZGzyg
LHnA5qtgOBceKjHbMGMlokyMpeMDS/503xF00TJqd2NPCW1RfRu44KSBstsrH4bZ
wbmfzco8Fv02ixjbl50KfrKodumwA+/LrLJ1rYPMT9Oc/yUE96DI9n9kxU4kJRF2
x9Hw4IGtJ2qOe3CSVAaqclZhi6SjCE4hwyWwESJJb+JZP7PkTFrPDYTcSRfGwoXL
UpxJc4sxFbMc5Tx3YX3AiKGdlU9T7Bq26KJOKgJoo9yuYpBc3SKimEnbUa8bDqGg
TrKx2xpWYlbtEVQMmDE+yOWFWvU2yixmM4NjVU8DLwEhR8FYq+PbjvRx+/oXu0al
9TSNieE3h6Xbb7Ju4lZM671AAyne0g5mAb5sZTicEdaiDhi3vaKWOuTz5mJMUUYu
7JkaGo+1G/ju8L9Vq2cC3TatjK09PF71h1FmAs/IUynLlOGQBSlrnbfP9QdN077s
fdnst5fylTlIKhOfOmmqVo5LaMsAGTmicNTOkur+tI/bdjyUHkg56QkkKWRC7jch
r0cmc1HtmlfuHEmKPVOOMwQU0f6GbUFmrIePxMTYSKqRBfUtr2Ec3ePweP+MfxdS
bRzrq7FUf1QDWagf3kUFz5v4h4zSWZUMBxxr15H7S9HjFtt/kzk/GiurGavvVLa0
xeQErTgmSyrXsI77HPLiFJVqnbwYlPsSsWfYl4EvEreqM8ZedbR8/80E914028jo
VXqA64yMeN2jk/kJImvtsNbk/1/5HwutxrRQZ+A0RqXMt7d6u0F53wLU8jmzyRwF
7jA4BNnPhCEVs01JLqUZ5nskiD/P0YUsuYTfyTd6mJDtF71W9ERYFyIFtrkZrXn8
Q2dIXAZDab/avzCmZalj/renijJnb70DH2/Rb3AMw+deaddTDNZe8xBpElrFITwd
466Jd5SatOk3VL27Kde7h7uJXJq+K/t2P7aruGkuQXdMkKS5W2Vwdv5RovpuZ9QJ
n3rqpOvCIRwpGw2u9r2mNRO3zny8Vlib8S9Sq5DAIIyAQfXkGpO7syIEEFuoTOPy
qw+ov6gy4zK103YLAai8L2SZAjz+3Ojz/CIIvq3N7di28gvW5lNZll2bqR6XTSzY
nKGdsPGG+H4yzqobTrcKRuERrBVPxeLpewA/sWkRzLLk+K1MnxwRonOh1EGxmLZT
63TJL+IGc4oDPRN8wz/pr+9qy32yBfEFhOK4jJUKoT73t/rMVUee/4/b67Be1YBU
n0fqz66JM6XteANMvTJB2lw++RCHaQg9EhumceB3lIQYH4wSpNSco1cDa10nx3oi
ILv8c3PHOxz+msMpO+Is7PuGRFfDuZWVjbCzGkw8V2PTce0W8wvFxMxhiiMBAak3
5vC3ZMzyOt3KdxlYKx5bK58V5A5iFytw/viBYT/wMt6vJoo+rUK1QP9YOFJF0wlt
EgUOH5+Io2ubKKCLuzaJjhy6ferhQwPURLNhS0xxkRWVRWdn3rncLM0MGWHkBZHs
7MhXGjAqZz1KfDsooL3CfHxu7KdpqlMvRNR6oIoKxyY83W4UNvoad2OpMQvXFg/t
GjMYa0unpMcD8agz1mCUG8zKnOelwZlfZk43qyi3Dl6SbSLGxnEdf6URmIrzoR67
iDmW9Qgvle9+RSCw2PFXBJcYgnd8uTvz/E7PDUje8ieyKSVOQKhFarYgJer/kYm1
qytetgHUXU8CMhRuCskEu91me84lPx9HTRqFoE3bAEqSxV3iNKV4w7wFms7c2bZh
4S5nKbWDUxGdgNhGE9OvGqZe12GlT8e9jcVA/ml2b/aL6+5Ogh0M7YYIYEozPVdJ
X7lR0Cf6dtv60/f9+DXc5UdGq/W7RcLtnPj1CZ4DnHWDeWHxeJe8ud3oGJErwG9P
wTVVsh4QdocTZnuSLVQzX26e8/QccSWcz1dEWmAy5lat9txYhnPEAa1NLvEVSExZ
7dMneeQdLsFVftxiDMIaTKzlt6YM10VdPVwKOQHYiwt2g19D1tmae7jipkxta1s8
03qM4IFZT/ClTh0j9LPd1bVzSqyD11J0NeVmMYOxTomw++Q8cXY7uKH8VpWiHSbG
cMdz/gE98VxG6PAHuhUBor/0xdRxFLzrxyStQeuOAhu3QMbstPoteVmWkzL7WAFm
8AJdpdTYgIlut2FGpjlVw9xhxYDBZP0Cd1l2AQfhxbEjSvAzCBOlhXZ1idhfXKMA
D1KOQYu/iat0FUD07XucQ1exTVlG5LDlXLcFf/S3hlfqJ/AEpvLKRwRMgmWiE29Q
5FfYoFOvn60JtUcdHPa6ARCLw37S8T49+lNGJhB6dX18KsoGYebKqS/6jo7y6Fdd
7Ig8tJDqx9/YQaK2Fb2oqkCYjGcbqMqaaCBoTQb9ijEyhzE3qbDJe9RcEpfaoVZd
sItebWqEkBF/kVlXnYfXWVKm3NDYqI5VbooaLY9o2IrCanXKH286u19Jrb3SajLd
XkozqnuAaW8QCWeiy9y2XPegOx0rkn/2mGK00VcvDrGq+o5I6qMhKQpGISQa5nrg
heLLkJbJFID1KWFfG0gulFlibvmAOtiLAVD66+4pKBG7yy2UhIr0EBBoIQGGtaKE
Va/i7I5L5QxWR6zf/igOMJiOKiF4QngFKIjwUJWt4NQmQ8h19NnqU+58t6p+lONh
pJUU9F0zUrlG8innyvDyKjb/uH2f+Hxj+n+Vcs3K2bBLYRkpuMNMTADal5YO1BXc
OzB+6qpkugIPEJREXA/FhHwTUvMgUqtObLMacI5BmFypwASwDMB9zU+8ES2P5YLN
Wr4W6edNB9IS23vZzgoWt/dQV7fe1g7ZmyV5w6WgeVhKbA6Mt6o0HOUKcht4kKDD
tj4vVgPQMcC7Dp5wPEN0aHJenEplPcIL5mHth0AW8vsg/eObP3RmF60qEUf0T3qv
gE4KMtGeiZePBOq/2X7HaedX7w8pwQiN3T4hWmTZGVcvCdO2G29lwFgxA8a2JzEw
AieIO2BUJDnGzM8wWdYZEWeo4/a/nxPFXf8W7tk0aSyd1uVRdRY/JegyujGTRnBG
+7m1F9te7wxoj9GdvvNrqweT45/59XKJ0TyfFM3UBdyDWiuUznwdMLefPHdbvHkN
DA9EmI/wbKpdSzEMN1yd5KorgYwxPLkGHNy01aSjns4lIcoaTtZ7SnjbLn3ErbIh
7HB1lFmGJGjzlqYlwjhJM/Gn//FZcx3mCWi3raTWypJSef/e8UuSYDK+q7wWRYzg
UJO9fX9gj15o0+QPAa9JUwQ82NJlD8NUnbXuA4NOBmomwjVRgHGTPH09TpFTt+ah
bsIzvOpY9Rk2Z7U+wCmwao6zpwYsTQ4SPH0PVJy1F+t53QXXvqnsE6nFTdUJSQOx
6Q+PBtrPjasIYmP3HkpByzixKxqInzOmqRXWT/QPAtDlmggu31AYNd9cFcW9qXyo
PlpolWwLF7YTiykeHhlKLH2SfQpXtr1LgY5jqIyDDQ7gV5BIGjKX14xFeQlhOIq8
4nazFX5D5cFRr6ZOZ/V3kQfRYghxW8A3fMN/JmhlJsDHjfYycyeN/xH7rC4Q7cEc
y8849iPP2PUeun4JFqatyg+URsaQTLowdKGMnsgaJdw+upxIZ2MhrQBEMgFd6P9N
kXH8YWQZeSTFPqH6QTp6o1lpcrDjWxgSc2yEvNXD3JemK85uyhJn75JKoVJYrped
nE6HjNE8+TBqtV3Xqcrw2GGrV/qpe4W8V8/l8cFIw8bLbUiXpQtNYakxk7KllnZl
OyxQIcwfCRpjp3hIDIqOh+udyTDuyq09ZotODLIZbT9cnY4M1JQkj38JkcT5+3va
AZWoS7lvUUYdPbZSMKQLIeqa42WIiWmSJT9Z2NckIxr0d3NWRkQWWDyczlONpjh2
xJ74o57lEFl2IFDq27ESpTtOyFYqCrDg0ucghNp+i1jCimPHd1hzz4aOhCte8J/t
QGx/R6m9ZGV6aUmFDn1N15kogi6vby/a//dsZ0obF5HMN8q4zzK79fpqtRD38Ex1
pSTwYsjbnp7pAVpRsuW4mZdPXaI6J9ER5T2Eu03VaZ1bF8n/5urGoKTjHnpkhtk7
F7nZ+X4ZynaGGWJBWBhSttFeP/o5x6ZSVEtKpXMVCK2YLCf38K+Z6D/5Bq9Co0vk
NCLAIdr9gpLKfLxBNabAqNa4pNSuIg37KOVjI5M0nIsnyRgJSPejj9Pjp+ltK2Fj
hIq6fLrJoADzEi4oYqJUuqbqXU7lb+TgxfLwPzZSNL6gs02BXTMbChPBx32YBOqp
LxsJ5CYbQITt3nQCGkg8Um6TugkNGarmJr/F4jyMT9nn5sV7AdDW1QHoTgW9TVpY
k9jnKuUnVsTQXODKGK3uldZ5R+Wl0hgBN2ReC9C4dRFaaezl8yQ3JPh+0jlvGePd
AwnUe8WH3jzVM+snrBCj1uWfnulDGUyZepsBQ+/61qQxseXUaAIXIu5JU5tE8RbN
PBQ+Fzimr/3V/mYEcCztqrjeg0jQPGMUViP0iXT65g9odch8WwLHHP9u+COq1fsF
Q3YnMhJlBfoF76nAJ42wicBMCxTX50udQiMCrGPtbYw9bXR+4FeoBKvp3ZUIMkW6
Et1q1nGW6hO+5fvYTdLau7o2m9v/PmCs1rOK7st8XxUcScfE3hdm85QvAjd3iHI9
ezLuOHtPnOtRKjk3AVaJH1qvEwsOwUzfo5auFiF/89S3/laWmee1jGkusyRZd2lV
gtcC6PQo3Fe3+vE1v6GI45Wm9XO8ITEYqaGwdrYrKGSCxJacqQkkZ6X9CV3scpY4
1a5nwxTNIC72th1h5j7eGdFUCoSC6WlsdjBT3CFZnGoYHvjpqRW8jxjzqWfR7sSY
ybGXntvW6qfUlN3yeKow8G05lIHJ15YIFYeCkOH019TkS9Xq5Z0GEsjT3XryEr2v
Y53w41jb37KgFP7SprTh8gskelrtdfUx5ueZsc0V7007f8AFG5MTMGjgi11KxINm
sbdaGNqr7pvJwMegT7zY89WiCfGgO/BHMjiSUsyNe4jmVxV+yW86Iy88YhVtVFaD
3NkscBvPBgCeW6xswPd3ToOAj9mwRHnMWpoZOBbwjZpaJadOeUyldTwuvI3s0KCQ
adez0Zuev6xY4gjiPdgtOUJkGTzoO/tt0h2uSJvD92sPVDbqeJi8GHZ48UrelZuV
ATOMDRZNs30oCJMDLqznzylNx40nKAPq6TPTJsPMJl1ciB9Jhay96V8rAwdiKqnp
zSo4hbdAWZ/K1bgFkknukVIWaTjL81uazfBGIZe/pSy0IrpBqC6QNncAkr0K1XGa
qmBTPOobUXOTAKm+FCGjnJq/iycvKiaeG0xzyu7K8rIUC30urdCSZtFdH62y05dN
K0BQahlQH1NvdOvNnU3BsHVoi2uQGrcp1rEbBupKBIMBTnG9ks1XJEMLtAL14h7r
u+Q6ZP7cNkHtPBPK6Qs2WU2pTXSk2miGWcGjOtfoMdWJj/10pGrr5CDcYreJw0ku
gBkP2I8SHptaNure3DR4y7M/tQTYcj6CwnAtCluplmu5xr9Xbk+obRyxccQLwTSK
U8HwmshXycnMBbigezQNGtfODY5mUUD80eWL4cDDGMXET7JRoNm80GBnw1CO6a3c
LaXzfKC2LyBSKJY+agi7c47JyySOXbRLEixtEPqZ+YdRkpVmBJMBAJHfqrc1o/ke
2GcX3ioge7MJziTqxRUHbdlRcYQvKMgNj5HaDggqCLbDPFyWDmBZDzoWQ8+rgrs6
iydOGhqC/CoVqGeGQyV/M+IBYPQSzZdNXhJhuPtWWUNHb3Cu19E2pzG+pBOcO0nB
TTOAn5gIzqSRg7ZCy9SdZQ2jQ7Cnw0zqBq5NGmIOIF/h+1smRMViOKTe2YpzXqA0
BRc/XFeweIODwE9URDi+ZwvVHPhx1Yd7zG0uyAOGiaNKkW9d6OWhfCXNNi45Tcsu
/9gSEszoZTO1Rn5ItKXcPmWN9HL82jPjaPDymkZzqnRGGwpBDhgRI6fesA0XFIg6
VgBTaA40Q53SvaHOD3PsWkq1PmdgOB5SLwr37+6qE0by80JEAw7bPAX5WQcpo0mo
QUtifRr1PMVEmUnzVmHyfZfHxuo1PfcOTsZ7zsn2DAnEhLC0SSdCySvFUdFluYRR
QY3Cl3++uQv+ygrTU4FrlAH9aDBUjC1+FvINgpdpjvEiPj0LCg4KV/wKJBZuNbEt
PDJLFl3nuPJyJ0XNfRVQeT0vu3oaXtVLv4HByR6q5yISnUb/GJnbnsnNAmiPOdBD
9hrwJTDCOKrvNc6+upKqWmjnXCg4GJG7QyFk1uI+a+XwMHEgWpn1m3IyVh/fg07O
o2J9DSdtuhv71GK7JJ1qjDBxjtScYcSWzagQEq9eMFO5Y6Vsm0d9ZXvk/bd9z8Nb
OV1UFw8PqPtrZBOf41pqHHETWZnK+duQNOKoIlenxdbfGER7Kw+X3JcjNdYNSw/M
iePJZmLn0C2eSJ/HlgSqJp4BEnepI67s40cLf+MAu1ewLm/XbgUQvquZXTKJ21h6
VABbUKURRhLEnBUVdYGrKDLp/0B9sPdWrpO+8rz9R2nkqihJVKuVtFL/mwiBsrRe
fiGALlkoNAMcqHglC6FwCpDy8VgUUEhfxktECSJFIIsnsa+RGZR0aeGw1LzqUYK4
WTAhZA4KiZ2ZvgBtDrdU29rSmm6ZOpKILT2NzpkfZVLJKIzNLCJRObxnymon0fKK
bi7s/vCl6MSDHGibLMjxziJ5rXsXzSOoC2OUpZwNUlfKkiJn9S2lFtw+iR7nDP3V
vQZmhOknZU/6+ai8oSHKspgLEXjat3jJ1BgeznV4knHvanarMCTGdAU3C/dUjv4Q
w5XDtqCzB1jESpM63A45/iFYIcXp5HaXvqEQBIXUiDSmdSTNAo1UgqhBS7e+gUER
Tu2ltOBfSn8asP0t3qco1nyqhdKWmOtKeWD1h2PHqigeor2ldJVpMH9O70bXf4jQ
45UvUuGqJxAcOy0jgLx/u2/ZNnIBWVtha5FMpzSPA99dOyePQTeDzSYHwivMEnOF
CIyJ49xVuHERdvcvB8ndJx+o73eORlChWV5QmzJFqkouRaerxTlzpDxyydkC5DWU
e4IoPr6nN5dVZcNMC4Rsryer3wfi4WaleUFhUoRtJLzaBEb+N/UiR8T2vdKbVoZL
3Oazi8qnDIGNj/mTltvSCR0a0EICIEjw2FAHH/nPHIUrwi0vqVMU2OWNfsuP8NWW
c9v7lpwlZA/O8UXevvMNqZd8+9mjTXh4UROwXMaysuZYVi2H5uNYPuYwDJ43JOGe
wAWx2AgSVrURvtc2So8wsAe4yAQaQ1cK73bZgrv4dfQx2HaCS3+NO+ktMRKB7OBX
wxzByHijY5MstpU4M15HKI1fyPaChualQ0+spEgveVTUWiZ2DFQe27+Zpg6xjkqh
0Sz4oGhSRuq8WS7o2EaxvzYMwcLVRU+gc7ngQEdepO6DnNNFQTFg9gCMsPtb8sDR
F3HA9pEXbz/F17hUzTFJDAl4slNNrIEIqMvhypNMGjXEgaZtF4KlN8nMAPyR58+b
DkxEcZ51M0ViiZn0R3Z3geZjy1cFvqcMGqGM3crP3RKe5ymQpo1TCaNHPk2YslVi
lxi7ilZKBii1XAEubZVGN4sppe1xYjn4C1AjQZ9Bjz9odkCK3F0qr3HSdZL5WIHz
2dgjYks1MOcbDxG/LmIfDeQoNYfFdEVuo22txlE6BX5ehgCHJZMIS/UDbSF7S1SJ
c9PFbbBnWMP/Dg+wIyEgOn3KyOPTPuLH2seHlDDd7wskGEMy8o4GYch3Mg1t62wC
BNwx4tARm+kNAN4RShieFbyLgvM7sYWQeuyQBOG9S41YDlO9Uq6z2Z9BahLwOI4X
D/PKwCWVANs7o+ooSM3UoT++DK0judx0ZF3YPgCwPqw/QsW6D+1Gf0vnFmRgyaM4
SrXb9M8EqWwBCAvTGGuI7G6Gnt3Sr8rB3yrAJ3yoS3a4N8wjOrENJ8JpHl9Zj99k
Rll/jd9i++MwL+UAmBDJfV35O4gnH626thxzTELwnbmBUnyFTmx45Ffr8RWu97bq
t8Zt93xSwPqHsfb5PAQ55kJGcpkVxxbaIqzBkHA637k2fbbTxrs6dxDzlH7X5bC5
6BSbwMlAR/dQJ2PcN9VRd9C7lWKY+85zjgrBSlXqxQYWBmwDR5ew4tKBtfZUQZMH
uq3T34Xxfp28CbJOqHUY222FX7YY2JX9aR/K5dueYW0bRiy10+J+BQVYx2JHSvGo
Ua+ukSmpEsFY0Bzsgjs9z0OJcFfqUFaeDS6wie8kOsecaUsHP8DxFZs3UhjnSKno
2TN9PdEjByWIyA1yNo+EAIsd/8B4qI6dKaGAP8cfHNPmKqzSQf5pPcnnYL8VqVK6
4strxQTG2P/jy747qMH/pPYWP6E/Ehf4l7dctLNglpCFjdEqbquJ29UEDxgWeX2O
HM0WtLDwy/5JiKC0PJIVGVBXD8IsOq1gn667QSYHfiU1APMwno1uF5PyxhbtnxSq
dQGmZs6i3kQkYB6EF5RzF1GkqKTtu1Awf7At4AMtFI84jsM66C1hnYWFZwkNf6Uy
NINtNzg/Ocn3fOSpWMf1MvxuWFFZZbVMtUgSBFrC13TaynBYYQnkCL7UBe6RE9rh
ylmbyjmYXjrSn/wT7DbFsooZGBY++EV9kc7Yijxnu+KRNcLn8tVRh1+kyvCnlnEF
xCwAyrl1oBK4xeYXwFO4LiigdYhJHFdQ6+GaG1+HL13GVpr3DwiqESzZTWs+JXTo
LSJicySEDpdtX1OFT/mWzNG3rDrdcgU3BeCKxFjmMkZDgyzeBkRq4vfwCNMB/C3F
Gakk0YAUxd5hoMbXdeIXf7qnPDJWyUQNroQp5RiulNLeRFQ5hZSJkpgRoI1oqPuZ
Wd/3tValvv5t63VNpTToqiWaPTR33Hza4MTpjeA52CtaiISTQyNQkitL84+zCHhD
glqF2R1PXtITnphKoo8CFfw7EEWzVv0UeyvIW5dFlLqRWaMpM9MyLtM9CFTjZtr5
xlfPmQL98gHZu3s1W2lo/7OJfkzKKYSTzfBkYnK3t1GWVmzakhju5XslvrBNGrD7
IXqKlhjvWXf339uhO3M+PpxW2B4sjMn6dAB0jO8nVRycdp0007DvyNpZJ51g7XBP
mUgeu5i7nAyUiUAwUsqWYQaEAgXMRYSAKpCmewMTgH86qqCcJieH9cBvz+Oa4aMv
GASrzNsWw+RNAcU02LtKyofVAk8zVkIiPYKSw9R9lgf6quhxGULlLNKsLjd6hhQC
bMsZrqksYAkjQkY94mih8t+9yzSFhnh7BTMFp6QRqJVo4+CHHSTkCuxIZGV2FyoA
8G3M8T/p1geNhJYbP1wwFj211ddWbFzQbOKcwtrC4Msrz5Nb5PdQF3gHNtN5RnqD
x03NXdhYjsiHoe5b+ND5Q3WItlVls1qa0j6gaHPTIX7cJkVgUpxsu1ywDl27yBJb
QeSdrp6YiYcqwpAafeGMfKE6vSQ8WnEmZ+fmLPk3G7pWYJc/RXyZ2JcuvpmGLoP6
suxUc6PCNAY49zeVFbEPZQ37QbTuxXt1YIeOREgGDRHuK+85sfUzDeUWMzR5H7eR
7ePb1aT5yZyCg5U42fBWCym+QmdCl6RPlb8aHQcNYs0/x3HVeeCY3NiSr9JHko4H
8QQ5JFBaoO2Q+BnWomHGBLRhlmIdfuBfpfb1k9hFnmpnudPFR0S/Frtuj4HTZy1s
lMLtGomp0E+jOuxDCq2ea9EVH04nfl8dhj7dSUwHvN7a3kSF8LQlH/yt/mzf00zG
3mAZRrC4rE0Ug/RkTihF1fyuRmxLUj1raivv0JE+WUMhQND0BONo1Kc1wCGiE9nb
sq8MtyFKnS0lnEYi2QH9VfaZId9mgV+Pqc7W8esS7QAo8ot4Ot285JqEIRj5kPp7
ZBIINZDeJnd+gXV3Ix8pJ7Ly+E+whljILbHjRRlnKOrgx2yKPBpOxT96fiM1lxBQ
rjK1EtGjm8zDJfCK56+geHyzP0AOoJRmt6hKzPMlBKNJkzJrFJCdeWQYgbPqEqqA
izJgdchI/fvMZmckNtPkDoQSr2rJ3QibDHiaeVLi74rMLXC8RGoVlPPTqMX1MEO7
9eAeQSdZ0lEHVLKP6cTH+T7PYsA4Cf65NKCBgqtlA9dl0hLOYCBou5YwGpgzl/nx
ExwTlcygQh8hLFzM1L8I5Mt1Im4a1vSTMXGfhZYvO6ZHv9SDPzkOpYp0882F9aA+
pU93GT2r7Sd+kEkinTAKMExqNhXM6KhadXWtOgKuMYXAijyKuPKdizYPUsNwdhr0
zcLgGI/m+V9Lq6YUhk0Eujfw3HMkrK6YqFsYMS136fJHaTLCe7+C6fLFveR6zkP/
Z2tZYv/x/1P6sv46fsz+cEue2sfRk6TbBvpC1jedecoEZDOPN0RifyzTIIDgsmBC
EBEDnpkMlWgT9dHVQH6DTJ5W9NEnwGEhw38DLbxTx41mwTWVsvZwhAhWlTcSKB7S
OeD6dHaqKqKWLBZCh6CsSZocAt3ZRoGkIqbuqW8gldYai7L/WVUxBR/mNeTAJSzd
Rg+cJVYHXrlHgNKyDMMHsfIQtLxC+V05BA23GXD51eT3UQMER/1kpxlz3vk+mn7h
Uh5eYctKGaLCeye6JdGWsiDaI66qEQf0cDAdD0H3lnD9YAswqAOed87nEEHS28xW
OpRjngXNr8coE8njvuNCrbnmPtboGEj2tmNLTA8CqOUQzmfXeOvrpMCWolmz79jc
p4/5l/+YgettsPaFGHMiYsa/+zHQSkUYKGmkGUk26qSmG6U3pTFVnNCWDDRI7BCX
OjXkeph55F73OKjVcAbslpbvT2bE9wbIjEW5x+LqWvXldjgRvt+mUbFgcak2F6QX
LpJ0UxVZtkU7QcqrektF2nb0yaT+xioq9a7iCYSNhIo4oLy6VunC6p/4nN5Ya4kr
ZLlqLUozc3sZeSkTlXCRQJ2sMvWrrtV3FEYmxhv2Z/+4aDZzbCVeqCD9tC4hrVFl
+BAzilbEHR7qCmYUM+huBQvcN6sqRFA53R56xinXL7o1hxMGKJ51EBMzozctfCwu
W711bCd+LSXbBHEyhdqOiW9mXFQmKzCTowACjzdYP8zvEs43HMHjxRHyKnhe3vDH
IupNtz1mcruBHNrZwHF1eW8pZgwjv4+7n5q7qfAPSQwFrKpM00Rtgtg53HEnWHSu
vYdimCU7iZo7CKIUpHkYbn7tOk0QN9qc2fwMQ4RkYl2yoPQ/Y4yV49JStjA2vAlt
xsmGGQStkJmTul5pGcftP7UcDx12TsXrNPZjFyPh2mPaMR2b3vAdReKcV8JM0UTE
LJmLSkZfqW6h8hPdBfeqzzXvyJ/XGywLCmSB6s+06De8rW9K8Hnh0PSqdnC7ZPIk
NPzrj5AcJphniZ7ix69QYEczrQpOf76fDgX/5nCqzD6rBJaAI1/5aw/cm7075TUE
7OdTDanby0EgvVM3OaOQQhLhNMu9brhiUw9lc5+zPJKN6XQOrVZS0kVunhsx0yjB
x/xuXf0Cy6WYds86bci+0rjhqTJAzkAUVU9xP6QqG6KU/JNa/brASJ211+9tWhOS
15Ia0/FL6r2i68oyfcp04U9Iaycau0ZToPnAZBAztqnBig4VRHgg/sJiNDMAsByg
71wMBFhywVBfhpYYPCuDNwgGZdZEnx4SstncOgTtVn8L7UES5k7U8LUh1DF2JVPq
ZXu5K381cPXsxTWrIWTtE1g9KU9ogYqZ3DBthphLu9qFjIeGK3Z0r7TCjNw+467w
ddP3Z6dvZKIGbUXBWJABb+X3YvwiNUMwLjGKxmltmfj+sjxvm/qw8FmL8Idnq5VG
s4hfTbZnVWnq4UYwl5lC+LPj4ilcrBApR4BStJ+tH26JdYug5aJDQHMcXvNxe4xf
uFWGR1qieT+tkPCVqrZy38DgNTR0uBg229DKNzRj/AAoU9QqkpviRWjH65H/Qkz2
L8LWM+4ViKDXWI3guHCYdu6BDcp647AdhojKT+ecHlBIT+RZjTwITtiOgIODhiJy
GGllfguRqd/g6LSc1m80rGQWzxIerxVa+OB+q85jb3D3fyWL1vj7rRXA2lzQcUSo
F1W4JvgeAExZh7Q+4cfaYrvr91E62497qZq49iD9weCwiZc8dMv9+K/NOZv5vCWo
rLdUAo7cHHJLLkKAsuyjU2NZP4e0lNjlGNkxjpT7AADhg4aXR2ld484PbpZzIxMo
5p8Mx9EdiGWYkTUpjg2+6EBVtiMH6lI3L18Jw8wf3BHNFbjsOWql7O+F53T8bmzt
cH4pZgAfYuisJCFZWaNKSQtnjSHc/ysUWmDS0SGSsbHKKUa2Nfns++SGj1bkY6Wl
RjYpQsgYkRD2xzgBqZMDwOFr1TteL/apCr/FTQKXh1UkJGrS3jemU8uRygIoYj0Y
iKGFXhw9QacXpUQ+JrtuHjNH/RZHndqkFomGZrUHRnkbZOPYrGpcJ1Quec7T/zAD
WDrSknfzQzFgf1cproDuiKax63/oqxDmboKq2T+z5C7uYKZCBmIypCTseF0/xn7/
Y5SWAx2H6NkNUd4Ohfi5aAVpn3579AuCWaEgUNcU/2UUYAGTrorlzOOWQ2LUDrgl
VCbZ7TntN41YFBr5RhmP0Qysj7rE2MgtFjPdLyV+DCwCPc1KX1C5JTUpL/2x8ryt
/zYUmXdWEMrhTB55KZ0wenPxPu9lS7e+zPQjDgxm+Wmj1+sJz9cCpisn0EzKnxoI
rTBVr9HbNM/EwM8Yipx2mWWuYDDrzRC46hAYoRwfjQQDEI4OKVT2XhCvu4zTPeDx
jRFCrcmp+zRFRgPrziZ9v34N7cAdq92O3SWvhprkOcoHM+fK3ehXxbONnjZBrjR1
fJs11791b/WFc/foo2VIx3mWRSCjOYWt8PXGe7yUwgZU6jNpSJueOkwnoqWW7TFj
7LyT/Y5W9kbMdJJRKgjbItWYqt3V/f5WsnHHC+psUwNZRE6+fYCv+kAeetOJ8hJq
W/R5MzeIQL2s+XO1EHe3V/86X2+le/ANgz/vfem1muQhCCtZXzYyI+v+Sbz+W6Ft
HCf2pS2PwcESjtXRuMOuiJjgeTf6nlr1gcXURpnpThzY93DKu+27CnLoN8NqUux8
GG4edyHmUbRwxi6/Pn6bW9RgmH+sfMPeGr8mbUn8yCQtSA7yr0Z6lYxxkDzrjjFo
8Yif/giKt49+8Xw6+mLs/iNjF26ooHay2V+wWCQWhqpSwLAAHHArZYTosyaRtme7
Vk5wEy+a1rWhemlvZMkark5A7eC2U4VzA+etDaE/Ue0CjHrBPv1f6yLZb9Vf5Z9v
TGluGhTg+Ya+/MRCmUmSVleQHKYgizId1P9DAMJDbJ1QAAAIzsmrjFBBLftatAcP
bMXNwRvu3BrkBQRrh7At1sAZuYg6j8AWEuKdEA0VOh9tmhrJtM2mZqTC/S7Wx3nY
/13fKSPRCVBtaiXV7BrB1tE4ncEsMB9cAxm+7CreVlNuJu4HipHUEWBqZkfx/0/K
9MTnKomknwGZYhMlfDg3sBoAQlncOWBHwSCYJtvUnb9OwYz6+lvIM0YjG9VZ0FXF
F98f+uh86Nfx/CBTqsCdvpKNcsXITUO8fkoothrUAn5PKSZNkmR/YqqMtfJNrpIP
mjeKOhSCoW63igPI99DA9uDYFLQin1AYJyd0eI12h8rDSHxzVYhlpKauqyNM2QV3
gUa9vyiiq/kqlpvCARt1sZJ67A227eBNs77hBVRlYYFysg5fDG9158R2jG0bAw06
8lR6IuhTuzkijQMCqmFrgOi5vTunDJgmsyyZSflDHeJd0IIdFLTH5obPDMo5ibxC
6f0OgwBiADuVv43JUVC1kEmfEz/iWuc88KAe7ux7T4ACo9gDCfHoRCnuiPAVKBxT
kK96fj5uQmdAJGcywmRxDPHxaZAc4j1LGG6yHFPERBVmRSmtJpvnwtrD/UEAadrK
XHy773rmRA1GFYQJ1Zu/V/3dxZeu8nyyLDp9Q+/zC/+Hjs4RdbpBGGkKmGDZ9gE5
SvSYjGHg/6uhBSCxlf5KtLpvL/jyGpf67DHNEx4JWk23cXatw2EUjFGYKE8MXCHi
F8Zt2zchit7hCqZT/MFcYq2lyIX3BnqhH6zT6a6lQF4t/mIaNY3ytaHojxye+TOr
lZs+bNZrGBPl/YE+DhV1Bal7NNqLLKRzU0pWZHErg0pNs+nPgIyT/KN1lrGklzGf
doq7lH8yyUjUQ1JG3i8Pd5zHk8WNozD4dpWVlMdr+n1U2ZYX/6bRodW6V7q0Tvsx
enm6GTNDR3+URnEpMrWKxOTqnRoj6BWp3PcM8DwgU4UAavKEmeYkSrMoJ+bP7lHu
1lIx1PC+m75gcQ5JtgLv8000t1GWwFzckXxF0avtMfTe5VuUEQ4i0yMNFfs9ugow
X3pEQwdqta7Wg3OKBXxVcsgwxvFEH47BpA86HHlvsGOxMMcPcTc3movKGNFN+vyu
xWx7jbSyZiE8VI/zVZF088JEvHcoWeKmEqxmOOV9NWhsuFTSWor59amlk+ofnnjK
R0oFJQtkZIzeZLot8cnPXhfeAhW2zvhng4d+18XK4XbA1kyfD0D9atnxZdV8jbYI
FkYtzTu8baBaoKiANLLJXueOhrHmDR0XTrO/2Ph/QF2h6b4py+pEsp/bvfQCr+Ps
DYFgqSOzpQQ2muFkRB/95WwBENJa9yj04dRE18tRnFO2mm1eKgzVra0//z4nBTpr
RTPIoLv46a/ljDYWyzMU3h/FwzNADZKCTl6XNdkB+GGQHWRSoAdhvbhg0/CSiMer
0P6j6OQ08hqdOpxm03RmTyHJcY90amG2n+FfgD5zy0ufBsAyI1NnbsTIRTxdiJZw
eqEG3hzgsZiVQcZB9OyEJQfQ3iPV4gRkBCre74XMuUf5sA4IucmpBsDJDpo8lJhy
/CHV4hxXYrvP0wRgcha99ga50BtXA7JN7msGYrmsQnL55MEuk2s5u5Qrn+rO8cEO
k0XwIhJi3+uM4cbQiIfd1raos4PuYC96gH4CB3/wLWDAHv1SH7nIBfRs2cQ//13c
fehhbmzakn25gLua21Vm5vzY8CD/HjjYCA/Wb/TiEvvWoRx7MafZRpBwkfLPwdxa
U7NhtRryiZeHOKZ30K+2RQgSh3GtvXv+pe4XEOzAWO4vd4BS69xUsSkT/5A0H+eq
OGWrSuv+F5IDws57ciHX8mCG7U6UazOCq/TojbEF9ur/wphEvQNGR11BtSFw/Bb9
onqO5F2G/DCVLmTeiPul3QWASTXzKH6b7JEq8Kq3ZvrIkGosDQSc8Pw0eAMdDe1x
dfj/Mibc2Yv2vkdFyHutVF88nbus/tYznYpxGj4nfrbCkWQ8m3uVdOlOStQGyoGF
NxcMkrgF2SWuTthVRrIi6E+0UkcrO9IgGv4wvEr0BB0r/3rFEKylFQZWOaVeQXyF
8HRasmICoie23M/DfOVJlGArnxLrAMM/6xKU3ea6MwKLTJvgXWbVwF6WOkavCl+b
AfdzDwfjv3LS+4E3460cp0un5jWGPcM+DJ5JR5tThBXalNBPJ3WHkBre9owdOi8s
ZwfGulQdDN/D4ziI9HEp5HLgNwnT7IyPD3bJpZnsYiX16ByDb6NW7Y69jS8sXMbq
/I867o4yeivkI98Fvlq43SiztgdpkGumKU1j9dXi5gaQjEhOkR6nXLWF+1qHyKO3
ekyvMKJ/n8dqijrVimCHEvciSR0XCPV4cYbDiwX9up/r/KR1OkFPLFqrjoxds/bL
nS5tBGeO9jg3dJPliXnRDuRxeAmJiHbMUP7QCngX/EqFoAt3c59rhBPGFLzIFfMo
tLMJueKOox76BfwAwQJ3nqJ5FeSk6Kwhwn6b+oxbCu2ksYPDUEjOA1Lt4aOlOotI
r3t30CiUbMelNI6HNbhW61pkpWNjgS9Gsn8RkX75ZLMo51/p9DSy3zlGEdqjhbxX
l6eCJyMBwOK7iUuFyBsBGLPXf0/iXR0dpqZAEcHYBI91UDLE+9hEXxRF/T4+3qEJ
NbMx5CrPVHGN4b17Zz99Grd2RK1ulwqMt5hg1baFlWoBObz0ZydLBbpffAQ22PwF
3aW1/u7e6tXIlwssQ0p+K9SUgC+7qPYpx+xhn6rSDLQ4Om0Bdw02w81qaOdUOqnq
Dz+HShydpNYxF4GJxnzgDkVm7QIPRQWMNO0q0wQdPwGeBcHuXE1cnLGyT7X4avit
m3ft1LgeTv5O0PAA405R07GnZ6xONQLfvbyIGM2nV+a/LSJUkwWDA9ZpgyUt1Gn8
FcuUtDzB+trXTiefx0Hu68rnN+ls17HF2AIOVoNuedxEsKMO6soEp5qyHTyxGZXa
NR8CBtmY0UUauu8PhHg5xwpa8cqJCSZ+f+YH3ah/+KNI2hBl+CkRHWg//KOm9AYS
1V04uFyzj8oYqVuRkHnm04NuTGSp6oKB+gqbh3eC8Il4Fob8lvlOdLhc+JjMC2Vl
7u98lETZch/EUeCK/egs03XuiuaagOEh7DTL5gnzLV/Q+ckEqOWBIoxwC8KJCNLs
OXLtF/eVRFemY6AUTudIKVjFHPgTJp/k0OjwLmx2mLUkxJF1VlgybXGaFfFwKlCH
BI4xqIyRWfbhnmoCA6i5uDoH34Ezi/a1JhnNMFVnXt9+hzZFeJmrzg7j8yx+hIQU
zLfpv4hk4PCxp7b+F5BYnC+Li6ZNmCMXABuEXdDgLj3bYZLeSbFn/pBXgsqNJnUA
Uz9Dop3xEGCNSOGBRA/MDbf8799xug9TMZ/j4ru1y3Cr7/4vwCtWJB+JgUy58svL
o8wQMerxO5V4lKFAvct5+k33wRf/lfDZZGpwT6YWhiYC8CJbafNfywZI3EnsWF41
UJxQ0nH7RIgPTCc9VEuhjrISxHQe756QWAw8gzLeMttB2lBFghDqwc65+U2BFtFt
gzh0k2XvQ2UcYiUqaQkNPjiySe6qJRH2bEAVn6Dgbs+WBHQ1CMw4gxrMBCx+TkQ9
lUcvREwiEWGSs0dBwhYR+7eERWl8oXZoBDH2OkSJOlYCKdozpOtvzMJaTyERcdDa
745UjGyPG7JFntrnuKBaltpla4VMH2v6/rgmwuT3HHy2mYd3gWigL+HHY/xpQFFG
+Q+IF056UqlXju6l6aE7I0mkr4P3SHSJhVmKEFKercDHfbZZ8omHODPOZfGvE3To
q35++6Aoer4GLtBDDhy55ENxtoF/QiCYK/d6FvfD8FgXE95HLQbYqNvdtG+q4NMn
5EAu0J9JR6RXsVkja38naSY2BZuEoS+MzODsX5L8gdwAPkY1n1m/jEYQ6mGm0KXZ
r5tNk/W7jUTcLakpCvuzauuR5KGzpB5UJiMHQWc4jzGuH4tTDYZblE4qvCV9u/6H
VfoXgOD3KtzWx0TcqcQ5OcOFu9a4v90RTEF8FrG7VJWCpGFqJW7jkr810l2g8gXD
Up5w25gTcFrC2Rf7oZR65oqs3nv7aFx0Re59jvzzbWw76OyM41c1xrzs/GXVD4im
hLNZeLPtyEvf/1Rd3dx+RtgoPVLK7h5JrRvXST9FdXmZpQSlmM5nxCr8recVDl+C
oFwz+7JkGeSvsVrTjNE8gzQPafy6XOpF+sRa0AE9uFs2XZr6mi+/iB1ixp0TbdSF
0iJt8/9M+dFNFSDOx1BIdsg9oqFUOguvXFbKtAk3qslFL0Y+XToq6H7VYqCebGN5
iJcIEnAEJrF7lFBDBfD8Xz4gMy8vFZzesjK0lXnNZn/SZbwA7Q0dSQKgM+Mkp/AS
W+ZCfvyV5vprFXAUy8sraA2avTDRbUQMaaV7lhny45cscnOE4LZ54SDRbOpq1dOX
4qJ441IbcP60pDiWzMqOReh+jW0tdw7uDNqPCf4x8hu+E4CfJIIurPknqPytwcol
igHlinrl7HNncczWlsHGs/Cywi4A1ql5oPJzPnXJVvH3gvD/FtFFfgFlWGvNpW67
QAywUTVdfz5Nay1xm2ur70qsMDGEoNNqs/FXB7hTomBeibb4CNM+aXPsaIHq0mbr
wde1f9ucC1uFHfxEPMJ1boXHAp1KIuUmclHNMXZUgxEni3djdz+pZtr6L5+mM2a6
96c3YzA2uEcHDBezBWsAzK6+nCvQ8Rq/bxp67rNnS9zXJ38BiViVBCXZVshQYxVY
ILJRvzOsVFGYeK3Sz2pFyUcqyQrs+ngNAibrT1buEFy8xpm8Hu0hAnVz9coZqqIr
IedWhYe0v6O5mhjtZ55+PnaX5R8FOekfk2ty/qITYgI17KH4FCMUZ/erBrrDL8ee
sdjk48j+y5+HijE9feEuK/UM8hh7IMQrDBtdHXzNlp0WEgJCrFbeN5gWo6g1jriE
AKbpvQ/FsMZuCaQmJBLbRfP77uMPQHoO4JC0YK/bn5BDwq9FYnzGbV1IWhoGv1UW
hPHxwq2HXqDdcEhKsHId2KgYEiFk91WSViNvsjuo4FVt/awdidOK4sBPDnSW1tmV
S29qbSFh+/UaQmwKwpIQ9CyPIVd9xftGtbwmTO4+CVhTYm8Iqz+Wmd+FtDB1rHGl
NDtWoLlogbH4oIWzOaP8goYon+4CIZRNZeRSd6L88+ZlFijMmKB3ERYPdfa6oazq
fO9A8zr6rE2rvuXbLlxEPZpGilvKNfOL0IyYgeMduHNzxuPD5LQe/uwXXHREQIAV
YUOLtjxAIeRYnTGEzAYiBL/IW+ffqObhZI0ctqXdATVF9EE5HELPbreSRhBrwXlL
o7sWxcUdTmNlZDpzMdfelGT0wzZrvavgcLGai8SmNXzVSGBwqt+0CCdttQEEom+h
qCJZqbyQreeArPVM4TIaw4b2ul9uQxBLXAS1cFTdl6LH23mCjE/2vPbHGeSmEmwF
Xyws7m9jvK7uP4feqgL3dYsENOJVD912iB14PuOV5ZsxXTS3AKgDLIVieIbZ9l9/
Gkz2HwTeGPMfkSoY8JnYTYVTFh5Bbtzc4JSii1uLnWhjpOby+sUB+ASxUt4irdXC
zonaOBuC6JyHraxXvydKljlgVIrujan2Ze/2jB1aikg/UcY4fyEvxGZ3lR/lkmGc
QfJopjLK1UhFT2GjbXSWw4hLoaC0HhAmE9DOfHbxptQxF/OZi9KwjhZI0TQfvSus
mWQntXb6ArkVCxyuUvAdPyJ2UqeW+EZtJYFIbmbBjOx1o6t5D63NDAcGGF+/5SZx
H9m09jAr3almWiqi28FxzKvTbgy50ziqntB6Z9jgX96kxEtM5YKPLTYnZ3lgfo6e
cU4P/vxbytK9+bTZ11Ptf7XpOdOF15XWb32R+aJp9jahI9BeFqQCJWUOagCW0Tfe
+uMXjVFjU6Ydyx9oGKHnaA6j3sT8blh3xpwaUSgFhMVRzodL7n2Ys3SA0oG10mSY
t+9EMMYMPNcvAE33lJ14dlVFPo6eaqd4bfUNFM/MQ++/7ylWNH121tHqeFQ7Xoj6
0KVfue5GsWe5DdPQ6uYYNHpXGvkPIlGFYf32fFFwVfw2dCqgBbyn3zkSnEye23sq
wDzsh9fcJmr5hksaAx8989jtK/0qZ470kZrV3LyUfNOQMCPpi//wb4yBvivivaZp
qrNTFHtbh64H6y2xDGuePsx6TjkKStyJv4rRYppTzXHd95WNnAKZl0CO/N1QIeRU
nGtNUyUoNpkyM4bB5PKrRB/FChSje/7pqPaEqB8u3D4JiicRlYj3HiqS0xu7gscW
lXLQ6uLFrPcgYBA8rF31+tTDMZnPmnx0Zwq9MXunyeKAqweNkbuuhvjPoOHGLM8C
VzdGuwa6GCF5uTvn+A+QYPfaJ3lBnKVc5XvOMTVcgQOBdbvxqKzk0FTmLIHYO9d1
NuHOwSsUc0aYcX2/yjQ9UF72wvOSV5tqXgBKJWhqE/I//Z04AmvUHa/sWSZBw1SY
GVYYHcMba6IMMhN9qiE2S+E7DRs/Y/H8ofNHlOMorodevwY9JDxJ5EZXW/+2cBQe
SGoyOTXdWhbT+3J8VhwVS6sSnVsCORmrEStWHCq+Q310G/zOomWfb/8oQ5oZvje8
jQ4mm55Vx/iPCFUHNI2Uaxvrs7+OPf+1fgeO7OYg0RzfH850j1l/rvF9grA5DfnD
I/5j68uEvZCMSJEmzTJ4wWLFqYQ+u9Q/u8TRC74jtw9R3JFp7z8401WLF1Af/PAd
R480DwUEpW193DBhvQFRrYCknYFUACSPMC1fdOyHtBZ1dtr6VC402Oo/F0CvfbeK
coPrYpjWONjuV9+N2xx+OPJ9d+AJqBrPY/9gAaqF9NVW63PWvb380ocwD3pPVo7E
4wNyzRr2Y3LC9dv6G6XYAhlctyCLlM7tSL6aZxSlknFtp5gfXIuMN1fh1N717A8h
LKLRYKSVSkn8Bo6CYFlrPiww6NN4uq8lPVt4zLOcn+GPGaYIfYC8aT5zUQEAxDLw
v8Jinq5f0eMQBCFj2Of2yVyCbMGnLOf30/8qoMoRp/8SgqkR0ctia1TtAXRhaasV
nAbGNosWvB9kjdyDimhLaJpESXnGNJaKnsE+0G9xblYGIoa6HSs0EJO+Nnl4QCY2
vVKcsA64CKWDoPapOQuIRoiLrrtxsnSsEuAQD7V0BfCPU7GbLursNfOBItL9nddB
eJWQYa5ntXi/0TU2UPhf3i4oYxOMvryccWRG3qmsoLjn8OHwSzcO6aleA11eEVe8
TQ8Bbh0v4kUaCn/nnZNnkhZhMkHbyhSiTDlVFiiuSZNf3C07BQwbDTFyXQ9H3kIG
OR7wd2FhS/Dgbzk9ynTXzoxCKXOISzseqjsXWL8cLU5/X9N29EenBf5peJYY6H0H
uC81sxNB/sXy4Mc6lLbzkQJum8w48PM4IsfXCNOsN6QqD2BtvyfIWi3SLzfAlis7
OAyTF191EnwPN9Wcpr2mjHJ08vj62HuCdJ2BYD/MrU78rtXY1Vz830VTXQD6lWrX
X/fCnypxzMtFuz4Px/7+6mNBO90sKjVvPyfkyxAy6ak/9BIL0GrdTqRWLio4PVzf
WfaNOWDFwnALGZVtpXHzrRhdVWmXmhGgr59G0MOFoBfZIsDy/xKC8eaBuRbjyk4I
5wagDogsV5AGphQxsxDpCNZww9Cz1CYh9nlqxd4CCXfy/J5rQXEy+44PxejwxYVT
AS+uS5Fv+Q5EveAnPLMhV016JTWOyVYXPQTJYMJ7ibvtzivYs0mZ167hKpr8coRZ
+1usgXAO0pDjf0L7g09Px64Kr8VUelSV7HTDsAk7zFCGxtvPt4bogkpXq6Nt1lZp
aBax2JvqG3QEEgxlVV47yoC4NeFMA2uWuLTlDrl6jeBMrRCw6yzXOKPU8IJJtinf
/3hIW24/TC388ZvGLhXOadEPLSxESFm7nBrCA3VE2RZbajl6Pi+4ag7oZJeK67Lm
cHLqcmn/1hq1eXOywlXHmc3xwQxL1+TpoGhHsIBCtVgUpMPMZ/oCsgCUAMAl0jZI
xnONm6jJvw40QjWtRl18iDBem+yar/OdhERhwDz7L4NGKgzUQgF4wL6jilL9Epc8
66ciJlHVDUdvbGoCHj+9Bj9k1UFEJZJJoAr9E8M5ZrNpDt0vow60C79s1LCZKrZn
H5zZ6zIiXudOj4sLCxbMWZwYCxwYDrkbJmjKCRroeR36Ru9F67bVHgeW22LiIe2S
2ADhUj5tmPRzLBke2JGwPq2345ahVTj3c6S5o2ZGjc1n6fGoPPFu6kVnS3/wUNRk
Q2N2C4lRc9Y9A52fCMzI9mtcigs6/SFBiCrIbcR8XRC+/CqyKJJxhOFM6nVynICD
NASB9V6674+Hez3XSc4uITdF+ja/+jD3bALn4u3msDVN3bsk75SQMf6HogKL8EeN
WThsymI4L9l1Utr/Im+wyzjBtKRvp+sO9SDwRFjmP9BjbwC4UuQ4prFK3mfLPXNS
1HslRkpd60KGolj/XrlHVS+N1lcgTkpHtz9XO/qCbeLob9c0RhiUqXOgjp5LSxXe
rXXPN1HaPY8Yd2eDXY/vInGFaRWjdpop7cNQOa503pKTjXryIG6egE4W8PA9HmY2
z8HF7j/sTR4v6M7oN3b1+3XsmwenKPoHRrl8iYIrR7K3vSbNcSPawLcLFZc/+Ex3
VIEirjDaTPBby3mwRbPJeshjCaeBHaO9oqGpWXt+yWJPCszuvY2ObOdAxWkkxYuY
rl3LHZhOldnyMfvFYf9RkkqQi6YfXRYKF38MaT5/1/c/61UOG7xQrV4WdfkUi9vL
hZEjen2U0Mjh/0lO2tBMMMjE8Q1gB96w4bseQklYMT9mz7DUx2zorlfKRyCwbUDl
nNvt60YOHWqOAIeD0jZT4vsgknGDVf7yJF8/yi30DKcTGr20AjSG9BiiTvqgIUoo
DCrz7WQCOyRFgGNhaT+pxQ75x0MpzBEwme++B4rKecYVsQ/gFIFNcKipJUL+xltK
U9gW5URFU7Wj8wBl5GXdB8wZ00lkBcsppejTRXjfDlrbXbFec0Qsq87bYTd9Mpdj
zk+p1UdCUZUExrYvpiYAOy5KCfeXPF76gy7nqgr59fSspysqDAQNdJ3Ej2Wcf6wY
r012zOksmewbmTahu2je0wDyhi1sevhrxmBbRdguYxWr4qyDebx9vI1w9tVxKjyI
nD6RMEgYSuPZA+1AW1JXilajS7OK4/Xc8tvWdOX2PLb5YMMQH/B3MTn4BDB9XF18
wnZB9SpuLZsrc1o/vZklhYb5b8HqluDCEmOLabvlwzNeyP8eZjB2ZOXIZ/bv6EkY
L98UvnGYB/JkZBGXJ014mu62dtGOGX8zCP1XN3cuCWj9p4dW50mu0eL+WiBEY804
h8UPTrxfVuhMNMvZerjQnXgTiYrG9yNw3UG9mPBKFvlFSLM/9zrCECJejoz7WmH8
0YCejS2Xj4jZe3XI3MkkcLn0gCCC8WXphJIX43g+mj5gzLmNyQc2ljSC+LPYRwRV
WT1NjGkj6fiMnjRGE5MRjbygbTqeq/q1aMO1p1pjnlUQ2oc+K6mPj8CD9gkEwe49
hLvMhA9S4c6ZDjnBMKbXtSXTDc/xsoVZjQCoGZN0Q/r/rFr6MvGLfIJCysGc5Gww
hEcxg5pJ4YMtSfaidcUxq+NMDzPRvTJZtCPR6wF4sNRVAA1V0KSqmmpO2tlq3NTj
vjerByp303OQ1zrn7TOXDSuCoYxeLUFFUjuIE9DZFdL2hEUEdqfJ5Pn3LRNL+Nu1
yld4iYoB37/AA1jww9hEzF/stw/tWnpaamy5NGM/R6qWNFEFTnphGQaCmu+8JHm6
glYJdSkAZ2+PZuz+BjC3m0yz6+ZXblmdzI7LCIrNTHrTJZ75Tvgmsi03bh+qRFp6
qSYc+aTyJLXQykguDtHrFPm6n8QBRbbjLkEnHhWg2XAre9lQE9EZspAb0illx+Ab
jnlCAuFaS57e9rUaGKswKP5R7S8Nv3fXdQVzXHUGfydNmYFq0dbjP/7zLYtX4fRr
uwjVN3w3Ngby78edb1CcTqsMKRM0TrYD7uobxFEprWo6TmuGh12xi3hUZoYDiSIh
DMte2wqjBtiW3tRafmwMOC/KsnKdFxkQBSORsRDvC/8hcHlwwnPrDyuIRZ5XcmH+
ePN1Voh5V5BjzqEuSBBV/Mneg7WqoUMoEqtNBPwFqjsl9Bgb4GyQ+xbT6R2ho87J
aH/97DSUJxpXOQIurb1r9p2kQIoWz2YDXa1molvSc/pGMxEyU1TETv8rUuDJCYWd
S0Jyz5HNJUSfQS0f7/x8RZnzpeVPGzg8W2bT4/URxO5eA/0zWE+syPUoesw9FAam
/TcAELb6F2n+nqxWT9dGQLpllv9MstmiKrf5pnJD8zkG47/4z9VdDmUmWGQhRLDn
t5/eecYAK9rGEGSXGh/CtqdcDHrbIQZsFwQBGX7vWwrXIznEbfevotFTXHMknwmB
UkEtDY9kDLXGSzMwNXh2dU0Vj1s1cFm66xpuXFW6ZX1xHeRQGd4xpduHNO3zDsg8
ri9A9PRLtdMz/+uq9xzQFKTf111wPICpoiN3HS9q/qxjxbN2cc6WvNJmAt/cqD3L
fXk1xqcbpP7iRE3jJbo8hsd9zkXLOpdA+tNVbsK2p1Ch5woSvpGjxAJs8Np8Wxqy
B+fKYwWRRtsd7WDYV0w1QtjBldlyW69+al/KvCuq/NUMSF5YnW+Hg0bpDyRqCoq/
cb8V4I2ugh8trrD1LX1cLJ7+ntu4N6miQx58fuXDpgEgi8rT7o1FZLUIkOZI5LPp
KVVcIc2crAI/6BYKPXdDqM/mZwj16nPk0NsRFnnkXN2qxPKAsONHZ3TNfeyZIaX7
ujh8bP95AoJ3Ie0XLd4plL/AgQfObymi2sQh/YKaNF9aULh0sj5Wi6LguWW/mI9c
6xauU948pNLk6IMT6la13djgMewJiY2eNcWh1stOT/yLgv5rk88alE1lF4nhCwYC
DFS5nnUUeY4C/D/nGov+XP5sW67TGZoM9GH4vQJxUsTvEUFfoM2wJvS3xrXnjkH+
UAUKFfdCsdg+drsyCZnpGPUhBATN2MpcGQwG4VEin58BX9kCgujokxq7Mw9HmOcu
4w5UXApN6wSE9zIQ43eEWPrkmbgEZ+cD6q56xVXrQEqsZCmdONaci9J2owUgUTr0
MLsZQqEiPOI39ONWDtYeLl3fmchqlEpnFGQRyr1UKj9me4+V6w32csXs6+y/yTpc
Y/CJdy/CsDTZTwBtvEVHspNePj2lpE1tu9wjrqUhQHMjeRWCUrxvFSia6dBLl24R
tUbl6SsDxxiRW1um/LVwDCIGXhFzZn9yK0uFNvmtLGnNISCdqmF7OAb0tblhiTqo
4s1F/Ay4S81KuzHW5aq/1aBWxh8fAJD544+tf1RUSOS6VZCRkpYWMNA0/Xtf1N+g
2oVVQGsHxZQk9xp1ADfUlKCRdqxP/G2765X2oyKaCqXXfGsLgpvsfJVqifGIm9lL
nSDQcB0bdAjJBJHP1A9Oxt6X5UtVQYDdKkeb6nsD1SRkEBX/3WrZWXsjbUozxS4M
xufpOPdyktMWEIvpTn7y2tayxfbnk58+9OI9AzWuUJK8O0d2r1Y+oenv4E4ZIt/b
SrzH4BJZEBQNED6veec9h5JRmCrgMTPnwKmtj6L+STgGuttlXd5+ZTW85i7sx33k
9gHwLK2czcY0MdVCIQs+OU7warSXC+v/rErKRlpHVbFcUeL7oMwze9P47RWRIzCe
yfyPnuqHCEXwzHnPfxJe+vs0Id9me/cAD7EtdCbCN+XUOXBGsGgglKdxSVG/3fGY
6UascTw9qwFBN58itZVjUbsSkzC3o4EyPy1GSteH1fB7JDInXeEjAztMTRuKMNy4
04J3LOLutHNR68t4/+XGLwupC1CG9a/VzcYWVST5fAmPY90DY9aX5c8V2mo+I85n
kJkESPWsQi29ITLBRW96tqDPgUYGcQIj4hfb158PYtOepRrK2ECGGphyUBcpQIWL
XGJRMW1diJTgYKP0Y3zgL5+9i6yxF2MoQYupJdEgJ9lo42d9Nw5JIBud6JPZ08A0
JCNBA6N9dDkFIWMXsciZEJeWT8leiQgxYBWdilENtdjaz3ZqXZlT6airQOuxLGN9
GUJlmb3t8bOmiJeOTMoqzVMZ3mn/7zOXGW6GszcFAotCuqfwtqY7DzerCZkmT14i
YUVZLVrOXedAckj5GS8l5/KCfKpxhOM3w+GLYndZ2btpt51zVbmv5ZBv3Nz9tDSP
nohYr9fILoSchQxkG0Y8yL9H4PUpRvl75/8t8POGBifMTznYUhfArv2XDylOFcwE
QeO5UqPtFz9d/WIK5FzYUWPag8YuJVdje25dtP+RbojmySUe0Xjd/WUv8Suqw7Cb
le0x9LK2YxVrcryN3irK0LngfJz5NrNts38GYkZs0KI7luZlNkdJPCs3D/BlA5fj
Mpk1yqYMypMHwSXjCSj0OQjN3f8q431sasMHYB08O82peiOkvfwWfDr05WuLwLp7
TnwHxnfzJ4A6EfHTLq3RtWc2WSwufaFZGqW2B+X6txSfR8zm661UOMZpylIM+QC9
MA+yB96Iox8yX741VIvbJKkXoQtk5CqGlKvMJrL0fRf9ZhkorScPRjLxFls48He+
Rtru0BMlMwUYbdvqZLmjZbajkW4+Z5iOk9Kg9KkOyEZYPCqi83ux9BnL4hUQypdq
HHjXophnclzBKlNHdtZsguEOkVclD2nRqoYAUYBUH9SFje84gcX44BmgL2rk7Jac
1Iqc8J2ITXkrmDFTWYdj8XWl9QcPyO1jLVqiCW3hslyZkJvxiVPjXkvGEBOdEr0f
Hi/as5YbQKjY0AJUuCGwooJk+32hDJ91vFj6N0WZtr9QxkFsF65AEvWa72FsC2ox
Oi2Qkt4gW2T6WehCuomiFEuafKaUWzaeMqy0kPSWjhRofLXDp1x9WkEeUnXs9CbE
KjZR9Sy4e7IKDQmGSER0hg+spX/YXsSkR47tsqrrg3PV+Pw5eOH1cBpINiWRcURu
mHFaFtAGyIyDDydloJ336bH8jphxk5SImEclbwb6aEgQK7Vyqz8OXumFzaq6mPGb
dK2LVEGVbWwdgvYhJNrnmBZ+MT0LFh2tjY1r39VjdPJD+1A2bcs3EpzHJrlDctLK
HuTxLlxDhjBBhqPqUuDW8TS0u8sCHe3yzEeNojXg+3Fj6ToEHF5BkXmnhjfLVmHy
HrzwLUQvIMGVscvj92L50/KNJ2FMUiNfpuOLrT7l5yBUR2ERJwQFYyvGptHwH53u
qP4k6bvCOMxfbEWa7Q48QHTn459jP6aQa7MO+5gbqGCOT71a3U//fy+OIsfPaVLe
+eUb+353hu3u2xN0zQP6Vv4uFxqShWvdFWb8F0c+UMqv1Dsfz2/dacW995PktWo4
+1yraA8exOqI83ezIz0kiutFlD8ogTtfQC9jfSbl2CbiuLkKrcA/rvfqEnk3hX3Y
cqNVLl0BEHgYCy3396kBLPf96WwgtpRaM+LFynCS9Gk1Jf7/nsj2HFbhEvWmHs3O
CWatDwFmXAZ7xDXMrzVws2ag8s19fWELz6t+JDeVsd40xCsg7BKWEjmQVAVQcXl5
FI8oI5U5kJ4hMC6CPxSC9uJGiK9Xwxf5rOPtzpJhVtimSwb0iJW/oQwFh31kw8gF
kRWJ2kO7Dcpaspo8+MTLRpVZoCynIgsvILEOcH7ubLy97xgmb+sJ/iiri/iN2VbO
B3a9ouwegYTBsEP8irzZ+s/8u4hAvnSfVX5OvC8r3QP6MMixM9CdW7s17vte/kBy
NvIVB9oRKIaSfiunFc0bg5B6gJZ9NcWyX7TdxcIzdL077Pi45/LjyokfKv5NC9tx
MoZ58ktY47FrwuYlcly7v4mYOcC80DkJ/xM4pw7ueDE8MRC6fmT9gZSc1FDYTllL
YG5qLYFlQEYe0QdOMVHdnCtqcbhiiy7VmrJhnjkiKrnAbT0o04DWEjaIKGObrdQJ
TeaPl3motZq6gqiVw1x7qO4Da1cQNXamSE2BTM2imv0vT3xMXwLPqfbMb3zrUi2L
VbELogSULRvXtT5nREJbomuMxx3F+LWLPxZfJsCIUBGaENq3iqmQEZPLDyESFmng
BHOUyYG73GqbX1vMzCb48bC3psXEo9EyprYY5rGW2b73s6V1Cp18Fwv3z4K8rkTa
SHdPwCQTvMQcdr8bK0jio1ocE8PvH8s8PiyEoBpEeh/R2294/8ueCHqPwQ0qXlZE
i4KOtSll14Vt6nad7iEuwFFpBaeOidBopjO0/Z2gvMqk8mLAjXCxL1y9qRibiSfu
mIFD5YFTJA6g+WB/u927+U/tC/QMd506JCT8tceX5IKpGXpaaGNYeT0Q+znC3Sdg
CokfYYbvRhM3QPMfkbBKrQT283vWa+BNlpL2O+XspKJ35AaFyZEdf4sRwYLJazDt
N8YEKeTmNAGV/ZwQVkCoz0DpaICf/liPyD+SWJwYlLZ1Hon7ZJr8ZnTBQV89aVW6
zCzd3aEg1lTB0cT/tiMhMRUOfJVAkFw+jHtE+lrvWvR9Ow3ermjOJI8wcJXJWNc3
NWwfssKUNDqfs114H7KOSRvMXOAiXW346Q/DUhhotwmOPwHSz1Q92QKtYUvDXz5X
potFMzq9Hc8YZfIFwts6K4r9urFw6lpYS3rzq5/iDmTmooNqPaH57WdTPpnE5WXo
MoKlneEQujjdG0NIrGV8Z0GwoFwp64aaU3KDb3YGZc2abT3jpySNmTfMAgnC9Vfb
iDQCiFw1nGiSwwQkpVkVqzBA684YXhpqNrbYu9bI9sFFU9KTUoTO/DuII2hAFryV
vAPN4PRksm9RGYcMex8Ajp53z0CDsU1Inax3Rvy2UnmUDRMK8RUG8j5IKWu4ai1f
I2tgS1E/i36tQltWIDhi8P9EcZWtvB4TOz/e0CSg1Df0XSAHM0hKJkNzy0WlPPSp
RJ3uH79wAVnUJfZN+9MTrZxIj2SIwiHPOT7XWz91EDMFQ7RehH+Lzb/lougyq0SU
6g0TTlbigvKgeBc4s9AKAUpdnM9DIzDaMb4MTXAp3TJbpj0xsWQvTcGAANxz4eI9
i9lGlR2XIt2TwzdlZO/kbQrcOiA7WnzyOMrFPZOQUSKXBGOj3ZzInx5lcdkiovXK
0Zeirrx5o1LgjCgy8xzcqi+Gq5IbX+iHE4v3XhGTx3GJHErpKBJ+jDQeR24SfQCA
X7Nyn/02ew5En/QS6gey50VQfdzi6ShjWW5a3KWv+LGpSc1+WBSMKPtlbDrQ3Chp
5goa0kPRSL92NHmf5sujIGvXnDCYA67gSq2yeKFfdZnOPmQtXyv5l8aD3S2UtxqA
p2SSq6sFViPt9nZLl8bpugxHVKx6X/2fNMHn9/y7ZtbTcSPNeN3THpSOzHs8xXn3
/MDhYcYNL1UWexyohEyxfGqT+46IEkQuGjLC5ChVEt00FPVEJwI2uXPl3qm1QGMC
2GWpk6tHqoKPwZwgZSsXKlpz0XklwE7ypKqeIdZdEuYt2u50Vtn253OEXGArZEnk
jWETx0T7KNu/SLwHMSkaQKcVNoUcYOJKcPI9uYpZeqrjLEHwoBaXRnOD6Ptgrq2E
8cORn/Buxm1Z9dIEkXYmIrhUXjJCR3pXtsPO+k2yiXtYhVAfU6uvamQC0gQFXgiv
TsPmFbWJI+tAQdGEV898BVQOSPLk38hVUMhbiOwZpeB87lvL0tFY1oeDIhOJv6YA
TxA7Ru/aoHgm7ciiN/RpNEIIheB4J+dGn2fTc+kmvCyBNsVM7CYlkDRzy0UwXcT8
5B4mq78OtVy56WowoasMlKwIdZt1F1I2JTmjbsWNcYu80TOi5E07zAivuEkqkICx
pn/vcimNxMy5mnPpG2sLGxtWG+eBiM+wFkwViZje8b+eOa/rjkD/lybnFVo964mt
6m2Ca3KdkwF7X5fZ4iQ91s0xvxiqw2qNo1LAHvk0nePY7Z3mp3p8BQNf7JxvBc5Q
OeV8oa78lWSgoZFs2zzMrfFbTelwOOg0QdtEB7xlnoyseIBMtlK9mvWr2GW00fQr
m4az5QViIwoD6ijKZbnKD7ZFedkcoXcFeGUmzKnS8eOElHpbkRvvHQ6NKz5+YiyY
Wsq9m6k59pHJgOJcowe3njYgjkhCRxYgb7okk+QUmXf7aYnd5/+7AQTaN59km+pF
ohEb7Wg1uZMipNP1q/5CLaVI0Jx1pZjxI97xKVhlRWR1Kjol1GHZH0T6k0DA0tCJ
Q8PF5F1NSiTInMQDcTf2O02BbtXlnBntEhPsjxrp3zFwgY+Na6ZRNsuNNyM53pDr
WtaGURBu2NKaA/0MxxHEgGx2oSejCqywXgDHAKF+w3l5MOYGWZgi9LVqlHZW1aUR
SfFD1vacPDWdOm1YUlNWLSMc15UsXn3U2KpAeHTro2a2maulgxUN/bgma4oKoj/T
j+s/P6mKFfZc0k3t1WY6qKfLH6DctFQj0u9UVdJXFsnMiTEysj1RJgQwzC/akdPg
zarcmGxzqZPDu18Ke/VNfRovfwB8xX2zsHjaolEh29XZr586SFlbKQ4opKxPWKxF
kXjHXWDm+fXjwp3sBb+fWS1EbuoF9TeaButailBtJmWg3Fn+Q4AxAcU1b43i0fKz
zFZuSrmJx7sLh8IihOn2fejUh4sB28opigdk35SgfHXTp6pbLGvIdgr08+8khHm1
CP8loRfW3IkHGduyeLyucuO0yIam3vUw2gUwl5V/pkwVL3m/0oKR0Y//g5LmRevj
4SMnsHXl8IOthFvl5ScOHIawk0Ut0AIgyyMdXbalnS0SxmS4VIJj83+DeFsz7Koo
36ubSOzPSC7aayUsr3SJBCm2wCtnm6tNRn+rAIDc3JwaUK1+MtXCvn6oJpdCc9vG
ZOrkt50hbQm7UuzqTtiQnVIEcN7Wz7oHFDCbwNz0govmPqpn4+EORIupCgfea03Q
kAHFVx8/4dSjQUQ9zCwGh+G4X1bfuFWk2MAM3+swYKrJope4VjGO9VydjYIIZaY/
vSaCSzb2OIEPE8dzyRgETI4H+DYgaE6alK/9N243CMo25bWlFgXokRyY7B4+Xisb
YRllk8bKq0uV/kPsiyV1s1lgGcW4Re9agmPV1yiBJ8A5/yU5agvpUmpHBK0U9Zsk
vsq8SCE3mjKuYs21K7xkqK1ith7v1kfZfj7GbMv1qchc8JcNmsWcsDZD9KzPXy/c
ozTzxWI0lj+ejV4QxS9HJSaWxQJnpvD7guD9I25nsr1o5EfOtCYNGDW2A1SkMfzr
R0KXdqVwHKuXINyUh7CxWeiPBc1x86FznafY+C6yVI6woOsPIFdRAmg3ns2BEZ7C
37wyBNVzcDqV7jH0zyWynRHZd1fcvCHs2tzCIKn4cz3glvdxibyN2WNkhpGEVNxT
IksO8E4fmGyGvBSiVCUjnYbhnjHwkqUTdMM9/pR699Xc+J8CQdW5EE/eBzu44poX
pX6+bIBnhweFIcR/tIbrH/JaUbfp7yEzIr+v/zGOfEp1OkQM70QFwW/BkE0CUj4R
H6eRqGiOxFZIH895SX9OSINEyo40lRDa+7LeymKSaa0qls+70XiYTf84DAM0lQfB
01DLHcfGHkreyFybyfWsOncMjuXtdsbwD87sMGjYu6+PHPG6XTtFEApm0WLZCpWW
JEW4nm98p8z1bS+KXf/niAPkqvlXgOjSMY7wkbEt9c2/ODxNELrr5QArVgBQNiI7
SEqZzSBcv5lLjaDh+0Lj3ryWMktkq7FeAeqwxZiLaBaXeP4Lo+RDpA6njv2U7zVn
GmXXnP+5deP2Cii0g9+sR9miRbbEde0AjHz6VLCRE9Z5qQZdQbRStXBR9HU3GQ/t
FS+Onxj4K8P+cYslHsKPU93xWZcBhUDILpGWfRHdQA+hkVp/aJL9Wwx8bjEzw6xl
dC4wALdMfibjriM/EGAN9ZvUbVAAxEzRCsTEed4h3hxJjQs8/np8w4xQwvdXdQN6
HLLkLn5Sjc1trGRwSQHPfwGerU43koHmfNxBy2hgPZsUBQXkgfLrvPH1AVJb2VfG
+4TfLEnJeb4Z6HgNyHlmHiNUbNuPwyoCAkM1IrFlAYY4d3nf+ZHQQZOvMBHqHese
fydsftCQH1ebi645Y362f3igEEeMlwbnRb7/iRggkMl2YrbmzUJWgAUMk6rXV+0b
C8nKBDm+YNLclsDAH5Gu70AM1NnwxC902E6sbUMU+e7JqSlc0whPxSNg3vgR1dnN
oVcy1hgjOQT0rXF1vBAzhMgPRtCuLJ33ku6UzWi4dWqp+oAabrUQiKhn1Wc2ykW3
KAetsvnZpyYxwKjY6eRCUAdPyLDKx/jWHqC5aC9/ueOCvk1/m+unto+r9BLH+qjj
drfGZ0ivHsXhv80O2AG0oEiCSdA/S3V7c48jMMqclzfJxm7+gBQoBIrb0icpx5oc
pcan5WkP6Ldoo5OWCGF5H/Qmo5T0BpOwDfEFj7+e792f8BZ76P0dRXc9XKZutmXa
fh+WpWJKVBifirFEsYEWqHrzx52+24z/6e3KCE8N9yKwck7bFG+byNXF/lsqk0f9
gufcAwzmsl1/HDcxbr3gXxHF0XRk7tUos08A7BeH5lIwcbYGXRdkDxbcQLYYm+6V
MAy6780yp4nH7szk6CLV67NuNUa8R4XHAsDbVypiBKzlazUcOFYSs60IEyPHa8QX
FhV91Q92KxUVRdLiTuXyRAVGqjLNgZ/L2uo/OpVXSzM2kXe5deKB5NtNRGQ0RbB5
XKJHZ/TnY5BfI1s6WISxQkfCbor8QgxslZD1jWBRqK0S8Y/J9hpiilbVCF/A38+7
V0sMxSagwlyk3xAAPdetx1d9nLDcAkYrWP7mhqCGV1FzXXIhIqcpDgkW6ols1qY1
wKP13T/NoIkQX4RtGmbAB9JMO2IG/ntgbblAD1CiO3nCal5hMiz9Pr3jYFxdxj9y
5LQEW0rWd4VyfuabUFE81RfllxSz1YvOHsGHIpgZ4b5nqyIq7QdWF8GW1mfS4O3k
J11cTs+iK9N2Uh8L4/LhwgPzm8lXJsLKWaP5xLtgytesMnbmBVtb1WGH2Nu4Fu2Y
cCmcJ7S2suMvaEX6QvXNl5fuyvEZDHgSNfXiUmfnyO55pkSj8SakxsUfNtABbGaU
tHrgH5DOB54mNFRNkgolLbn2L47WrrJ7ZIRkXvZC7mtqTGSzRqOn5V9Nti5cJ1lw
2LU+GcKtkbxqF6K6cuVQWkMQhsrlkpcjtPEbYQEIQDNoFeXVYIOIaa2UJa982NHa
j/x/W5kq6eOgRtVL3C3YVdgwieYcD5zdKZYVlGWeY/XYs2pR4JShnAweKZXhrh+3
DbyC+EbTNIGJVWo2yAklfuiZyOAv5GTGwbTLzKQ31/Y35MCBNeuslXmT8LbBO/u0
adVP2YZaRaDBqr1uAcCdGTJKU6P3szOZqx/XAgKeRyAcexSOjT/MiygFxBUBKbhO
VujVSPiYQ2MrKb9GyOEFLR5FWTAN+7eCBcGwp3ZXkeZAsjoO4v9msai9vnNHWsKp
cyWpaiC8HnrVb0wxpeneRh2WHksZZeEq2VrdIH4bCYMreOUQsehZtJPpDsDksghp
iFmCwlQjaLLxhiu+Ucrppwy765Dw8661PAEezM53MBi6gkEMlSKf48zBOcrx/qYz
JW+fCDxZJ+iUBFwPaLU3ZjcDG3kzCbXj2WaxvC/a8yyaRxDxhgLwNQKuGRMni8qJ
geXnYRKGMTR5wiUUVKiwyCSxBOMoCiA2Lt0wZMzIxPEGYsc+kt5v+jseta6ww6sn
OeA31UfCGHd7tnzNpDaLz3qm9ei+twv7hAOGwaY0+9K2H5my403L++qAZKm+yBRz
ydhvhKSUlIxJ3KdrDKUZhwJ2FeYf/MY8wQH4WL5dAhstapGM6HbrUSTcUdL1Xk27
N1eYBdanzWGPbZRlV6kVD4sWbbpOmnJUiNdzTpgNpE+069Xgakiexc028/1yZhcV
mq/zO19VbQg9I/MeTo63elSFL9F25hgsLp5sbwFsBEy4sxZA6i2ed0tFB6sosljB
Iq+ZACPJW42xwQ6bcullpYm7s/PHMJJ8YXTmWozSURP1qi9tNP+1mxqq8cPFimTv
3wcY7sxy6J7JAI8wyLPLOqUPGE6ltQHrHNRa1hg6nChFFYowyH/wvsWVn5L/R4QC
bbeOfzeqd/baWU8f247ExSKn5AmIBv6Kif81yy1pGaPpl7hSl4Ue5W9cCHg5xnwI
xNnCE5QA+zz9F82K6rsPs11nBGBmocEO3sG9F8mLvXbujd4nLgcIa/sWIj3ggIX0
3vTmQXm+NUK5g+iuW+vqATFuNWLXfFmfLH45YhPXl/adlr5PBBUj0Oxa0+/3OUZ8
ga2ILs09MPymm10DrnrOe87D9G9T7sksF+9Znn5NYCKm3t9UpEYQMlXC3zo+zGhV
pck4hjhaU27ZJ/x9sHE5UAoeGsDDGPC8/lwrXMd48akRNetJ0eUD1TIteUxai5Ki
SC/lq5baNZAqet8elQervk+yYZ4zt5/Tl/v7aqC48d9YwwsJFXJAlhW+q2udwq75
egVw7OECqJy0oKPFqVeod0rSgestFuvgohjw81i7kjzvte8B1y1q0Qz1qI7/M0tl
THKj5oRBs/t/AjmfQew4c8KvpBYWYGBwRQK527sAc08ToSgeoiBcprWy4cpQAYX2
a+/eYAIKyXFNf2hcNhEtGgHoTxB2TXiUX1SLs2rWOK23VFFGOWx/ct3faZZJ30hO
cMXmWkfxEIGuMHFitlEh5Mw295/1dM8mNRDOtkuoQhJWtD5lVg2JOGgA3zq5aJ8b
qFdVSGfByECJPs/76O6SAj46ar/SLTWHKykslydU0inYXZ2Gj3LE3oRxtlwC2Erq
KjXZ7ASWRheTmUy7ICR3BZOyTrUCoNnH2D37/DwnvDz1fuk0mMLiVgIfxqS2cD3G
tj746j5JIsrRCBlzeKVuZiF08SvhXuly42fxepbQxo6al1O4/YRWQMBljSHXdbfg
c0eAzoxE8iFhX/C8z3iUkrPo9cFMNXciwTfDjSWRzdwjLTrclK/RXTwe3RT3PAT7
FlVjnxyHR2EUImC/2WSMZ7XaYR9rEhVBOPA8xaPxCW9JXgUhE5se48f8dss8y0A4
qq1yJEUJPIBMaJtxfodQipCXRWxqcbp2UX/HIDK+L1mfn65K5dbYYgeN2xtmOooA
3u9Wh/PqrKOe50Hah4SKNwk6RFE5YdBkoL/9MnyqMsW0IY85qWApAMcUY6MmYrAA
lQQjltWfBHhYsiIcq4rqkijavfuOTdU7up171t1oq08iRjrUw36x8nDNTGhDt1ZK
Ushxcb8r4PJmM4zqVOBL3LzvSA3ogG9CiZBJln4tSfOY1dlTS/ONRhw79Dyx01Es
J0Z5t7WrZppGUxe7Xl5KDLqFuPExsgHeoUDFRkxOTV/TeIAw0tEq/OGvr3BaazNO
qp1kq/MMT3l5OJbchcwd5PAHoNxCsCyAY8AScR+huaMa5BOfyoa/KE4/frVV90GY
uE3ATYgKLNuyunHR03MczXokhJig1VdmciwOjvO5uqqrtgRBacXAC86Oe4iRt+R7
wGHXGIa0PAZUndwla3iIpR1dZzK7wlvyRmQgggNVydisFdfsaJ4H5Zr2NvxwQv2I
JCf6M/eFMy+PNpoHD5q/UmZKoe9Uo9mysHEEPJoVeA5WlhTECO2UGdpf82OMKam7
wY+zN/qN7fpmpQFHvpI8qtdhWaKd42vklE3h0y68/ldiVtmxE6c1jOumigqTMluq
plz1G1s6xVxGBGdq9/91p15XyR+q5eIu2NOj1t2vsxBZhsC1L+fxGhzFJH7CTBun
080cSrbYyISpqqyHKJ08sUfxAT2FrJZR0xKRIyK1czT1i61r3VNTzKi8KMJX13bq
pAzLSBuU/ePM/zfw05+vqM1rh4K+xGlW2qryCsI0rfswKtUt/9a2QfbY3w2hmR5y
IjZpXSh9pyBp3GfEndNEWJysk1vCiMgnepzmUZzPTg28TkicmFMZHr7DL4hxwaKV
B0oZIdvpkM98SbxxsvJMumvZBtFsP+Oi6of+y+lrJ71N8GWmhTlutN9NAL788459
red0yhQeOeCLFqmVWuqpen01+X8z2SZfFiSwaFQK5ciaWG/sBZE6Qjy3xWRXq7yC
C4LN2X1yKlrRPno7NRkTnWqz3TVnAYDpMfhC3AUPYBwSg8pCQMXcZtRIbkx4GZiD
AZXxcNAhBeTbfFTsllhasrWvNL4JO4SIsv5GYemlw8rVkFjfP7u9sboxl7cVJt02
9Pnn3pAXSVI3cWUZVUyWuctBTU3DpoGfnMredLMb/DvD8TbnjMs+ubx9qNec+rsP
ARbboTbUjkVg4l+nAoy5kZwQvzup0R90BEAH6OPduERXfwMIy+wKK0JOlhudFAkN
APYM2AiV3M4F9k5TVPaqnDbjwiLqOBU53eLOOulrPpaiVtE+4LH1+PLBaqpK5GJ0
eT1OoywQAbd845rBCkTE5mjCFJprFs10i5iDkN64BON46UdI+oaiyd46yZbViOgl
FWvfAV32Dai1k7o7HNrvpHl5Xdk2riYQ+jHRcqvVioAwU7aTUHShShlndV/iUteN
mYVt12CD7bjFkD9wbUOE8AQwo3SKUvdsAoqnRegA3JLPv2u2e2+klibaMQsv+V21
f7Cz4xmtGc3tZxXVWbf9pXAsqM8b1o5eTWp42k/poUcWtTKkO9pNDJUUKSBDxSmV
7ZMr1k9xEXBnthTVMU0yU2dL/mQLD2N3M/k6hv/Ck4JVLx+qKkskPNst1iPmTpwZ
YrNyWyQT0nhR55MlQ4rulXa4KG78B0+tYMPRL5lG86BQXLR9zob20FKj9AYKL5eN
bPIqO5+coexORZ1dkTH1auWYcDqD8XP7Z5w6kPgmsxs7IkEHbMs9eslyDZbgnii/
ex/AjZjDpd2N/0vlvKW9gtj3XLxv7PkFiFUl4cA4hUtaoR2P6QBf6yKm+htxK2jA
UNHaml+LeECrIqft9rd9V3Cmux8DpYelnMHXzUQ9mb9C976k+hgHyUHMMfaAa3I/
hbwchMZfngMVhmKfwL4OQtwS+ylrm18m/V3SgMSD4G2Jan4DhZKuVLqmwHWU71zL
nsZFRWzWfFz2xT4xLaHcp7DHleiHk3nUbpjCnUOmVgIpTXxCDCARFE4IS/B11c1x
WUC0JuxwhBQOS3U25vTunpztuwiu2S7zLxAAzt4aTOppelm8uSOMXPbMKofRsGJC
sV+w0VDoGxB9XuJRsBgU+zXjrcn/90svV1B/wbkNbyi/Ib6yOBiowF6ARm34l2gH
h+ZhyOokGEbNIYmYYar2mE3waAZrp3UY/O2PeyjiW/MYXkjf9iZKWZbU6xbQ63NK
KLLqEegzw2chETxyta73KxqdDATqpuZMsFoYZR8c7RVVuvqEbY61ZRDFll3WFZ9s
ozGxIjPQFfUfoja6KuucbSloIulTt4fvUse4Rs9viYdr0lbZkUkQewVH9KkuGuue
SGIbC4+M5GCBE8s2xWq052TKakzXzqE3wF+CqPeKpYui8rs/mj8Xw2pbjQNrEoQr
ZRl82HYHXppcjP9/mNWLgaSNBcNHBcFpgtro/a4fUPUiA0gVAbx3LiNXY4K9YsFZ
y+v6Z2qeJdszFvhUjgLy3n98qqdweMXpvFO4kgKrlccOV6oSD3HTiApyWP1mm/K9
3fchoLti5u4CQ57Qt3jb1klEDJE1RNP8amFykCztZZCyY1+aSdph+V1b4kQWthY7
SPZqDLTiKlE8PAdbdmP+Fo10p/f02DZkk+84o0GX4eABb+OoTQKwh9nr4sU/uDFw
HgYwwkMa5tl+9M++qPdFE+s9bu+fe9lxg6kdU4rjHUU3gEoZ5OsVd1s9t5t3cQ93
9XCiHf12XRkEvwCoHunFieg84yLn6LpwaGdXAmcfT277uiytD8mZoAtPQAr8oQu4
lZa0fc3Ui03k8UVDk4rj5WQwRVQ+dT2oE3wkKYsqQ45eQzKSuPZdPrVCzx142czC
U51uuIlIY23qGdZuGcZHWkZTg6PGuxOJ2DbhwsqpR8q38u/K8j0AYhiwNfTiinEv
S32s4LO6VZUMtwaf50W6fh7xow3yiMfI4eapei1YwUKYMqflqqQ5d7G7eS9z5J+N
5LUBjzF5sHiXZUZ5CVMHy8E43eWKcbTOTt57E2MCz1jwlaS4xwTfUY5nsPf24Znb
IC3QKCNOiVzSngHHECzcYfTtLkuWKcQwTpDIjkdthsF/lNjfIc05D8YZmLTRXAaO
kYjOEvmFkzB9BNK3rx86er1g/9VEdI1tJs9bDCWtRNW7umGfbRGzwGEfJsUmDUWa
X/sUuYJHi/x0gutmKSatGr3peNCEwwBhLIzUotEZ8VdrICKpQOko8h3Spd8kfPHD
EL0gPC8+EHzBsy/sqUIP9/yLjxDHWLUnxCYid+5nxUm2BmOvnjkBwY1E8jsqaJyd
OE0+0wJahPTqxA3Fk+JntW6AexTraIgC+RunEmZom/Top1Cp9d33VUhL4yyZAikG
NuqjGc4ZtkqqJCQ352Uj/K7bH4vhvtg0d6MZVLYHpkv7K03U9X1cwfo3Ls1sUGOA
aHRg66XyZdZgy86mVnkkF0+d41rrW980oHuz4v+2S+/6jId+bH7VaIFo2FaND3La
n1fNyZJbFH0aNJ3SoJQLiM40ly/v+GjXW9M4ZENOXATC7EVoIPT4Yzdeks2nTQFA
T/joMb/jpYcJ4YiSci39Jl01i1b2GCRVEiU+kR/02iBucQUpx/vdu3CIhWaeJNe4
+L/0JnH8yCnTqUWeeuKHzzK47W9PVZNH2dAPEc3KyGxvqC+kBpPWR0kACIOpItD9
M5kK8SPvDu2mQshcaRnPM96DLWvLuqEnIU1O5HmO5isIK8dqYITDzI9tVUt7Tn5Z
oeSDIAlqtrdMNdXDOeiMkw79JuGB7zhBSp4I3GdIXEUuGiGZLIdN4GqZ22h31/Bf
h+hw0GcJSw+GpfrZUrxi1+hYfIPFTs1WBM+iEIjmZTnnT3JNgLvzjPil5SAVM3Px
DMWPf0nFUVz/o3IBU7zS/1A0V0TUt0GVNbo3JrGXWcmJ02jVjP5D7rCrS6mz/udR
N6QvHBkYDy/6DQJF1Y3CWpz+o1BtcD/+qHH+cs5kJorPwc4N1p5xtMw6zXgKcMRE
E2tHaTML9u0KnosF1FYsb1dHxaxJ5gZy37MnXfV2Cley+OVa2XcFdzgMv8d7IAVf
PDQbNYf+crwXBGGtxB8QD/nbcU0f9ne5glRx3DXLaeFDycbT9bWxf4oSfRpPKmsP
uU9F7pkcps9Ogw2o1IXq9+oZgulwqxxz6i+Nkb14PQkXOLyuSdHwll1LpD9hhFkU
fELIMs4/q1CN9X7JDltKD4YNvUM4D9m4MR05QuCvqE8mNBdfBu4ZmgedXL9eKSP4
r/hJC2POZa0pzBa5g5Nby4VtOvzWiHBoc+orOHXoTF/J0ZswAuLhGd1vuFpkOlzU
kUQdHYnshx35ShhGbT2044gG1TYCnav/zAPurCAsyDr/oyYKsTSy3N3MjQ32vADF
fCjk+rn4MhxsYnx9PQDSSSJ/c/+M2EM5R+qkjLOvFJEpgLBkp2FUR86IU96eQ76k
oc5D7he5smbjlKKYtPKSKqY+i2PYIo7PGJMcblJJyF2AMj8wC1MhXdlAAgE8jSoR
b9pgt5XAoETCNfTH31JdxExZIYE8DC+9XatTcM49448MfVlc3fxqbLx+Pkxfx6D8
mE8v3ty9fxhD9BRECHrXWMOADVgXb9LEsmPCykmCvOe9l8D56uTPv7yc6IT2RRV/
BlnvdLGPlgXONI76QJQcPOXq1szY3zbq37ub3UFtl7210o+nmTObr3BpHPDCWwnN
d72ACA08+kMTxtsjpqf5T2jIaDUWpGQPN5AqU38P4AxGhYLpeK7/N976URqoD+Q/
wwYdqHev9dvaDTghhvKXs2qcfE908cI7ynd9BTO5QlVSGAyw//LKkvPpZ9NPr4a2
hR18sYidllrkRPhtHg+a1Odeqk8c4zEKvwwvxfBDEYOeJRC4RR3fioHhaQsi0g/r
xbOfw2RaWHWycJygwGzdNiOxVGfxsdBORtGo4AExOWYjhQLUtGoZk/8JdiCguH6i
EvM3BYp/khmpK/HB7aMMdJV3jjtbbyzR7f+akdzwuh0fHB/wLkVpw7n0f6WB5k8d
R/QRxbI0Bs6dcEia+Blawwwl80LXdfszYNS3rhwmNtSlz1oZPQ0cRqoTquY9X8b/
EwNMM6ryt+HWTKqWlgI30L4VBifBhfgiwF45SccefTn1PD7j7c0uExokjd9s5W/e
iKtfXsH7LcMNiXf9USYIwuozIF+A38k7fb6eSvVJj2rQzzyvkZnLwhZ8Hrpr2GhK
LAfbeN3TQz7dSxkn7DxljhmrSgzL0zHHcpGkdkhgfb40fIiV29qgtK+T5tg/lGM/
TSdQKB6IieFdLsL8ckwE5HGxmUKK6nUWrVxBwFCDG55nLiRgH12mrWbl5+raYXu5
yzCOG0Q+HosqnLL0xV0kWp2madbw+UXhqWAvlBdXEF6ZKU0dUjTkQQm5d5PCuZzT
RX/VgJPD6lyrIY9sRoo09IdF6WcgFsNjhc21tZKz92SnhO+2LXCSpDsICcaW0AjM
AAGZ6qctd5OqF39Hv2RwpRyfU1ll5lkEUjOVKyU4lhQcGdpECq4OsdLwzNjX+qb9
msmhExqiUSu6ZOavMq+4K6BLTmpFIs4R6RksI9u0v/05x0/Sokn+YrGJitnzPFZa
ffwetJ1I/gyytUPolopQC+kxmNPdoIr05pqBJyqoEtbLXhRLErBa6ph/aGtq63wm
R2mOeR6tjtHa99AO/nVO1AM+uaanhY/cEU+L1iMdc4QJEJYE4wuHfAvkkyCsGldF
Md7IQEZHk7xEJ7WtzJeEMy2SD4GuqyWsocLPt7ykrvKH5U6ecrWRW31nU8tasawl
BrU8NHOE+jAdwqHIfzvXR9QZGBXvRnsKUgcdnO9zK5hsM30lebRTl+1e+bvxDdt3
jAKYpdXKGqozS2xHi7VRqIms1naRLIpg6O3VVG+Q0CFAK6/MMVlAP62OMXMjWnkx
WFzSKfVPz+c+EmxFS7mIQWN87Nkh4ihjuCp7/YlrKW9iWCkB9mWuaKlC6JLbpEpc
vpkBZqKPnJH8Owc6dYMm1Mzg/m6zoxJi0qCew9P1FMQwiKgMdHEYU+egxUNf3f1Z
RA8aHeF8cApg/q4CK5q/gwFAXXvPbV9lzWOyWVwli7+GIPAipC6hAXcStz2c9Sz7
daqZgyCcoXYF3n7ktnwQfebBb34mkLNpFyqYjjEikQs3X2mHvIko+/O7t7sKtY5n
vuWseKCYEcKFzqBglmDEXFalNN8xNi8q/RcZnLksiGNx3kmcGCFQhGi/WNaT6tzr
NZgaxdHdpPt6npMlktg5gxdD90VwxW50mv0cAQeuP8Ln+Kb4gcaVBOl0vA+WcwKZ
jpHLdEdJHagGbqDjc9VqGDny+w/gh3NQMU8Hdl24hSBeKuQES3A4Vd+/574oa1vm
/8y7lTgA1ssmH8Wb9F7Qd3Yl1XtT2FrjCbK74tYrVhKW3tBWtADNLNd2dHdkq0wy
ESLcPng83bO09vUzJ6Pvfys90RG6pxSEtk2ZgqRECmUOvXdWiAJuHhyxJ868t55L
/Nj+6dz9QvPOpnbRp59ulw2RcpInMtLnYyo9Dlxii1a13ycvV5nC2fnqQxBifJnu
6bOxHKa6M/jnFGs8NSwgY02Q3TZu4vm3uVdIVLV6d2RAN1AdNoGeFLYSdP8uZ98b
fIuPwQm3q3KAosX3OMAWnUpdTJKNmaNYRIRP5fzFF1LuLPKvi+M4UHkPzAhr3hDn
dVp4D8QmVyCXkErQOYDkoVGE83R4zpixiFCYZ15EkCOXCXHbcnDtRoI8rE1rk5oo
TRCuZbnm/6ydwXZMyg1h1J6y6RFMrQqPMAY4YeJ5DKzrF4fWmDjfsivbmnEfvog3
kNLPRrOKNcsT389StZlYd+Nvjd4AZ9s1inFxtc0KBs33xvAdr7jB6UI4hNza9OIl
08zk4QlJHRxqgf0omx2FOHLWFm8p6Nl59hMec+TMKOBBjw9hVCPnQioauZ8wpnHh
iWm8FNCgxcR7MnBqiZJB7CFrbA1MhNOGvsvSaF2X6XwpazTJn4Ggo0ZzHWt3ZXjH
AMg5jEcIgD3yOVbHewN/b5iIhLb+TYSZ3Q3TGOR7i2m3gSUdtcR9bZYWGRWQ+SKE
`protect END_PROTECTED
