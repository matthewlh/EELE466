`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
Tx1G/WPgi4VEdUr0PFUVmeIYSWbyDs7d1//Fq1J/HOEOxHCzt092V/OJ9GA6qXNj
DYY0xME5bQuP5FYUj3hhhmLKq9DtArmwvtBp3Ay6ltDHvisMWFS9zXgOD+vYqoTB
8nx9J1dkPePesPotQgcvGc5W25GSPYrFn1lnzqj6FWXtctJENS9ENaxl6R1ZYxJK
vgcHnifsqefK4BqTsvzfDWUkhtsqJBuboA8kwW6Z4TmCZTY1jCfc/HiNnDN1Xrop
6ZQds7dzwDV1p5x6iJJsn3miPmTcoN6+OMi7d/x+AmdBRpA0N9/1wPwv6jLNFbn7
1jyhkel5fod2Eun/RIuBPN8wTLUJ2WZoZoOptIwJcU5vVWLcy85Pf4ls1aKxvvl4
9p1ze7kYQmNRN8oEdmqD124PIual+u/BpRs69AmgYv0Lw+U0uY5HBOz75d5Jx5aK
825niza74QWwfmiI8NzVKpsDAqHCyM7f0SfLcVhWZUlCbBOLq6BbOvspzqI57+4D
2iwGKkxE/rAwQUfGx85/swApzD4igb3jsGlogN1923S/V+gAoGoLecbpiYC9ExDh
G6OxKQSQKyo3ZCbTvPShweGqeTEDpz4mnH0yg+C2uLK/O4hpja05WzIxm/gGcxmU
DkGqd/9Ay5eNn+nklP20JByKlHEPJysTIW/FqdlOvF2D+P2I/k6miy/1+TOngf03
W7oTTnPy15es2fgDkbZpSDJ4PZ2RQGGbPc//fS2OcH6AS/0SRciErdrC2QLziHrT
K8KfZJkJ9CnJARPK+P/5X8B71Bg2KKHbgKcRWxyG1ltA3bkVAb4FU31D6Ivszh5R
68oAthBIz4ZahJKb0eAYpmEMFtY77i0rjT2wKQpVE7372vRGMP2mB/XS0MENs4uO
fNP3rGl4X+nXxOVzbvw8/m86XrRcrY7LS0KrYmm6oc1e+7lylKSQ6AJnz2sK3fHm
9bxz0wUzPWIkJg0T8xmY8FeXN6xFMv+qrMwQw7S6ufrmn42QwyOUDdSbZWg0CFH7
Cs5iqmepKqwy5H4ZLEB2Rolus2MNxHT5kLsumFaowRfTpKb6lnpvri93fnLmyFGv
dOrmWA5nmE7kLzzHVOx6VDn0YPX5+PMmn8cunrASj+5JrJwsNeodXoxD9bI21Aox
B9FT0JqaPb2Rw54j7MZ78UpnQfd4w6wLtMz5xUdALgppa3AUfstFXOGsSxFhfd4D
P+oMV6uFVX93kQjLFkxW0Fira1ljCFgJquD/7qHbwl1l7LaEGmEJGiyC9nXPw5EF
qRRJYNm0rAzrnA3hsSrCqwuSS0EMPOi/f4PDZkaFXxWFo7KvgJiy2ydUxNd9MEYi
BipS1g4CMloUIKZsnI0PmTOl4TyGHH1ctMzrrShkTfARJ6q2Myzh7uGQNHQAMc5e
EtkACPZnLYLQG/9fcca3KCn3aSkf84mxoypV/eWnQwtBKPDNeIB9F/SNdor0rt43
u1I4KC8nJqbnCr6D37zShARZzBrFq5SgTDLVSx6hJCFIBbVroWnU1Q5TsElvHSw3
HSRL4WMsghhFHGrOgJtY4eSCQQtTZZ0pB5j27nWdXDCti86IRg99VFAoVJFIyGYN
pwBo+KAlBARmR7LtM6GRi91IGzgsYR/Q/eHMgHYx21M6xmjQCxfJpDv+yRwvC4gh
WjrMkkM8Zm7gRhDB69pv8KV9ZTU5suqiVcmunLWFKfj20vQRjGnFfFEpfamCPNg1
CpdhpDqLoR0TdoXSBn//ytoaooSkBsY5lEJI89rnkvxE6PKPvohGt7LTrf6C/OuI
R6FCMMcy+HKKlj5Rkab8U0rAS5Uv4WtdZRaKySJKeWihxqhCdTPuBMeV30rxErg3
W2liXA2ki9bOEOA/HFXq5WGuYGpdkn9lznFKP6u1JZ9q1r8Fihjym8EBzIzxr5kA
FbcEVc3czxAJwv6HZXGpYGtkf1H0xwWuKyIsvyuOU3hZJx9n4wLgamdv6X1NMz9g
/rKDer2wNd00JVpvsF1G/I/vzS6MYovYrTBAnT7m8Fms+lxBABhDwRGg0t0Ttb6z
yDzXZeJPPPkRPBwqKSGwKNbi3wIuqdE6HUBptHqgh3KCgYoVBOWX/qrik7Grelvc
Km6ZR89uGCuMEswYGI5asBPzcDqn9BD0li1ZJ/Kun4cQhSRISh+SWc9GfhWR8zj+
80Xa+5EkM266Yq6YDzUdgaKA+DNynS5jwH/WHpGgbff1OmQVpE1sH5WgRs8iurLt
FhREXlmia1qrZjJ+gayPMRRibYntOXbEV+vdfybwjuNXYm7H2xYYnYZxJNBywKgo
vGFPTdzbQh+ZarDQjec+OKJ6My0zHICZUhLLsaaDVxnHwUp6eiNEPasy1BzFlH8P
Du7DkCx3TnUBfYs4XeUjq0h5R+LpJv1idaJHYmXhCwOyVaijQMVsEE5P/HMZpKmu
9Nlm9Zw1OAalsV2lQJIngkjukvYmM9Xy1LVlwqk8t1WtDZrEyLRa+QJm3nMz8hn7
RVVLT91IPcSGJmwWA10NJh2K3ULY7spbTUBw2D8tI2QOY3uj204r4wnIzsL60/EK
2LoszH4PRqQnNNQ3B0nczoX++aZ9vyPgVtXs33jxpwHP196GEPzKv5WUxnizECD/
d1qkiwOvk96/n/ypVQSanUs8MU0LXQcUj9eB1XTNFe+5BJmA+0dg25U4b6H8P4Hq
9GWvr3mHlhvbOuDvDzUK6Y6heVostCA5plJeR3J2hZefpmtE6/D9Fua8A3lmWN/e
refctnJznjmJ5KA4eNdhtOSoRHMZgxbaXhoyQyPuAp3Q0z+S/vcXjb9i2QblehqT
rCKesX1jBzVwMz1zs6n1LRk33VMODxRE9lnVaQZgfxIDifHG5SE82MxdjdjMdOc2
FbMLF+vqyHmM1hcIgnGAkSUhX2F08TzyqIGUYzoR6t3Wydq/q397++gykNSDMCOJ
eLvTJhCp/fC3GUra9EEIReH1Oo52Z/GeayLE0W1Wygvd87rU1SmXJ0Nc9nEIzK89
DmvMzccWcp6rufO5ICeEk5DsFs4CF5tiih7g3nIho/VE+yL4/x4eyxLlXhTtGVIb
REy6wRoG4J/Vnq3Vu2nbNZTQp79nLwHOTw9VWWdFalhoPGjdRWT5+pOJ7KHY/VwC
3qLQ+j/2WINtUActATc6TeZG+15yLW/lld32x+lWNMjGASvupvcRAkVrBMnVgOsO
6AXHAQ27dN8bysOha9YKlrSIWF2yqlZ5f1sN2yUm0/i6h5/S32ju0fjheAqCysD7
R392M6DqC9OrH0iCcVfXr3/wWM7uNzqlcBvlpzZCtWz0tZvVVoLiTphvx83lZcdr
/ytravdbzjK9gzMbnbBhMLd7rxz7aHRniJ+vRzcGnKbVtz69ULoZpcwbv965DXhq
D9m7+IbZwHF0i8Ga84Y6IEMnTSddYyvjQvB7rCeRXyhQUDTEQxSxxW80VLTG6iHV
EyBunuqUxCveTbhKg29M+/qHBf1nG38XWGFocKVdwAgTvISHk2kZIMGHyfnZJBWa
Oj+incmeZqYPoAbRxcyp6wunIFCIPiHKFQhJMawZ0qnbGNgkgNfdSDjfUegMGVpI
ONVCg/Ph7Gyc6WcxJaSSCM48yQ7jX818v1jJLlCY8BAfu529bzFu4gXssUtgmtuy
ydFLPlGxoVEUfesJZ6D9AuBFSxVfSrRGfA2IQ+zuPi8X6IEllOEv97QrtakKjARQ
bQTjp5QgRwkw8M9yjXpDF514JN7JJaSofCG56e1qCmwRckSCHJzdeBdlyk4qWzP/
pILb1qrLwSE53MWDoqiczDCay23uHk1lMjtLXLto/BeHb694HQFgnHkOsNQxTn7w
dnfN5wEhm6S5OAK6lCC6DeaKv9/glyhoHE2aWX+JHX3PBXIxm+8X7RcmSPp00FuT
Vv8x4nXPTjJmt7sBfvU720XECQCbu+5mYvYMGSkeTpt5yCfn2ov+NKsmJkNNqHFO
g3keUyHEO++TjGQNie5qrrjhfk0tfEX8T+MNs4bf6e3VkR735pAq+sKBNvs7IY2I
P6vdaYded1E898s80hO5Bvnoyjzz9rbSKl19zNlwT9r8Nq37jpG0EYiqIO7o0NAy
tr3vQGoioKcx6bzGxC6UoAvcktoBHjTobR0KGmu0zTKGZZdy8Yj2J6WTG51fs/R6
5MXHTOnXe9Q2wZIrkWWpzFwMdrcC5mTIpg2AgdvQ8ssr6dDUb5j6/RsVEIQKVtVv
tvAjqYWDCVGW90FcyO3EeBrHH8Y0bnf7XV74PFc7rT4sB/WCe/mPjxhSuwvc+1TQ
3bzNtBMWfbmKNmEjwv1IPq8oBqEiuBkZVSLuqBh9jU7ID4TXNv2FMUFvbwkolp5J
lE/NHn4G2oyc5t/xifzVqgozNsoKAFUXc8n+183ZuwpVB0vaae8c3Rp0Lc4G8va3
cPup/Ra/SqfDAcjl9tpPj98cJAt51yNqBZp3sHRoob53GhcgnjviSIZV04Y1IWtP
z0Ga+/i7IEBoH8kmTjPlH+kCb7lwkV3JCq9svh8fTW5/T49I2zjLnUDpMFm0XfTM
63SO+Zr0s1LLSxF0/hsxCDjs0k5l6bslr5cqwks+ucrKaOR0dI23NiAR7Rn8rbiz
ERFg59oaSg73DV65TxDIXO/lrZ43narFfk1boZ8Ng1kLbLp0DuamwZB9BzPf3ImH
LDKRPUqM6O4WqAaaCJ8LXwkOlrgEbWw2ZtDdRTuf9O/SIEEdtzw5lq7nEHe6SL0k
2TH7zQz2UdBg4f/74dgeLi6cufSKx8mw6G+izoJP1lgeTHqyNk9iuwEBIQslm801
tqGhHzcC9lJEWDueeX6EFOj+dMorHC+eQ9mNtlAz2xix2XhNkvrthAqr/mQDW+w3
q8anKv+pRKw+quUzzCh+2jHEZd7b9TnYbck3Mm+CGqyq7yhi3/0+GLqzkSiJOf7f
vppiVIInDNxz/0Kcg4/rCil6yDsfNLTeeaTNxmC7z9hy3uCuTX5euwvGentV+XYU
ea7cgq19xw8p+Nr36bv+wxKhF74eOzhMhHk0wLhAvKkvxrqbtPaeS0550I1CCLFH
MmZ4dx4+3rDyukfk0JQroBeZ26y7rndNoCF44l6nvylVF8phC+UdbiWAn+b2Czcg
OO2cV+T/ArPnD2aKJYbwq3qd+hAUqZQgi90EiIUc7gpAbAomu4Q3boPs6ibYIQ9j
wsTiFYFliCLa1liXvDQPHqm5Eg7UTEKioitaSSVhZTnaXbTfhhZYe3DJxGUOQVjD
QmROygHxBOQV/F0o7bRHRw1wiV6yJIdS5DeMixLD+rfNodE+EJeL94Sc9A1AZyDR
BmbsT6iFcuK6DQ1Hgu3opSGeswBQ1VlmHFzeSLAlbJ36jqyP7XuBkpXyESwCQUk+
oUEdpCR81MHNDcbFPBs96tNxm9fsPgG2QSoBbFhp+0CwvRb0fWT0khuZs2XAbBJj
mw55bQ+QDq00/vDu7GwuUKaHPmz8vrTo4Ze62jXMAIVPI6wHBug8nridJYblmFVS
Blyszh1//YmcYg/MAJBaXDOgGc12Dd8BY2eJpnmpnh7Stk0zDBLzfqNFT/WPzMEZ
UCpKj6QVbfpQVe5R9lqU24jpqNoA2TfQH30JIWQeCmOU21ShJa99YeisJGR9zkeS
vJwBDGXlPAVVtgxKtYbnCOoWrPWGi46pw4AqABuNwCLzfn1w7wYFxHvjCQ7Wh/LC
O50krqw+Tt4IMRjoHJ89hxt8KWeTssQM03PEb7EuzFULjSI3uvxpKW6ZR56E4ZoN
N/+uKmYP33JEakogRbKNR9FUt85KQ5xN8EJqrooh4ziGf5MYypSA/aSgF4STsXUz
5xi9vG3R635vxVdhebseDexIjnpJFQ9v0YIu1MKy153CC2I8Xn1isIHMnOORsjKt
+54btqVE7AHtpUZfDQ4PRNL7vETjL8TdHUzU3TuXZX+lBWchi9y7Ot/+YqlffxxI
+0XwaBxFdSGfj7w2XcUN4VzwVM9WwqxIG+ZL1YsNmnxN4abxEa++ILRyJNeRvobO
bC9AC2pUqttNW+KaB3o/C2mWaCG7d8306lHSTEVqNiorztVv28eyQBnyKDJmpE/i
f2DCFOLOIjHUCpVZ6GH1n7aUJgT4i49fPgapk7eIzkPMJhIZH5xg7lTAucKIuwWB
h3AAIkcKgr7t7yIc/A5h5Ub3QD2E1TtR2n68trnqj8apPVU2HSJz8Zn9JEi9RFKI
k3aDAl2YWDZY2YDmaRd8cX0vTtg2EnPGHINInbfW7nkNdirmeyEMwr2Ix0iE3pZB
mNW1jgN49KlDfA+AQjVWyuDWUy1nLjgfrsAO/o+IdGNY1BaBjq/L+QwZtM3LxtIS
4Nqe+/N5mOpAo7a6EXZ6OEFWDsg8n+fYMeqpwD4gR2HLtZBZ5e3bv5kmgHv1GXON
Ug0xWJJFBLjzgKfrHar1LCxaHfj0bRadC4N9+bZD8ps9+FZknEl2do2dkE1zKqYz
MqBFPAGYBFBYCxjv3Yqd+MdNexyh8Mb73MlAFuUimIcdPL61ovVLYVqXqcUbZUZP
z2s3p2eq4Qxa1rcdtaxCRyiH/vzMf/uoRFeL77n7b1c5btOR95jsxZm5S3DldvCW
z6r/DBN1iO/Bp6oPey3TZFCKJWDQVEEa+tPIHUnOTl3DtPEjI50IHy1+u6eXQTti
oBSuq06drqxXaqb1cXivcPLEqksif3Dem99pyTwguMW4ctyoaPJehaQH4a4PDypM
aVhxMCaW9Di9RISb32NIr3wxx4trsxbv6ulCv0RF9hT1GCR1qY7cvaRnQX3Vufso
faUydTKrSMfU5jRYBbNjitu8HD75Jp9UxHPm19mh0migyts81Ict+izSxbLk5Kao
Bn0XYWxlczVPv5qcsZlUPUNdfyy/zN5rQ3VuBHjf7S15QDFWtlOjCrbNuPgf5Z2n
ZkMAp9oRJVgqWiUys3H4TgHx7ZYGUcdqDP/g9IQ7+dFC4Oh1ryKK9mrtRrlO/3aX
CE5kZI6qC/LfinuWY5HTK46jsEaHO0rfuHHocxYcYIS0TijA2af2CPNQv2BSOmPo
DfjHCZlRlfwBoskRoj6E5qDrSHdcIAXRTDSBG1SDj7TquclTpR/0Y2hMG/IkVSk6
QQHIjr84M/oiUC+L8Rx+HvYi/Ts/ggNWRUWzt2lsiKgUIUPgmBKbzoNqeBd5ba/t
rx1iUVDWJvKnbNFZhyIcrPYxknEbkaqbabqN42XrDNjWYQxG5pspqsBaKkudvmCT
fFPTeKyxqO9aB+76YopBHHjVZy9dcGoBVTJZ//XIb1vzB6SV3sFquHTplwmaFTg/
zi85WSILleAAfYR0UeKb7mGSPJ1KIMZOBpm6XyTK0sNtuKa7+6hjwUwNVFnDvgHk
SeC+wCuyCQsYxfv7JLhhn6jKs2AyPIGmFlyFS8ZAqM7qmj/SiJnnKm8KKwv1C9qj
ZWYGBYxkZL8yf/ucvySfV0z8TRlNLTpo4WQRTGq0hwT9KRYnRsFzFuPVfnon3R5r
naquL34cRyp3kGZRY0rrwSeFo+l7Fo2cknzBz4pH43K9V2iNKlTbXfZEBSnO3lTj
gEKA6wqkc1jzYiwdMxcNMFTGAviTJ6sf+QQgFjDn9Ocs8yhhKtAxK317nOvlksQL
yyk8//+C2mpVp3/TOn/OAf+aPiO6+X+l4LJclpPYZgpqrWC+IzhJ71X28jlXFw7u
pqRd7vwuQfUr402m9IW4UZoXuRBb64GUeoITHMD74RIEvJK2J1nBEQvHlLZIheW3
rElHdWYhA1/FQmPP5XqcvrzP6ahhIDogXzNEWvCIqCVnyx8nyvtGcp6Wp7N+JluZ
7Tiksibq4p2pANJeV9/++egHjnM4LnViYXnr58x1tdkNKBK+/6WNwzwrJmksN2nN
FJHlR25wzaNw6FW7iHVrZRgzoK7pitMaoPsBI5v8RWenK263mFdxhhh3r2oDt13d
Q3G6BdNh2O4ugJruhUWqIpLZZgl2qx8aIOyCuxj5JiHL07Mr6zs5Sgr6J6B2IB55
sMvIe0WgADyma+OkzupRIArBsnVzBoYW34ZNFEQVHKw8mQkowdDROFdlTiWjypmb
gK02xmX+TqM+A2w4Zt0hcrua4VRsfpbEgeu4SFDqRX0JP4iAN98cwcty4ZwT6gMI
+5KcjXcvLXpLXk/eQlhlD/hTNP0fyJpq626dBAitQfGyAluQgnGVy160yp75vXAx
cvlfB99yvS1erlHT3uZKIwKBGrduHPdAhEI+BVBp7wsTPlDcpyG1nHpWx4q6TgdF
hqAnzdAV6EconsEx/VSeR/CZdigWuQ/+RphsaWt8pKafQKAlH7hXzZ+pUN2+v73w
EOZbhgLIHiYDdVMeOJvFUBvOl2XPF5XUMSimBYW/mRomZJYt0X8nZb7rcjEBh3+o
9IO1i4U4QDKeJspprwVC/jOKyn0/BWLbcupp+TueH979IZdTYWCoG2NhYyHJ3mTx
ZNsRsxCQDrvd+7xgfWgnN5AAI4JVQdrnTv58y1RWRzBSmeuCI+hjvucmg4zTirKR
CDKcSrUHv1RvvFXovC5l6jNo+PqBuyIms+3bhfg4dDbtR/RUlcTEsOfqhHhJGF39
wBm6rsdTUBxL4HR4HMCW6jkKlYHwlHCmfmmO2swIpjfTGsMFh0ISPkOuk2UlhIBH
4StJYBekRO07Yxe22Z5KazJtBPpNHUuYdBxhSwWpwK+3ohpA6J1NzmKlAVrufr4p
iK5dG04oxm4tjlplsTLAPwHiasCJmXMmvwjsBP8llFiFM4oGatV+R9KLAuHX7CXI
mT07XXh/a6INmwYoDIPu8G67J3P0jFwmtK3nqRGVyYzwMrX93V8nd6dv29YGKZmP
plCpmcomTeK04ycHQ5PXg1ILTjvRRk69tpHijWBo+f7fbrcAlmqAPn1qSecun5AA
X889Ux8lWB5CKijeZQnSg4i1XBcFiuTydbVmyepvK56LEV1WwyJQHUYlIUX4dhO9
9lVKNHciuxLF6lYiEsT9s3OyiG8h2Kh4ja34jCDUiePXTdG/R8uneekt96y3hZFD
/OdIftTgjPDc/LnOJUsjqilxFSwVR8vxytj7W7IiJcmWpC18rdFL7qKGvNrPye8g
Dh0q1knkhrM5qynvxOItDoGhJVY/mVAuLyYqzJnzkc+uCD9gs+9v7B3VY57jyahP
qyTrOKl2IkxSbivs7UuKiFTd+NeixCxU8n7PLEF0e8Kh2K7E51so63Gq3Q2w1P6B
WJkPvV5WIIzJRPjBh8qzBsf43Vwq+oSk0tWnQ7OPqJJhS52WYkmgkeKiUEBLF5hk
Mz0uksvaxl6eaGBCRKfuQXzfd9xIj8B1oS98UEvRAc7/BAKnkPdDXm0JlqQrtadi
fP82dbRoubw3W9Gu4Ef1Wn6ULbBmSkglOpj6HDWsMgQmVUid/m1I2uEkK7r2426w
G2E7mzTJfmEWmsTc+jirTTNrZM42l8hdOpa0PrvwTy+Vobh0wTMxrHrownlMDF0e
25X546TDrl92Lbw4kFvkf4jTtcCxOppXPJtkAHJkd1dNdw0OvNy12YfCDsdThtRe
FZZaO8MqTQ/1RXsPPNP/CQ3/A3DreTxM5W66cRlLVBXBkEDMrSzjiatOAtWBOTaV
iRdXTZn8TiyslfjrrxnZq1mvgoV/LIKEcWj9YiVpkNw4bbV+BB4htiWBtwoQxZVn
3dbtnXKTUexWTdW+upGK3XVsLkLkjnKVlvVMHFO/jhk+o84wm6maOJNiVVjwjDKm
68k82wr1n+3Y77xadX0qx44PuK+yBIROP60xUGUmLX1IlcSrWjAYI5YI/yFE16BC
EcqjDSa0fgRpN0Qi08gdMPud5RW8SA3lS0nz6TATHHRvd0xb1To7CV1v+UsonlFY
dBOnJrrnmP/Db5JhDFjp5i+KKSIPiUyMNLadLfroxncWjWMGcWFLJsi+C9m9bxQV
jB8oPOstdqr6BDzRnnxiz4QV0Gwwzq2b+W+CdVz34tLSGDKQpqnzgJJkZFjnJiwh
eXdz+vEk44e/6GEp9/z3o6vvxikfZShmdFmNzXIeUfMhCfJcb6V7Vq0z5IeCNZPO
x5H+cCBkXuk1gF1DfnjvkKjlHA6hS7bXpOd6jg9TZBV4uAnBko4Dnj5xMD451R+/
9K/65qgtlC6M/4T6qZZ1kmHMfuVx70xCqptdG5cWQSO7z/RhEcxm6wk4xzeusNJB
6a8VTDHl7PwJVFq1wKfM+Wle8GEjQOMzByXqGJO5yvx2CLZBHxk9udbGROLu8Ylt
1rAQMyUeovKbLnDQsNv1ASZowbn2/oPanKkFzcOvCUchd87QbR4ihIT0C4ZyoMQd
GSvdSMPTqd5TMQz/l/PhDVmtjSk+cc6nemeCuuZamb4aucPLARuzTGO4QTKeB6rC
FR/Qhc33/WgVDCtaBgR+DDFRhbicej+1gyfUXg3i2po0CM6kG/Fj3ApDZObumssK
u0EQMqmT85yctdlooJ4pyKCt0oG5aOh6FP9/3kFSKOEhp4+1VsG9mzKEUjNwcuzV
SAmuR1Q8rSapgUmnf3Etwp4YvoJYhMhRkp2HICreR5lfoInXSGYgyXZPdXq1RbxG
mY9bS3Qm646njPltwTA68EXtTnZLTYUwxjLK0LVe52TcIqVfIPQ/ysG53kVwHhDO
L0ZCGmYwRQ1I3FV6EAVYSrDUraoVqmq7ISKcbfKVp5pX3t5nNzSu09hFhP6Tl4zK
wgpNBXvxz5r+8ZfMdCrm/9LwVTkwlxL3yoPbOt7yJceAW8ZVxrzIcSbjg92LirPx
58F4AAbzsiCqM9Mko+FK8ewbCBWpGicclpxEUfVp/POC/imgF/4S4C9nebSVfG/f
YkrPOe0BUuw12SuH67qrDP4q3f//JmOK04lWEIaUhQBftt1Pr8bjy7Nga+sbp46E
FvSfrybYob7LeGVPvUFEvW2ifS8ML0TmRYCSzcaZ9DEoHA3Ccvd8YZ45lkAaJ1hf
9RI4lIGO18//CCXE/8l49D0qRdotxMviJZDErCIbPnM+cFh7//tS11Y8UCCxqSKn
6Mhnkb+VbqHoJMZYkOrtfXejYUO64K51A52DUsd27+QV4jJbGIPLx3gjBGAiszow
Tb841bfbU1se5Ze+ogZ2TM5FzYDJLt7++/PCbbxPImf3bPVC+Ov1pP2Sm96W/o5R
wwHkOh+UZFe1VN7qNqusuCfiECFOoUbND61GdkD8Dr92ntXznTU0Kz76qDPhUq5P
MTuvPTWDmg1cxHdLRPpOOd2goy4YTcTyNv0wNC+YipskaZ49viAC44SB6lPthlDo
I2L9GGEJ1qed2arZw9//TsR0Bu9l1/2Fbz90v7/swfvDYRQzzT2OHs2dHL96xIKR
qYKAO5DD11GT6fXCrMtBagHXUTPmCS2mdQFZazAq4sLkR8RlWCMyCg/cqEU69FmT
bYxHVeQlNnrHJxOEsQMk4agyMQFc2RSG1rFxmO6Nw7i1LL4TVB0PEZQpWzWVZQc7
cUEVLf/cJQ/60WI8L+NazB3DNW2AIUNvjSOpAS11zjMyDFlsdjlhLraxQTI720pS
/72FkSbTSQ/MtDzDSc8YhuWCq5wsb31nBIocj00xXAK0cFY8Vix6wnSaBrCn/Vtd
r47kypmzqRth+zBPPnqxMPsTcReTMbowbYmsGVx/37nYC0Iy+rMJiuPXxX1D4u2z
Hf4/EnCswCdtBevKd5cbPhSJ0f54wsNxvJQFc9OxX5x29+l739ty7vCD5mkjmrdG
iQaXl8kftSF4oOxtFkD8A3bc1ub5aDWPFWLBqXL7UJ0lFdQY0RbtY9QWW5oRbWaV
PiJ09XyMqNW44JMBF1l+RczY2QAEJUDX9dBmBei1H3/5LlXmWP64Z1k8qRvWkk2J
hrAXY0QsU4Xwho88HgXPfolA6wqs0l6yxGRHXQk9HaB7TbvpXxy5/Vfm+Wi2JZyn
SfuKG9mW5tderdS1KO0WBZZRAD4/W9wg+2vNewlyviu9uE5adcCR11R2vYA2WlCc
NSEc9Cd4Qu//htdCr13DrtON3XL6ouYeiA+01RdfRlp0JX0GjAJqOopy6LvrDLEI
Tf0PUQGxPHXVtnWrvf5v4O2VHg5qEo+7Qn2adN2qBh1VT3SUJ96mlvuEJfmUKEU5
VIrMuFVohnQuhHZcTcxxtO112DUciTy3V3y6UvFKMQCCUqkYRtxUBzwP0HZdImwU
KSpGfSb4PT5kFJVL+RYN/qnACs/Sg1dP/721xKSrjLUNbzxOD9pdMkgzAGErep3W
FojbNTbIwrfPRcJ1wlqgC7AqWjh2uE1u/9juwByHU9+Jaz/wRkwNU3j6Ac65u5Fo
lDsKegKOr4LfNTOxV26G+hpgwJ/+8Wj8BCsuyHXSTpTuNVVOIojD0Hba3QZpVOYQ
3Q3tx8rO7CXb3QlwGqAbKl1jFq8cbM8PLwUXIV2jcOeevMjFhwtx0MxfbkYUAAF9
BzBLWeKQuWLRZtRfphJU1YlUpo8eP73/ds+dE85bIKFr9UTE1SjKJbmaADC3GP1y
NJha4qxTMlUZsfF+UrcshghQbQf/4dfjtMIxW6cdwFU=
`protect END_PROTECTED
