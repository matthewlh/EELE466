`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
fxy+R8NrzandM1rv/qjrh0MQgqiEm3M2Olhx81DHXv9F0P5vaSr6k/s/lyJIcZXF
dAB+PlAIPSMVy75M+AciccYsLwooQekGiBMNBJvEaPeVnRdlpy7jvk/W9EvipzVF
z7HtvqROgAuSLdAFwkDEM+dBEqajF00iqej5x9jzPL7lZb/v2yqTA+5I1poNabKF
GBXj0opnafFDnnDTg7rJUkuv5QLqHpmga0GvmfQtnSrgJ0RqtjGZiQDiGVw8MdeS
avZCwmVN2SUvNQHhNtVu0yiKKTPuZDlV9tXXqvXbxqnp25aryia1nPlFaTlZXGCO
pUUJXZE1faaeQw+eKneQn6+66tQesuDsaA8qh/1LMyz4jtTXsnj4aS+UpvHqCi12
XYzVokXMZPYzHytkEJXq6dgvTcSl01OvO2va4OIhLl/4oWDWh81OJFcUAfuls+Br
4lV2VMTHDkRZdSX6iZbjHxq68vT/21hwnppSz+j0s5oE9Edj5Jo06RGxxAtFVuxV
m0BeF+1Ehezoql4XfJcFOkX/tmhQQLiiy0U7PK2Bc45ARQkfgEhxuGJwY7/T5QzN
+huLjb7YpOFzDlq1KnbFaVOOMRAGiMu4EIkBR2PtO9K7cexSTXTpF07P/WByu11v
d8pb4nxHsAtFXZheJgwvLqDmwW44iIssEKffz983lFD86qMAjYoDkRw10l9uiRO2
v5qp7TLI/GjeGyax+vh2ms8N1Hv0FPsOeC2piA0Z/v29GSIlnS/nuuWl36XXqZbE
OQBAbCntJkQGEcsOlDje2geyCbpKHEXE2o99Qmd8PBfGlwy713+r3ejK73qU+Iw7
FKdOICa/wfEkRdfyw1CNDcqOyCsxLuZmUuwnznXU/mb2b3IHh5vDmHX/ke/0yKtW
Nps0eWDkegKGzsh2cSHLLfbW6dgh/9bKvYroesXN8kR1H+oUclfouJ54atJ2iGZ6
6IASXTamuROfZZ227mKQp6BqSKB74z3UTw6d62IlOnWSZ5gRbMrB/6hRUthfZQRY
pabYXoTJnBZ87UAJaysHOgPIkHYL7f9gF2k8V+deu6VqvF3hFrVaVJ5Af898viWz
AfhlCSOrpWwTyKsZhCcl1SpEkYzccSHoS4g5w9IVJjtD+mbI9E4AaeftdBegTMsY
rQlGU+WUns0ymbZBw4Sirm+30Xn56ls3OaS+l7vSereQuPgAfwf41x7qdmSxz/kp
jjHCkjYSABAVTZMoe4Sc5kEwzdSYD9qTLDotAREVELQB1C4SHls1jRURECItWXp1
1fTkoARWegKjuLK5JRXXh2iK1/rrHnUczVRJ422Ripp5IxFIRfa3mJ/FGPpLeNO7
+CYPjyOIaPe7UxxcX6b6KN9E+RiPnegKoTua+AcPDvIH3tvYfi3pW0mrpgPhGP9y
peJaSzAvof8q9oPDpnzQQxV0I6mXmbHTYxXdNWqRRtHw3j0JzaTGnj9ubvTOI1UM
b3Jk10L2WWwbxmDFphfz4aLFyScQw5BUcdCDN6qJam055HKytjPWI4gSYLiR6N0M
h5I+Is9jfJ01XyVSZNTBSlnYq1kPXuMbmPEIvOdXLsfJrMYJ8Yt3hfQ6RgNequ/P
rvgdxGWWg6JlfOA9SkZNieRb23jZrKIiCJj8QS8yexFkRuMCpvC3q2XDqIR7okUA
8C56sb0qHkbj7H2BX/EH/V+S5+A4hx2BpTNSqVrnxBWTe5a0QceRnfMiXqD/ayHq
ew/DRzoufhmvwaGIkEO3g3DAtpFYcTACw4LOUdIP3W4qtzWeh/47hplaKnS/+Jqm
cjtWggdbrXeFRY23H/EN04rJsNGmZDpPe/gAzJokopvPAabUHn7C58SrWC36iJdh
esCwU6I4tzU1V1fSoGnEfSIYtqWFK0tQ5gbE2H5freREdzf9yi8eSqYDOM31svMC
2wQZW/bmVHbayVSH5WSquxIMVqiVbzaI1dO8xa6qgNjBSSthito7XwvJLXYzNy9f
VkSfHlUdUPNwpbOUH6cypPtqxrDebXQL7rDhnz+rvzIYHpqYEg3qWBpPFtcLEvfu
T8iSjmSMZadpcKSFi74hIsx8SvwfflEZdRK3yryZ2EVsawJLqd4RARW+TPQrInt+
ZoBkhQ5lBVVWrsYRctsn3jUBAy5Y6Jnux3dbYbR2J4e0nkIrzDqe+D8XF0DwUUY1
Z2bSlNnKmVMHWHrMYyyYO9g+x12kXZO0BNg7nxkuG46gFha8AIsspQasYUw16Plo
6way5K9beE/Zv0xzLUsiNSPN2sPBTKwn7TKN7f3/R1ATBmS0m00nACfGrdVSOAyJ
6Tzvd24BNnv21lPVlMTH0ELd92en6P9cVx3sobFFOteKybR7POHtUQ9oKZw+0qjT
q2zLC44bFMar9sk7fT29UGSC1PUALV5KzM7iFEPd0Hw+VnW7qJ0jdPrN3QC7/yad
/8KoJ/pnvbILoHfeK1pdP9uf8/SSVIrGhAsoue9e3JodpcuzMzFPj1SzmTfsdMgy
+SpaX3jPi48Z+kgBmefOAsZJK3s6JCBDEq0aC+jgIKaGmyyXzq6VhBqWdAoATcMn
EBmAMZ+3v76lLqjQeh1C6JDzhWD6qCT5T7lEEOUslL4=
`protect END_PROTECTED
