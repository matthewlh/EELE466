`protect BEGIN_PROTECTED
`protect version = 1
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV"
`protect data_method = "aes128-cbc"
`protect encoding = ( enctype = "base64" , bytes = 168 )
`protect DATA_BLOCK
G8S7XU7wIUfsUKIA6zT0GcvEm1kdxdaa+TB+3/uGpZEAXLEsnRUEncsOYHC8Jtns
IjD4SCVAD60kYhxQDpSy6QrIt+el7W8XjmmsOyJ5idgq+rMVbRDvs2ju8y9h8QTm
qAWQ/+InXE8v2ESutgiVxR1xIVqsouXGCmNo4iO3JARXVEi+3vLwrNfTQoB14Gco
Rjj0iuM4tQDrxOh84PZuy6/d42jTOUlWHDRRV5Zk9cUjcr6+Cv4uhhtHh5cfPwdp
QxQ8AwQac9hDZTNYYYwYC91YJSUTdeJYuRCjPMTxZWZHsqCF+j7fqnHZ59RGbA/O
pN2o60Qlk1rFuJPysg2h9vEuA4NjblSgQ+ellmY5OEaPijCbx7TomaChekFA4cT6
MDUdcS/LKreSc6DxDlI/VcX8LZiYSheDOPB4QL8sGaE8AJcRCFtNu8TOE8Ky0PAx
wqMQmJhUL4Og0HLCu8OeUzlUPBCaEWBA4Vs9fFqLVe8h21MBCt5hCj2qwr9DhsXA
N+C3tlDic214VsZ57iDJ+1YSzCNZQRhMmwUOLwdPnrXArLLeAj0K8IIByz0rRLtq
gVyBbhpyIGYCcEwHw+lfAryyncsFIUSO81tMGOUKotMCdHK1fuVW8KRsdd8djBC/
4+n0XURDrQ73PJ+vOAtmTqP+vCSLof1Gg6hvlPcgHa7+6/cvFJHMVVCEM37mQ/VD
rOHb0K/UoMSeSA7SaNMgFq8RFl2mk0W7kbiZX9osJVs=
`protect END_PROTECTED
